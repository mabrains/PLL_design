** sch_path: /home/ahmedelbadry/D_FF/conventional_pfd.sch
.subckt TOP
M1 net1 RST GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=2.5 nf=1 
M2 net1 REF net2 VDD sky130_fd_pr__pfet_01v8 L=0.2 W=4 nf=1 
M3 net2 RST VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1
M10 net4 FB net5 VDD sky130_fd_pr__pfet_01v8 L=0.2 W=4 nf=1 
M4 dn_b FB net6 GND sky130_fd_pr__nfet_01v8 L=0.2 W=2 nf=1 
M6 up_b REF net3 GND sky130_fd_pr__nfet_01v8 L=0.2 W=2 nf=1 
M5 net3 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=2.5 nf=1 
M14 up_b net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 
M9 net4 RST GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=2.5 nf=1 
M11 net5 RST VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 
M12 net6 net4 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=2.5 nf=1 
M13 dn_b net4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 
M15 dn dn_b GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=2.5 nf=1 
M16 dn dn_b VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 
M7 up up_b GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=2.5 nf=1 
M8 up up_b VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 
M9 RST dn_b GND GND sky130_fd_pr__nfet_01v8 L=0.2 W=2 nf=1 
M10 RST up_b GND GND sky130_fd_pr__nfet_01v8 L=0.2 W=2 nf=1 
M17 net7 up_b VDD VDD sky130_fd_pr__pfet_01v8 L=0.2 W=4 nf=1 
M14 RST dn_b net1 VDD sky130_fd_pr__pfet_01v8 L=0.2 W=4 nf=1 
.ends







