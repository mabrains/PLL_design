* Extracted by KLayout with SKY130 LVS runset on : 17/11/2022 14:26

.SUBCKT integer_pll_2 VDD dn ibias_bgr ibias_cp up ibias_vco vn VOP vctrl vp
+ vco_out FB modi P7 P6 P5 P4 modo P0 P1 P2 P3 REF GND
M$1 VDD dn \$4 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$2 \$15 \$53 \$19 VDD sky130_fd_pr__pfet_01v8 L=0.6U W=66.6U AS=19.314P
+ AD=19.314P PS=139U PD=139U
M$5 \$9 \$53 \$122 VDD sky130_fd_pr__pfet_01v8 L=0.6U W=13.32U AS=3.8628P
+ AD=3.8628P PS=27.8U PD=27.8U
M$14 GND \$11 \$280 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$15 \$107 VOP \$280 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$16 ibias_cp ibias_cp VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=40U AS=9.5P
+ AD=9.5P PS=61.9U PD=61.9U
M$18 VDD ibias_cp \$174 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=10U AS=2.9P
+ AD=2.9P PS=20.58U PD=20.58U
M$21 \$11 up \$19 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=10U AS=2.9P AD=2.9P
+ PS=20.58U PD=20.58U
M$22 VOP \$309 \$19 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=10U AS=2.9P AD=2.9P
+ PS=20.58U PD=20.58U
M$23 \$96 \$53 \$282 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=1U AS=0.29P AD=0.29P
+ PS=2.58U PD=2.58U
M$24 \$11 \$53 \$284 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=1U AS=0.29P AD=0.29P
+ PS=2.58U PD=2.58U
M$25 VDD \$122 \$15 VDD sky130_fd_pr__pfet_01v8 L=0.6U W=66.6U AS=19.314P
+ AD=19.314P PS=139U PD=139U
M$28 VDD \$122 \$9 VDD sky130_fd_pr__pfet_01v8 L=0.6U W=13.32U AS=3.8628P
+ AD=3.8628P PS=27.8U PD=27.8U
M$31 VDD \$122 \$280 VDD sky130_fd_pr__pfet_01v8 L=0.6U W=6.66U AS=1.9314P
+ AD=1.9314P PS=13.9U PD=13.9U
M$38 \$282 \$122 VDD VDD sky130_fd_pr__pfet_01v8 L=0.6U W=8U AS=2.32P AD=2.32P
+ PS=17.16U PD=17.16U
M$39 \$284 \$122 VDD VDD sky130_fd_pr__pfet_01v8 L=0.6U W=8U AS=2.32P AD=2.32P
+ PS=17.16U PD=17.16U
M$42 \$330 vn VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=60U AS=10.625P
+ AD=10.625P PS=69.25U PD=69.25U
M$54 vco_out vp VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=60U AS=10.625P
+ AD=10.625P PS=69.25U PD=69.25U
M$66 VDD up \$309 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$67 vn vp \$472 \$472 sky130_fd_pr__pfet_01v8 L=0.15U W=250U AS=48.5P
+ AD=41.25P PS=301.94U PD=251.65U
M$68 \$472 vn vp \$472 sky130_fd_pr__pfet_01v8 L=0.15U W=250U AS=41.25P
+ AD=48.5P PS=251.65U PD=301.94U
M$77 \$501 \$439 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$78 \$502 \$455 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$79 \$349 \$439 \$571 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$80 \$571 \$352 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$81 \$352 \$501 \$572 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$82 \$572 \$421 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$83 \$354 \$439 \$531 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$84 \$531 \$358 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$85 \$358 \$501 \$534 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$86 \$534 \$386 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$87 \$503 \$467 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$88 \$366 \$386 \$513 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$89 \$513 \$369 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$90 \$369 \$500 \$516 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$91 \$516 \$407 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$92 \$372 \$386 \$519 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$93 \$519 \$376 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$94 \$376 \$500 \$522 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$95 \$522 FB VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$96 \$500 \$386 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$97 \$388 \$455 \$541 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$98 \$541 \$391 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$99 \$391 \$502 \$544 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$100 \$544 \$428 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$101 \$434 \$455 \$547 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$102 \$547 \$435 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$103 \$435 \$502 \$550 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$104 \$550 \$439 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$105 \$447 \$467 \$555 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$106 \$555 \$449 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$107 \$449 \$503 \$558 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$108 \$558 \$442 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$109 \$402 \$467 \$561 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$110 \$561 \$404 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$111 \$404 \$503 \$564 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$112 \$564 \$455 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$113 \$472 ibias_vco VDD VDD sky130_fd_pr__pfet_01v8 L=0.5U W=1000U AS=147.9P
+ AD=147.9P PS=1034.79U PD=1034.79U
M$122 VDD ibias_vco ibias_vco VDD sky130_fd_pr__pfet_01v8 L=0.5U W=200U AS=29P
+ AD=29P PS=202.9U PD=202.9U
M$173 \$407 \$411 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$174 VDD FB \$411 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$175 VDD modi \$411 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$176 VDD \$372 FB VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$177 VDD \$420 FB VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$178 VDD \$366 \$420 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$179 VDD \$386 \$420 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$180 VDD P7 \$420 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$181 \$421 \$382 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$182 VDD \$386 \$382 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$183 VDD \$366 \$382 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$184 VDD \$354 \$386 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$185 VDD \$427 \$386 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$186 VDD \$349 \$427 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$187 VDD \$439 \$427 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$188 VDD P6 \$427 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$189 \$428 \$432 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$190 VDD \$439 \$432 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$191 VDD \$349 \$432 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$192 VDD \$434 \$439 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$193 VDD \$397 \$439 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$194 VDD \$388 \$397 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$195 VDD \$455 \$397 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$196 VDD P5 \$397 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$197 \$442 \$446 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$198 VDD \$455 \$446 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$199 VDD \$388 \$446 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$200 VDD \$402 \$455 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$201 VDD \$458 \$455 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$202 VDD \$447 \$458 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$203 VDD \$467 \$458 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$204 VDD P4 \$458 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$205 VDD \$874 \$871 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U AS=1.45P
+ AD=1.45P PS=10.58U PD=10.58U
M$206 \$871 REF \$859 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$207 VDD \$859 \$872 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U AS=1.45P
+ AD=1.45P PS=10.58U PD=10.58U
M$208 \$860 REF \$872 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$209 VDD \$872 \$873 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U AS=1.16P AD=0.58P
+ PS=8.58U PD=4.29U
M$210 \$873 \$875 \$874 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U AS=0.58P
+ AD=1.16P PS=4.29U PD=8.58U
M$211 VDD \$872 up VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U AS=1.45P AD=1.45P
+ PS=10.58U PD=10.58U
M$212 dn \$875 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U AS=1.45P AD=1.45P
+ PS=10.58U PD=10.58U
M$213 \$875 FB \$861 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$214 \$875 \$862 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U AS=1.45P
+ AD=1.45P PS=10.58U PD=10.58U
M$215 \$862 FB \$876 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$216 \$876 \$874 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U AS=1.45P
+ AD=1.45P PS=10.58U PD=10.58U
M$217 \$611 P0 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$218 \$611 vco_out VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$219 \$611 modo VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$220 \$739 \$611 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$221 \$739 \$622 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$222 VDD vco_out \$614 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$223 VDD \$739 \$616 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$224 \$616 \$614 \$618 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$225 VDD \$618 \$620 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$226 \$620 vco_out \$622 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$227 VDD \$634 \$624 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$228 \$624 \$614 \$626 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$229 VDD \$626 \$628 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$230 \$628 vco_out modo VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$231 \$632 \$652 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$232 \$632 \$739 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$233 VDD \$632 \$634 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$234 \$635 P1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$235 \$635 \$739 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$236 \$635 \$652 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$237 \$740 \$635 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$238 \$740 \$645 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$239 VDD \$739 \$702 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$240 VDD \$740 \$639 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$241 \$639 \$702 \$641 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$242 VDD \$641 \$643 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$243 \$643 \$739 \$645 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$244 VDD \$656 \$647 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$245 \$647 \$702 \$649 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$246 VDD \$649 \$703 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$247 \$703 \$739 \$652 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$248 \$654 \$675 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$249 \$654 \$740 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$250 VDD \$654 \$656 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$251 \$657 P2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$252 \$657 \$740 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$253 \$657 \$675 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$254 \$741 \$657 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$255 \$741 \$668 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$256 VDD \$740 \$660 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$257 VDD \$741 \$662 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$258 \$662 \$660 \$664 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$259 VDD \$664 \$666 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$260 \$666 \$740 \$668 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$261 VDD \$679 \$704 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$262 \$704 \$660 \$671 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$263 VDD \$671 \$673 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$264 \$673 \$740 \$675 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$265 \$677 \$706 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$266 \$677 \$741 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$267 VDD \$677 \$679 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$268 \$680 P3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$269 \$680 \$741 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$270 \$680 \$706 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$271 \$467 \$680 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$272 \$467 \$690 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$273 VDD \$741 \$705 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$274 VDD \$467 \$684 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$275 \$684 \$705 \$686 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$276 VDD \$686 \$688 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$277 \$688 \$741 \$690 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$278 VDD \$701 \$692 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$279 \$692 \$705 \$694 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$280 VDD \$694 \$696 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$281 \$696 \$741 \$706 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$282 \$699 \$447 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$283 \$699 \$467 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$284 VDD \$699 \$701 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$285 VDD \$18 ibias_bgr VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5U W=200U
+ AS=30.74P AD=30.74P PS=273.48U PD=273.48U
M$317 VDD \$18 \$18 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5U W=44U AS=6.38P
+ AD=6.38P PS=56.76U PD=56.76U
M$357 \$31 \$18 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1U W=40U AS=8.7P AD=8.7P
+ PS=60.87U PD=60.87U
M$359 \$25 \$31 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1U W=40U AS=8.7P AD=8.7P
+ PS=60.87U PD=60.87U
M$361 \$36 \$30 \$34 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5U W=90U AS=15.225P
+ AD=15.225P PS=107.03U PD=107.03U
M$362 \$34 \$25 \$37 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5U W=90U AS=13.05P
+ AD=13.05P PS=91.74U PD=91.74U
M$381 VDD \$18 \$30 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5U W=20U AS=2.9P
+ AD=2.9P PS=25.8U PD=25.8U
M$383 VDD \$18 \$25 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5U W=20U AS=2.9P
+ AD=2.9P PS=25.8U PD=25.8U
M$437 VDD \$18 \$34 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5U W=4U AS=0.58P
+ AD=0.58P PS=5.16U PD=5.16U
M$589 GND dn \$4 GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U AS=0.29P AD=0.29P
+ PS=2.58U PD=2.58U
M$590 \$258 dn VOP GND sky130_fd_pr__nfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$591 \$258 \$4 \$11 GND sky130_fd_pr__nfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$592 GND \$10 \$62 GND sky130_fd_pr__nfet_01v8 L=0.6U W=20U AS=5.8P AD=5.8P
+ PS=45.8U PD=45.8U
M$594 GND \$10 \$57 GND sky130_fd_pr__nfet_01v8 L=0.6U W=4U AS=1.16P AD=1.16P
+ PS=9.16U PD=9.16U
M$596 GND \$10 \$58 GND sky130_fd_pr__nfet_01v8 L=0.6U W=4U AS=1.16P AD=1.16P
+ PS=9.16U PD=9.16U
M$599 GND \$10 \$63 GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$607 \$107 \$96 GND GND sky130_fd_pr__nfet_01v8 L=1U W=1.3U AS=0.377P
+ AD=0.377P PS=3.18U PD=3.18U
M$608 \$96 \$174 \$107 GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U AS=0.29P
+ AD=0.29P PS=2.58U PD=2.58U
M$609 GND \$96 GND GND sky130_fd_pr__nfet_01v8 L=1U W=1.3U AS=0.377P AD=0.377P
+ PS=3.18U PD=3.18U
M$610 \$11 \$174 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U AS=0.29P AD=0.29P
+ PS=2.58U PD=2.58U
M$611 \$62 \$174 \$258 GND sky130_fd_pr__nfet_01v8 L=0.6U W=20U AS=5.8P AD=5.8P
+ PS=45.8U PD=45.8U
M$614 \$58 \$174 \$53 GND sky130_fd_pr__nfet_01v8 L=0.6U W=4U AS=1.16P AD=1.16P
+ PS=9.16U PD=9.16U
M$617 \$63 \$174 \$10 GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$624 \$284 \$11 \$57 GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U AS=0.29P
+ AD=0.29P PS=2.58U PD=2.58U
M$625 \$282 VOP \$57 GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U AS=0.29P AD=0.29P
+ PS=2.58U PD=2.58U
M$626 vn vp GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=100U AS=19.4P AD=16.5P
+ PS=121.94U PD=101.65U
M$627 GND vn vp GND sky130_fd_pr__nfet_01v8 L=0.15U W=100U AS=16.5P AD=19.4P
+ PS=101.65U PD=121.94U
M$636 ibias_vco ibias_bgr GND GND sky130_fd_pr__nfet_01v8 L=1U W=250U
+ AS=39.875P AD=39.875P PS=278.19U PD=278.19U
M$641 GND ibias_bgr ibias_bgr GND sky130_fd_pr__nfet_01v8 L=1U W=50U AS=7.25P
+ AD=7.25P PS=50.58U PD=50.58U
M$648 ibias_cp ibias_bgr GND GND sky130_fd_pr__nfet_01v8 L=1U W=25U AS=7.25P
+ AD=7.25P PS=50.58U PD=50.58U
M$649 GND up \$309 GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U AS=0.29P AD=0.29P
+ PS=2.58U PD=2.58U
M$650 vco_out vp GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=4.2U AS=1.218P
+ AD=1.218P PS=8.98U PD=8.98U
M$651 \$330 vn GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=4.2U AS=1.218P
+ AD=1.218P PS=8.98U PD=8.98U
M$652 \$413 \$407 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$653 \$349 \$501 \$422 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$654 \$422 \$352 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$655 \$352 \$439 \$423 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$656 \$423 \$421 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$657 \$354 \$501 \$355 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$658 \$355 \$358 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$659 \$358 \$439 \$424 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$660 \$424 \$386 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$661 \$388 \$502 \$433 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$662 \$433 \$391 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$663 \$391 \$455 \$360 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$664 \$360 \$428 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$665 \$434 \$502 \$361 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$666 \$361 \$435 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$667 \$435 \$455 \$395 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$668 \$395 \$439 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$669 \$450 \$442 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$670 \$366 \$500 \$412 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$671 \$412 \$369 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$672 \$369 \$386 \$413 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$673 \$372 \$500 \$373 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$674 \$373 \$376 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$675 \$376 \$386 \$377 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$676 \$377 FB GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$677 GND \$439 \$501 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$678 GND \$349 \$425 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$679 \$425 \$439 \$426 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$680 \$426 P6 \$427 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$681 GND \$455 \$502 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$682 \$447 \$503 \$448 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$683 \$448 \$449 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$684 \$449 \$467 \$450 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$685 \$402 \$503 \$451 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$686 \$451 \$404 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$687 \$404 \$467 \$362 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$688 \$362 \$455 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$689 GND \$467 \$503 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$690 \$611 P0 \$767 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$691 GND \$411 \$407 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$692 \$767 vco_out \$768 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$693 GND FB \$409 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$694 \$768 modo GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$695 \$409 modi \$411 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$696 \$739 \$611 \$746 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$697 \$746 \$622 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$698 GND \$386 \$500 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$699 GND \$372 \$415 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$700 \$415 \$420 FB GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$701 \$632 \$652 \$749 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$702 GND \$366 \$418 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$703 \$749 \$739 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$704 \$418 \$386 \$419 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$705 \$419 P7 \$420 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$706 GND \$382 \$421 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$707 GND \$386 \$380 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$708 \$380 \$366 \$382 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$709 \$740 \$635 \$752 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$710 \$752 \$645 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$711 GND \$354 \$384 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$712 \$384 \$427 \$386 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$713 \$654 \$675 \$771 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$714 \$771 \$740 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$715 GND \$432 \$428 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$716 GND \$439 \$430 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$717 \$430 \$349 \$432 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$718 GND \$434 \$437 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$719 \$437 \$397 \$439 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$720 GND \$388 \$440 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$721 \$440 \$455 \$441 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$722 \$441 P5 \$397 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$723 GND \$446 \$442 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$724 GND \$455 \$444 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$725 \$444 \$388 \$446 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$726 GND \$402 \$453 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$727 \$453 \$458 \$455 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$728 GND \$447 \$456 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$729 \$456 \$467 \$457 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$730 \$457 P4 \$458 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$731 \$635 P1 \$769 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$732 \$769 \$739 \$770 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$733 \$770 \$652 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$734 \$741 \$657 \$757 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$735 \$757 \$668 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$736 \$677 \$706 \$760 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$737 \$760 \$741 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$738 \$467 \$680 \$763 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$739 \$763 \$690 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$740 \$699 \$447 \$776 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$741 \$776 \$467 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$742 \$614 vco_out GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$743 GND \$739 \$778 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$744 \$778 vco_out \$618 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$745 GND \$618 \$781 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$746 \$781 \$614 \$622 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$747 \$783 vco_out \$626 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$748 GND \$626 \$786 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$749 \$786 \$614 modo GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$750 \$634 \$632 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$751 \$702 \$739 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$752 GND \$740 \$789 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$753 \$789 \$739 \$641 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$754 GND \$641 \$792 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$755 \$792 \$702 \$645 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$756 \$794 \$739 \$649 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$757 GND \$649 \$797 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$758 \$797 \$702 \$652 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$759 \$656 \$654 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$760 \$657 P2 \$772 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$761 \$772 \$740 \$773 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$762 \$773 \$675 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$763 \$679 \$677 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$764 \$680 P3 \$774 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$765 \$774 \$741 \$775 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$766 \$775 \$706 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$767 \$701 \$699 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$768 GND \$874 \$859 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U AS=0.725P
+ AD=0.725P PS=5.58U PD=5.58U
M$769 \$860 \$859 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U AS=0.725P
+ AD=0.725P PS=5.58U PD=5.58U
M$770 GND \$872 up GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U AS=0.725P
+ AD=0.725P PS=5.58U PD=5.58U
M$771 \$874 \$872 GND GND sky130_fd_pr__nfet_01v8 L=0.2U W=2U AS=0.58P AD=0.29P
+ PS=4.58U PD=2.29U
M$772 GND \$875 \$874 GND sky130_fd_pr__nfet_01v8 L=0.2U W=2U AS=0.29P AD=0.58P
+ PS=2.29U PD=4.58U
M$773 dn \$875 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U AS=0.725P
+ AD=0.725P PS=5.58U PD=5.58U
M$774 GND \$862 \$861 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U AS=0.725P
+ AD=0.725P PS=5.58U PD=5.58U
M$775 \$862 \$874 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U AS=0.725P
+ AD=0.725P PS=5.58U PD=5.58U
M$776 GND \$634 \$783 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$777 GND \$656 \$794 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$778 \$660 \$740 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$779 GND \$741 \$800 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$780 \$800 \$740 \$664 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$781 GND \$664 \$803 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$782 \$803 \$660 \$668 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$783 GND \$679 \$805 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$784 \$805 \$740 \$671 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$785 GND \$671 \$808 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$786 \$808 \$660 \$675 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$787 \$705 \$741 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$788 GND \$467 \$811 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$789 \$811 \$741 \$686 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$790 GND \$686 \$814 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$791 \$814 \$705 \$690 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$792 GND \$701 \$816 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$793 \$816 \$741 \$694 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$794 GND \$694 \$819 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$795 \$819 \$705 \$706 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$796 vctrl vn vctrl GND sky130_fd_pr__nfet_01v8_lvt L=8U W=17U AS=4.93P
+ AD=2.465P PS=34.58U PD=17.29U
M$797 vctrl vp vctrl GND sky130_fd_pr__nfet_01v8_lvt L=8U W=17U AS=2.465P
+ AD=4.93P PS=17.29U PD=34.58U
M$798 GND \$36 \$18 GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5U W=4.2U AS=1.218P
+ AD=1.218P PS=14.2U PD=14.2U
M$808 \$31 \$18 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=20U W=0.42U AS=0.1218P
+ AD=0.1218P PS=1.42U PD=1.42U
M$809 \$36 \$37 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5U W=1.68U AS=0.3654P
+ AD=0.3654P PS=4.26U PD=4.26U
M$810 GND \$37 \$37 GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5U W=1.68U AS=0.3654P
+ AD=0.3654P PS=4.26U PD=4.26U
Q$817 GND GND \$203 GND sky130_fd_pr__pnp_05v5_W0p68L0p68 AE=3.6992P PE=21.76U
+ AB=4.3681P PB=8.36U AC=4.3681P PC=8.36U NE=8
Q$818 GND GND \$25 GND sky130_fd_pr__pnp_05v5_W0p68L0p68 AE=0.4624P PE=2.72U
+ AB=4.3681P PB=8.36U AC=4.3681P PC=8.36U NE=1
R$826 VDD VDD VDD 17264.1509434 sky130_fd_pr__res_iso_pw L=30U W=5.3U
R$827 \$10 \$174 VDD 23018.8679245 sky130_fd_pr__res_iso_pw L=60U W=7.95U
R$828 \$53 \$122 VDD 11509.4339623 sky130_fd_pr__res_iso_pw L=30U W=7.95U
R$837 GND GND GND 1620.94607173 sky130_fd_pr__res_xhigh_po_1p41
+ L=7.07137723794U W=8.725U
R$838 GND \$30 GND 100482.269504 sky130_fd_pr__res_xhigh_po_1p41 L=70.84U
+ W=1.41U
R$846 \$30 \$203 GND 28709.2198582 sky130_fd_pr__res_xhigh_po_1p41 L=20.24U
+ W=1.41U
R$853 \$25 GND GND 100482.269504 sky130_fd_pr__res_xhigh_po_1p41 L=70.84U
+ W=1.41U
R$865 \$16 VOP GND 6468.08510638 sky130_fd_pr__res_xhigh_po_1p41 L=4.56U W=1.41U
R$871 VOP vctrl GND 90553.1914894 sky130_fd_pr__res_xhigh_po_1p41 L=63.84U
+ W=1.41U
C$874 \$16 GND 4.97289984e-10 sky130_fd_pr__model__cap_mim A=248644.992P
+ P=35680U
C$1066 GND VOP 2.5120144e-11 sky130_fd_pr__model__cap_mim A=12560.072P P=2004.8U
C$1076 vn vp 3.64e-13 sky130_fd_pr__model__cap_mim A=182P P=54U
C$1151 vctrl GND 1.74227e-12 sky130_fd_pr__model__cap_mim A=871.135P P=118.06U
.ENDS integer_pll_2
