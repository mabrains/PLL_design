** Test bench for ring

.include ../spice_files/ring_cir.ckt


.lib /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice sf
.temp 27.00
.options tnom=27.00
VDD VDD GND 1.98

xring Vin Vout VDD GND ring

**** begin user architecture code

.control

    op 
    save all
        
    print all

    tran 2ns 4us uic
    plot Vout
    meas tran tperiod TRIG Vout VAL=0.4 RISE=15 TARG Vout VAL=0.4 RISE=16
    let freq = 1/(tperiod*1000000000)
    print freq
    
.endc

.GLOBAL GND
.GLOBAL VDD
.end