** Loop filter circuit model

.subckt loop_filter_3rd_order vout vctrl gnd
*old
    * C1 vout gnd 14.8p ic=0
    * R2 vout r2c2 18.5k
    * c2 r2c2 gnd 261.1p ic=0
    * R1 vout vctrl 163.85k
    * c3 vctrl gnd 1.332p ic=0
*calc

*NEW
    C1 vout gnd 25.5p ic=0
    R2 vout r2c2 6.6684k
    c2 r2c2 gnd 504p ic=0
    R1 vout vctrl 91.9513k
    c3 vctrl gnd 1.7642p ic=0
.ends

* .subckt loop_filter_3rd_order_ideal vout vctrl gnd
*     C1 vout gnd 66p ic=0
*     R2 vout r2c2 3.8k
*     c2 r2c2 gnd 1.32n ic=0
*     R1 vout vctrl 100k
*     c3 vctrl gnd 2.4p ic=0
* .ends
