* Circuit Model for  DIVIDER

*########################### 1/2 DIV behave ###############################

.subckt 1_2div Fin Fout Pa 0
+ TR=10e-15 TF=10e-15


	s1 Fin fin_int Pa 0 switch1 OFF
	.model switch1 sw vt=0.9 vh=0.01 ron=1 roff=1G
	Rout fin_int 0 10K

	are123 [fin_int] [fin_int_dig] adc_buff
	.model adc_buff adc_bridge(in_low = 0.9 in_high = 0.9)

	adivtest fin_int_dig fout_int_dig divider
	.model divider d_fdiv(div_factor = 2 high_cycles = 1
	+ i_count = 0 rise_delay = 8.5e-12
	+ fall_delay = 8.5e-12)

	abri2 [fout_int_dig] [fout1] dac1 
	.model dac1 dac_bridge(out_low = 0 out_high = 1.8 out_undef = 0.9
	+ input_load = 1e-15 t_rise = 1e-15
	+ t_fall = 1e-15)
	s12 fout1 Fout Pa 0 switch1 OFF

.ends 1_2DIV

.subckt buffer Fin Fout Pa 0
	s2 Fin Fout Pa 0 switch1 OFF
	Rout Fout 0 10K
	* s1 vout net1 cnt 0 switch1 OFF
	.model switch1 sw vt=0.9 vh=0.01 ron=1 roff=1G
.ends buffer


*########################### 1/2 DIV behave ###############################


.subckt 2to1_Cell Fin Fout Pa 0 MODIa MODO

	************************************************************
	*need to have pa and para first before

	are12c3 [Pa MODIa] [Pd MODId] adc_buff
	.model adc_buff adc_bridge(in_low = 0.9 in_high = 0.9)


	ainv1d Pd Pdbar invd1
	ainv1c MODId MODIdbar invd1	
	.model invd1 d_inverter(rise_delay = 1e-10 fall_delay = 1e-10)

	abri23 [Pdbar MODIdbar] [Para MODIabar] dac1 
	.model dac1 dac_bridge(out_low = 0 out_high = 1.8 out_undef = 0.9
	+ input_load = 1e-15 t_rise = 1e-15
	+ t_fall = 1e-15)

	Xbuffer Fin Fout Pa 0 buffer

	X1_2div1 Fin Fout Para 0 1_2div

	XMODO 0 MODO MODIabar 0 buffer
	X1_2div2 Fin MODO MODIa 0 1_2div



.ends 2to1_cell
