** sch_path: /home/tarek/Mabrains/Inv/New_crystal.sch
.subckt TOP VDD GND Cout Cin out
M11 Cout Cin VDD VDD sky130_fd_pr__pfet_01v8 L=0.15u W=240u nf=16 m=1
M2 Cout Cin GND GND sky130_fd_pr__nfet_01v8 L=0.15u W=240u nf=16 m=1
M1 out Cout VDD VDD sky130_fd_pr__pfet_01v8 L=0.15u W=15u nf=1 m=1
M3 out Cout GND GND sky130_fd_pr__nfet_01v8 L=0.15u W=15u nf=1 m=1
R1 Cin Cout GND sky130_fd_pr__res_xhigh_po_0p35 W=0.35u L=177.84u m=4
.ends
