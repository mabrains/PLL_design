** sch_path: /hoM_pfd_e/ahM_pfd_edelbadry/D_FF/conventional_pfd.sch

.subckt integer_pll VDD GND p0 p1 p2 p3 p4 p5 p6 p7 REF FB modi modo vco_out vp vn up dn VOP vctrl ibias_bgr ibias_vco ibias_cp    

*******************************pfd************************************
**********************************************************************        
**external nodes:up dn REF FB

M_pfd_1 pfd_net1 RST GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U nf=1 
M_pfd_2 pfd_net1 REF pfd_net2 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U nf=1 
M_pfd_3 pfd_net2 RST VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U nf=1
M_pfd_4 pfd_net3 pfd_net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U nf=1 
M_pfd_5 up_b pfd_net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U nf=1
M_pfd_6 up_b REF pfd_net3 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U nf=1  
M_pfd_7 up up_b GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U nf=1 
M_pfd_8 up up_b VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U nf=1 
M_pfd_9 pfd_net7 up_b VDD VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U nf=1 
M_pfd_10 RST dn_b pfd_net7 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U nf=1
M_pfd_11 dn dn_b GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U nf=1
M_pfd_12 dn dn_b VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U nf=1 
M_pfd_13 RST up_b GND GND sky130_fd_pr__nfet_01v8 L=0.2U W=2U nf=1
M_pfd_14 RST dn_b GND GND sky130_fd_pr__nfet_01v8 L=0.2U W=2U nf=1  
M_pfd_15 pfd_net6 pfd_net4 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U nf=1
M_pfd_16 dn_b pfd_net4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U nf=1 
M_pfd_17 pfd_net4 FB pfd_net5 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U nf=1 
M_pfd_18 dn_b FB pfd_net6 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U nf=1  
M_pfd_19 pfd_net5 RST VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U nf=1
M_pfd_20 pfd_net4 RST GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U nf=1 


*******************************cp*************************************
********************************************************************** 
**external nodes:up dn VOP  VBN

M_cp_p1 ibias_cp ibias_cp VDD VDD sky130_fd_pr__pfet_01v8 L=0.15u W=40u nf=4 m=1
M_cp_p2 VBN      ibias_cp VDD VDD sky130_fd_pr__pfet_01v8 L=0.15u W=10u nf=1 m=1


M_cp_1 cp_net1 Nbais GND GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U nf=1 m=2
M_cp_2 cp_net2 Nbais GND GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U nf=1 m=1
M_cp_3 VBp VBN cp_net1 GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U nf=1 m=2
M_cp_4 Nbais VBN cp_net2 GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U nf=1 m=1

R_cp1 VBN Nbais VDD sky130_fd_pr__res_iso_pw r=23.0188679245k   m=1 L=60u  W=7.95u
R_cp2 p_bais VBp VDD sky130_fd_pr__res_iso_pw r=11.5094339623k  m=1 L=30u  W=7.95u  
Rdumy VDD VDD VDD sky130_fd_pr__res_iso_pw r=17.2641509434k     m=1 L=30u  W=5.3u  

M_cp_5 p_bais VBp cp_net3 VDD sky130_fd_pr__pfet_01v8 L=0.6U W=6.66U nf=1 m=2
M_cp_6 cp_net3 p_bais VDD VDD sky130_fd_pr__pfet_01v8 L=0.6U W=6.66U nf=1 m=2

M_cp_7 cp_net4 Nbais GND GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U nf=1 m=10
M_cp_8 cp_net5 VBN cp_net4 GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U nf=1 m=10
M_cp_9 VON DNB cp_net5 GND sky130_fd_pr__nfet_01v8 L=0.15U W=4U nf=1 m=1
M_cp_10 VOP DN cp_net5 GND sky130_fd_pr__nfet_01v8 L=0.15U W=4U nf=1 m=1
M_cp_11 VOP UBP cp_net6 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=10U nf=1 m=1
M_cp_12 VON UP cp_net6 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=10U nf=1 m=1
M_cp_13 cp_net6 VBp cp_net7 VDD sky130_fd_pr__pfet_01v8 L=0.6U W=6.66U nf=1 m=10
M_cp_14 cp_net7 p_bais VDD VDD sky130_fd_pr__pfet_01v8 L=0.6U W=6.66U nf=1 m=10

M_cp_15 UBP UP GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_16 UBP UP VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=2U nf=1 m=1

M_cp_17 DNB DN GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_18 DNB DN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=2U nf=1 m=1

M_cp_19 cp_net2_ota Nbais GND GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U nf=1 m=2
M_cp_20 cp_net1_ota p_bais VDD VDD sky130_fd_pr__pfet_01v8 L=0.6U W=4U nf=1 m=2
M_cp_21 cp_net3_ota p_bais VDD VDD sky130_fd_pr__pfet_01v8 L=0.6U W=4U nf=1 m=2
M_cp_22 cp_net3_ota VON cp_net2_ota GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_23 cp_net1_ota VOP cp_net2_ota GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_24 cp_net5_ota cp_net4_ota GND GND sky130_fd_pr__nfet_01v8 L=1U W=1.3U nf=1 m=1
M_cp_25 GND cp_net4_ota GND GND sky130_fd_pr__nfet_01v8 L=1U W=1.3U nf=1 m=1
M_cp_26 cp_net4_ota VBN cp_net5_ota GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_27 VON VBN GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_28 VON VBp cp_net3_ota VDD sky130_fd_pr__pfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_29 cp_net4_ota VBp cp_net1_ota VDD sky130_fd_pr__pfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_30 cp_net6_ota p_bais VDD VDD sky130_fd_pr__pfet_01v8 L=0.6U W=6.66U nf=1 m=1
M_cp_32 GND VON cp_net6_ota VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_cp_33 cp_net5_ota VOP cp_net6_ota VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

*******************************lpf************************************
********************************************************************** 
**external nodes:VOP vctrl

C_lpf_1 VOP   gnd sky130_fd_pr__model__cap_mim W=25.06u L=25.06u MF=1 m=20   A=12.560072n    P=2.0048m 
c_lpf_2 r2c2  gnd sky130_fd_pr__model__cap_mim W=27.88u L=27.87u MF=1 m=320  A=0.248644992u    P=35.68m
c_lpf_3 vctrl gnd sky130_fd_pr__model__cap_mim W=29.5u  L=29.53u MF=1 m=1    A=0.871135n P=0.11806m

R_lpf_4     VOP r2c2   GND sky130_fd_pr__res_xhigh_po_1p41 L=4.56u  W=1.41u m=1
R_lpf_5     VOP vctrl  GND sky130_fd_pr__res_xhigh_po_1p41 L=63.84u W=1.41u m=1 
** R_lpf_dummy GND GND    GND sky130_fd_pr__res_xhigh_po_1p41 L=4.44u  W=2.82u m=1 $ this dummy res is compined with the dummy res of the bgr


*******************************bgr************************************
********************************************************************** 
**external nodes:ibias_bgr

Q_bgr_1 GND GND VBE GND sky130_fd_pr__pnp_05v5_W0p68L0p68 NE=1 m=1
Q_bgr_2 GND GND bgr_net2 GND sky130_fd_pr__pnp_05v5_W0p68L0p68 NE=8


R_bgr_4 bgr_net2 bgr_net3 GND sky130_fd_pr__res_xhigh_po_1p41 L=20.24u W=1.41u m=1
R_bgr_1 GND bgr_net3 GND sky130_fd_pr__res_xhigh_po_1p41 L=70.84u W=1.41u m=1
R_bgr_3 GND VBE GND sky130_fd_pr__res_xhigh_po_1p41 L=70.84u W=1.41u m=1

R_bgr_d1 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 L=7.07137723794u W=8.725u m=1 

M_bgr_15 bgr_net5 bgr_net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5u W=4u nf=4    
M_bgr_13 bgr_net3 bgr_net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5u W=20u nf=4    
M_bgr_14 VBE bgr_net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5u W=20u nf=4  
M_bgr_16 bgr_net1 bgr_net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5u W=44u nf=44
M_bgr_17 bgr_net6 bgr_net3 bgr_net5 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5u W=90u nf=6      
M_bgr_18 bgr_net4 VBE bgr_net5 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5u W=90u nf=6            
M_bgr_19 bgr_net1 bgr_net6 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5u W=0.42u m=10      
M_bgr_20 bgr_net6 bgr_net4 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5u W=0.42u m=4             
M_bgr_21 bgr_net4 bgr_net4 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5u W=0.42u m=4             
M_bgr_22 bgr_net7 bgr_net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1u W=40u nf=2     
M_bgr_23 bgr_net7 bgr_net1 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=20u W=0.42u         
M_bgr_24 VBE bgr_net7 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1u W=40u nf=2     
M_bgr_2 ibias_bgr bgr_net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5u W=200u nf=40 


*******************************cm*************************************
********************************************************************** 
**external nodes:ibias_vco ibias_cp

MBGR ibias_bgr ibias_bgr GND GND sky130_fd_pr__nfet_01v8 L=1u W=50u  nf=2  m=1
MVCO ibias_vco ibias_bgr GND GND sky130_fd_pr__nfet_01v8 L=1u W=250u nf=10 m=1
MCP  ibias_cp  ibias_bgr GND GND sky130_fd_pr__nfet_01v8 L=1u W=25u  nf=1  m=1



*******************************vco************************************
********************************************************************** 
**external nodes: vco_out

M_vco_4 vco_net2  ibias_vco VDD VDD sky130_fd_pr__pfet_01v8 L=0.5u W=1000u nf=50 m=1
M_vco_5 ibias_vco ibias_vco VDD VDD sky130_fd_pr__pfet_01v8 L=0.5u W=200u  nf=10 m=1

M_vco_11 vp vn vco_net2 vco_net2 sky130_fd_pr__pfet_01v8 L=0.15u W=250u nf=5 m=1
M_vco_1 vn vp vco_net2 vco_net2 sky130_fd_pr__pfet_01v8 L=0.15u W=250u  nf=5 m=1

M_vco_2 vp vn GND GND sky130_fd_pr__nfet_01v8 L=0.15u W=100u nf=5 m=1
M_vco_7 vn vp GND GND sky130_fd_pr__nfet_01v8 L=0.15u W=100u nf=5 m=1

M_vco_6 vctrl vn vctrl gnd sky130_fd_pr__nfet_01v8_lvt L=8u W=17u nf=1 m=1
M_vco_3 vctrl vp vctrl gnd sky130_fd_pr__nfet_01v8_lvt L=8u W=17u nf=1 m=1

C_load vp vn sky130_fd_pr__model__cap_mim W=14u L=13u MF=1 m=1 A=182p P=54u

*L1 vp vn 4.022n m=1

M_vco_inv_1 vco_out vp GND GND sky130_fd_pr__nfet_01v8 L=0.15u W=4.2u nf=1  m=1 
M_vco_inv_2 vco_out vp VDD VDD sky130_fd_pr__pfet_01v8 L=0.15u W=60u  nf=12 m=1

M_vco_inv_3 fout_dummy vn GND GND sky130_fd_pr__nfet_01v8 L=0.15u W=4.2u nf=1  m=1 
M_vco_inv_4 fout_dummy vn VDD VDD sky130_fd_pr__pfet_01v8 L=0.15u W=60u  nf=12 m=1

*******************************divider************************************
********************************************************************** 
**external nodes: p0 p1 p2 p3 p4 p5 p6 p7 vco_out FB

** divider  cdl


*FIRST CELL
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_2
M0 fout0 2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M1 fout0 1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M2 fout0 2 net1 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M3 net1 1 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M4 31 fout0 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M5 31 modi0 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M6 31 modi0 net2 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M7 net2 fout0 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M8 3 31 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M9 3 31 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M10 finb vco_out vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M11 finb vco_out gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M12 2 vco_out vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M13 2 p0 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M14 2 p0 net1_nand3 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M15 net1_nand3 vco_out net2_nand3 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M16 2 modo vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M17 net2_nand3 modo gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M18 net1_ff1 fout0 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M19 net3_ff1 finb net1_ff1 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M20 net3_ff1 vco_out net2_ff1 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M21 net2_ff1 fout0 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M22 net4_ff1 net3_ff1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M23 1 vco_out net4_ff1 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M24 1 finb net5_ff1 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M25 net5_ff1 net3_ff1 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M26 net1_ff2 3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M27 net3_ff2 finb net1_ff2 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M28 net3_ff2 vco_out net2_ff2 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M29 net2_ff2 3 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M30 net4_ff2 net3_ff2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M31 modo vco_out net4_ff2 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M32 modo finb net5_ff2 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M33 net5_ff2 net3_ff2 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1



*********************************///////////////SECOND CELL\\\\\\\\\\\\\*****************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_2
M100 fout1 201 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M101 fout1 101 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M102 fout1 201 net11 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M103 net11 101 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M104 3101 fout1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M105 3101 modi1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M106 3101 modi1 net201 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M107 net201 fout1 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M108 301 3101 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M109 301 3101 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M110 finb01 fout0 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M111 finb01 fout0 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M112 201 fout0 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M113 201 p1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M114 201 p1 net1_nand301 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M115 net1_nand301 fout0 net2_nand301 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M116 201 modi0 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M117 net2_nand301 modi0 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M118 net1_ff101 fout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M119 net3_ff101 finb01 net1_ff101 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M120 net3_ff101 fout0 net2_ff101 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M121 net2_ff101 fout1 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M122 net4_ff101 net3_ff101 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1	
M123 101 fout0 net4_ff101 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M124 101 finb01 net5_ff101 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M125 net5_ff101 net3_ff101 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M126 net1_ff201 301 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M127 net3_ff201 finb01 net1_ff201 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M128 net3_ff201 fout0 net2_ff201 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M129 net2_ff201 301 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M130 net4_ff201 net3_ff201 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M131 modi0 fout0 net4_ff201 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M132 modi0 finb01 net5_ff201 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M133 net5_ff201 net3_ff201 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1



*********************************///////////////THIRD CELL\\\\\\\\\\\\\*****************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_2
M200 fout2 202 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M201 fout2 102 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M202 fout2 202 net21 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M203 net21 102 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M204 3102 fout2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M205 3102 modi2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M206 3102 modi2 net202 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M207 net202 fout2 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M208 302 3102 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M209 302 3102 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M210 finb02 fout1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M211 finb02 fout1 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M212 202 fout1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M213 202 p2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M214 202 p2 net1_nand302 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M215 net1_nand302 fout1 net2_nand302 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M216 202 modi1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M217 net2_nand302 modi1 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M218 net1_ff102 fout2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M219 net3_ff102 finb02 net1_ff102 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M220 net3_ff102 fout1 net2_ff102 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M221 net2_ff102 fout2 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M222 net4_ff102 net3_ff102 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M223 102 fout1 net4_ff102 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M224 102 finb02 net5_ff102 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M225 net5_ff102 net3_ff102 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M226 net1_ff202 302 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M227 net3_ff202 finb02 net1_ff202 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M228 net3_ff202 fout1 net2_ff202 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M229 net2_ff202 302 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M230 net4_ff202 net3_ff202 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M231 modi1 fout1 net4_ff202 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M232 modi1 finb02 net5_ff202 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M233 net5_ff202 net3_ff202 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1



*********************************///////////////FOURTH CELL\\\\\\\\\\\\\*****************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************


** NAND_2
M300 fout3 203 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M301 fout3 103 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M302 fout3 203 net31 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M303 net31 103 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M304 3103 fout3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M305 3103 modi3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M306 3103 modi3 net203 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M307 net203 fout3 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M308 303 3103 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M309 303 3103 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M310 finb03 fout2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M311 finb03 fout2 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M312 203 fout2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M313 203 p3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M314 203 p3 net1_nand303 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M315 net1_nand303 fout2 net2_nand303 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M316 203 modi2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M317 net2_nand303 modi2 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M318 net1_ff103 fout3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M319 net3_ff103 finb03 net1_ff103 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M320 net3_ff103 fout2 net2_ff103 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M321 net2_ff103 fout3 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M322 net4_ff103 net3_ff103 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M323 103 fout2 net4_ff103 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M324 103 finb03 net5_ff103 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M325 net5_ff103 net3_ff103 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M326 net1_ff203 303 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M327 net3_ff203 finb03 net1_ff203 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M328 net3_ff203 fout2 net2_ff203 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M329 net2_ff203 303 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M330 net4_ff203 net3_ff203 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M331 modi2 fout2 net4_ff203 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M332 modi2 finb03 net5_ff203 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M333 net5_ff203 net3_ff203 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1


*********************************///////////////FIFTH CELL\\\\\\\\\\\\\*****************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_2
M400 fout4 204 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M401 fout4 104 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M402 fout4 204 net41 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M403 net41 104 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M404 3104 fout4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M405 3104 modi4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M406 3104 modi4 net204 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M407 net204 fout4 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M408 304 3104 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M409 304 3104 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M410 finb04 fout3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M411 finb04 fout3 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M412 204 fout3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M413 204 p4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M414 204 p4 net1_nand304 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M415 net1_nand304 fout3 net2_nand304 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M416 204 modi3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M417 net2_nand304 modi3 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M418 net1_ff104 fout4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M419 net3_ff104 finb04 net1_ff104 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M420 net3_ff104 fout3 net2_ff104 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M421 net2_ff104 fout4 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M422 net4_ff104 net3_ff104 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M423 104 fout3 net4_ff104 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M424 104 finb04 net5_ff104 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M425 net5_ff104 net3_ff104 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M426 net1_ff204 304 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M427 net3_ff204 finb04 net1_ff204 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M428 net3_ff204 fout3 net2_ff204 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M429 net2_ff204 304 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M430 net4_ff204 net3_ff204 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M431 modi3 fout3 net4_ff204 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M432 modi3 finb04 net5_ff204 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M433 net5_ff204 net3_ff204 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*********************************///////////////SIXTHS CELL\\\\\\\\\\\\\*****************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_2
M500 fout5 205 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M501 fout5 105 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M502 fout5 205 net51 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M503 net51 105 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M504 3105 fout5 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M505 3105 modi5 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M506 3105 modi5 net205 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M507 net205 fout5 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M508 305 3105 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M509 305 3105 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M510 finb05 fout4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M511 finb05 fout4 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M512 205 fout4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M513 205 p5 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M514 205 p5 net1_nand305 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M515 net1_nand305 fout4 net2_nand305 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M516 205 modi4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M517 net2_nand305 modi4 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M518 net1_ff105 fout5 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M519 net3_ff105 finb05 net1_ff105 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M520 net3_ff105 fout4 net2_ff105 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M521 net2_ff105 fout5 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M522 net4_ff105 net3_ff105 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M523 105 fout4 net4_ff105 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M524 105 finb05 net5_ff105 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M525 net5_ff105 net3_ff105 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M526 net1_ff205 305 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M527 net3_ff205 finb05 net1_ff205 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M528 net3_ff205 fout4 net2_ff205 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M529 net2_ff205 305 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M530 net4_ff205 net3_ff205 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M531 modi4 fout4 net4_ff205 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M532 modi4 finb05 net5_ff205 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M533 net5_ff205 net3_ff205 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*********************************///////////////SEVENTH CELL\\\\\\\\\\\\\*****************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_2
M600 fout6 206 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M601 fout6 106 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M602 fout6 206 net61 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M603 net61 106 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M604 3106 fout6 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M605 3106 modi6 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M606 3106 modi6 net206 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M607 net206 fout6 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M608 306 3106 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M609 306 3106 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M610 finb06 fout5 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M611 finb06 fout5 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M612 206 fout5 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M613 206 p6 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M614 206 p6 net1_nand306 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M615 net1_nand306 fout5 net2_nand306 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M616 206 modi5 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M617 net2_nand306 modi5 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M618 net1_ff106 fout6 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M619 net3_ff106 finb06 net1_ff106 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M620 net3_ff106 fout5 net2_ff106 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M621 net2_ff106 fout6 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M622 net4_ff106 net3_ff106 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M623 106 fout5 net4_ff106 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M624 106 finb06 net5_ff106 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M625 net5_ff106 net3_ff106 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M626 net1_ff206 306 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M627 net3_ff206 finb06 net1_ff206 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M628 net3_ff206 fout5 net2_ff206 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M629 net2_ff206 306 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M630 net4_ff206 net3_ff206 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M631 modi5 fout5 net4_ff206 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M632 modi5 finb06 net5_ff206 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M633 net5_ff206 net3_ff206 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1



*********************************///////////////EIGHTS CELL\\\\\\\\\\\\\*****************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_2
M700 FB 207 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M701 FB 107 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M702 FB 207 net71 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M703 net71 107 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M704 3107 FB vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M705 3107 modi vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M706 3107 modi net207 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M707 net207 FB gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M708 307 3107 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M709 307 3107 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M710 finb07 fout6 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M711 finb07 fout6 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M712 207 fout6 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M713 207 p7 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M714 207 p7 net1_nand307 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M715 net1_nand307 fout6 net2_nand307 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M716 207 modi6 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M717 net2_nand307 modi6 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M718 net1_ff107 FB VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M719 net3_ff107 finb07 net1_ff107 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M720 net3_ff107 fout6 net2_ff107 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M721 net2_ff107 FB GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M722 net4_ff107 net3_ff107 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M723 107 fout6 net4_ff107 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M724 107 finb07 net5_ff107 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M725 net5_ff107 net3_ff107 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M726 net1_ff207 307 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M727 net3_ff207 finb07 net1_ff207 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M728 net3_ff207 fout6 net2_ff207 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M729 net2_ff207 307 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M730 net4_ff207 net3_ff207 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M731 modi6 fout6 net4_ff207 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M732 modi6 finb07 net5_ff207 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M733 net5_ff207 net3_ff207 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1


.ends
