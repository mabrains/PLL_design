* Circuit Model for PFD


.subckt PFD REF FB UP DWN FBS REFS
+ CLKDelay=1.0e-10 SetDelay=1.0e-10 ResetDelay=1.0e-10 
+ Out_initial_state=2 TR=1.0e-10 TF=1.0e-10 + Cand=1e-12

	* Analog to Digital nodes Models
	.model adc_buff adc_bridge(in_low = 0.9 in_high = 0.9)

	* Digital REF
	aref [REF] [REF_D] adc_buff

	* Digital FB
	afb [FB] [FB_D] adc_buff

	*Define the and gate
	a_andGate [UP_Signal DW_Signal] RESET and1

	.model and1 d_and(rise_delay = TR fall_delay = TF
	+ input_load = Cand )

	*Define the flip flops
	a_ff1 d_d1 REF_D d_d0 RESET UP_Signal UP_Signal_bar flop1

	a_ff2 d_d1 FB_D d_d0 RESET DW_Signal DWN_Signal_bar flop1

	.model flop1 d_dff(clk_delay = {CLKDelay} set_delay = {SetDelay}
	+ reset_delay = {ResetDelay} ic = {Out_initial_state} rise_delay = {TR}
	+ fall_delay = {TF})

	* Digital to Analog nodes Models
	abridge-w1 [FB_D REF_D UP_Signal DW_Signal UP_Signal_bar DWN_Signal_bar] [FBS REFS UP DWN UP_bar DWN_bar] dac1 

	.model dac1 dac_bridge(out_low = 0 out_high = 1.8 out_undef = 0.9
	+ input_load = 1e-15 t_rise = 1e-15
	+ t_fall = 1e-15)

.ends PFD
