** pex of divider