
.include divider_cell.ckt

.subckt divider  vdd fout gnd p2 p7 p1 p6 p5 p4 p3 p0 fin float
x1 vdd net1 fin p0 float gnd net2 divider_cell
x2 vdd net3 net1 p1 net2 gnd net4 divider_cell
x3 vdd net5 net3 p2 net4 gnd net6 divider_cell
x4 vdd net7 net5 p3 net6 gnd net8 divider_cell
x5 vdd net9 net7 p4 net8 gnd net10 divider_cell
x6 vdd net11 net9 p5 net10 gnd net12 divider_cell
x7 vdd net13 net11 p6 net12 gnd net14 divider_cell
x8 vdd fout net13 p7 net14 gnd vdd divider_cell
.ends

.GLOBAL VDD
.GLOBAL GND
