* bgr behav

.subckt bgr_behav VDD ibias
Isource VDD ibias 90u        
.ends
