* SDM behav subcircuit
***************************************** 1-BIT--ADDER **********************************
.subckt ADDER A B CIN S1 COUT1

+TR=1.0e-10 TF=1.0e-10 + Cand=1e-12

    * S    = ( A XOR B ) XOR Cin
    * Cout = A and B or  Cin and (A XOR B)

    *Define the and gate

    * AndB = A and B
	a_andGate [A B] AandB and1

    * Cin and (A XOR B)
    a_andGate2 [Cin AxorB] Cinand_AxorB and1

	.model and1 d_and(rise_delay = TR fall_delay = TF
	+ input_load = Cand )

    *Define the or gate

    a_orGate [AandB Cinand_AxorB] COUT1 or1

    .model or1 d_or(rise_delay = TR fall_delay = TF
	+ input_load = Cand )

    *Define the xor gate
    
    a_xorGate [A B] AxorB xor3
    a_xorGate2 [AxorB CIN] S1 xor3

    .model xor3 d_xor(rise_delay = TR fall_delay = TF
	+ input_load = Cand )

.ends ADDER

***************************************** 1-BIT--ADDER **********************************

*########################################################################################

***************************************** 5-BIT--ADDER **********************************

.subckt 5Bit_ADDER A0 A1 A2 A3 A4 B0 B1 B2 B3 B4 S0 S1 S2 S3 S4 COUT

	* A[5], B[5]  S[5]  , C[1] 

	XFA1 A0 B0 d_d0 S0 C1 ADDER
	XFA2 A1 B1 C1 S1 C2 ADDER
	XFA3 A2 B2 C2 S2 C3 ADDER
	XFA4 A3 B3 C3 S3 C4 ADDER
	XFA5 A4 B4 C4 S4 COUT ADDER

.ends 7Bit_ADDER

***************************************** 5-BIT--ADDER **********************************

*########################################################################################

****************************************** 7-BIT--ADDER **********************************

.subckt 7Bit_ADDER A0 A1 A2 A3 A4 A5 A6 B0 B1 B2 B3 B4 B5 B6 S0 S1 S2 S3 S4 S5 S6 COUT

	* A[7], B[7]  S[7]  , C[1] 

	XFA1 A0 B0 d_d0 S0 C1 ADDER
	XFA2 A1 B1 C1 S1 C2 ADDER
	XFA3 A2 B2 C2 S2 C3 ADDER
	XFA4 A3 B3 C3 S3 C4 ADDER
	XFA5 A4 B4 C4 S4 C5 ADDER
	XFA6 A5 B5 C5 S5 C6 ADDER
	XFA7 A6 B6 C6 S6 COUT ADDER

.ends 7Bit_ADDER

***************************************** 7-BIT--ADDER **********************************

*########################################################################################

 ************************************** 5-BIT--SUBTRACTOR ********************************

.subckt 5Bit_SUBTRACTOR A0 A1 A2 A3 A4 B0 B1 B2 B3 B4 S0 S1 S2 S3 S4 COUT

    * Set Cin = 1 and get the two complemnt

	ab0 B0 BI0 invd1
	ab1 B1 BI1 invd1
	ab2 B2 BI2 invd1
	ab3 B3 BI3 invd1
	ab4 B4 BI4 invd1

	.model invd1 d_inverter(rise_delay = 1e-10 fall_delay = 1e-10)

	* A[7], B[7]  S[7]  , C[1] 
	XFA1 A0 BI0 d_d1 S0 C1 ADDER
	XFA2 A1 BI1 C1 S1 C2 ADDER
	XFA3 A2 BI2 C2 S2 C3 ADDER
	XFA4 A3 BI3 C3 S3 C4 ADDER
	XFA5 A4 BI4 C4 S4 C5 ADDER

.ends 5Bit_SUBTRACTOR

 ************************************** 5-BIT--SUBTRACTOR ********************************

*########################################################################################

***************************************** SUMMER ************************************

.subckt SUMMER A0 A1 A2 A3 A4 B0 B1 B2 B3 B4 INV0 INV1 INV2 INV3 INV4 O0 O1 O2 O3 O4

    *[ 0 0 0 0 c1 ] ,[ 0 0 0 0 c2] , 2's compl[c3] , OUTPUT [5]

	X5Bit_ADDER A0 A1 A2 A3 A4 B0 B1 B2 B3 B4 S0 S1 S2 S3 S4 COUT1 5Bit_ADDER
	X5Bit_SUBTRACTOR S0 S1 S2 S3 S4 INV0 INV1 INV2 INV3 INV4 O0 O1 O2 O3 O4 COUT2 5Bit_SUBTRACTOR

.ends SUMMER

***************************************** SUMMER ************************************

*########################################################################################

***************************************** 5-BIT--REG ************************************

.subckt 5Bit_Register D1 D2 D3 D4 D5 CLK SET RESET OUT1 OUT2 OUT3 OUT4 OUT5

+ CLKDelay=1.0e-10 SetDelay=1.0e-10 ResetDelay=1.0e-10 
+ Out_initial_state=0 TR=1.0e-10 TF=1.0e-10 + Cand=1e-12

	*Define the flip flops

	a_ff1 D1 CLK SET RESET OUT1 OUT_BAR1 flop1
	a_ff2 D2 CLK SET RESET OUT2 OUT_BAR2 flop1
	a_ff3 D3 CLK SET RESET OUT3 OUT_BAR3 flop1
	a_ff4 D4 CLK SET RESET OUT4 OUT_BAR4 flop1
	a_ff5 D5 CLK SET RESET OUT5 OUT_BAR5 flop1

	.model flop1 d_dff(clk_delay = {CLKDelay} set_delay = {SetDelay}
	+ reset_delay = {ResetDelay} ic = {Out_initial_state} rise_delay = {TR}
	+ fall_delay = {TF}) 

.ends 5Bit_Register

***************************************** 5-BIT--REG ************************************

*########################################################################################

***************************************** 7-BIT--REG ************************************

.subckt 7Bit_Register D1 D2 D3 D4 D5 D6 D7 CLK SET RESET OUT1 OUT2 OUT3 OUT4 OUT5 OUT6 OUT7

+ CLKDelay=1.0e-10 SetDelay=1.0e-10 ResetDelay=1.0e-10 
+ Out_initial_state=0 TR=1.0e-10 TF=1.0e-10 + Cand=1e-12

	*Define the flip flops

	a_ff1 D1 CLK SET RESET OUT1 OUT_BAR1 flop1
	a_ff2 D2 CLK SET RESET OUT2 OUT_BAR2 flop1
	a_ff3 D3 CLK SET RESET OUT3 OUT_BAR3 flop1
	a_ff4 D4 CLK SET RESET OUT4 OUT_BAR4 flop1
	a_ff5 D5 CLK SET RESET OUT5 OUT_BAR5 flop1
	a_ff6 D6 CLK SET RESET OUT6 OUT_BAR6 flop1
	a_ff7 D7 CLK SET RESET OUT7 OUT_BAR7 flop1

	.model flop1 d_dff(clk_delay = {CLKDelay} set_delay = {SetDelay}
	+ reset_delay = {ResetDelay} ic = {Out_initial_state} rise_delay = {TR}
	+ fall_delay = {TF}) 

.ends 7Bit_Register

***************************************** 7-BIT--REG ************************************

*########################################################################################

***************************************** Acuumulator ************************************

.subckt Accumulator A0 A1 A2 A3 A4 A5 A6 RESET CLK CO B0 B1 B2 B3 B4 B5 B6

    X7Bit_ADDER A0 A1 A2 A3 A4 A5 A6 B0 B1 B2 B3 B4 B5 B6 S0 S1 S2 S3 S4 S5 S6 CO 7Bit_ADDER

    X7Bit_Register S0 S1 S2 S3 S4 S5 S6 CLK d_d0 RESET B0 B1 B2 B3 B4 B5 B6 7Bit_Register

.ends Accumulator

***************************************** Acuumulator ************************************

*########################################################################################

*****************************************--SDM--*****************************************

.subckt SDM A0 A1 A2 A3 A4 A5 A6 RESET CLK DIV0 DIV1 DIV2 DIV3 DIV4
    XAccumulator1 A0 A1 A2 A3 A4 A5 A6 RESET CLK_D C1 B0 B1 B2 B3 B4 B5 B6 Accumulator
    XAccumulator2 B0 B1 B2 B3 B4 B5 B6 RESET CLK_D C2 BB0 BB1 BB2 BB3 BB4 BB5 BB6 Accumulator
    XAccumulator3 BB0 BB1 BB2 BB3 BB4 BB5 BB6 RESET CLK_D C3 BBB0 BBB1 BBB2 BBB3 BBB4 BBB5 BBB6 Accumulator
    X5Bit_Register1 C3 d_d0 d_d0 d_d0 d_d0 CLK_D d_d0 d_d0 OUT1 OUT2 OUT3 OUT4 OUT5 5Bit_Register
    XSUMMER1 C2 d_d0 d_d0 d_d0 d_d0 C3 d_d0 d_d0 d_d0 d_d0 OUT1 OUT2 OUT3 OUT4 OUT5 O0 O1 O2 O3 O4 SUMMER
    X5Bit_Register2 OUT1 OUT2 OUT3 OUT4 OUT5 CLK_D d_d0 d_d0 K0 K1 K2 K3 K4 5Bit_Register
    XSUMMER2 C1 d_d0 d_d0 d_d0 d_d0 OUT1 OUT2 OUT3 OUT4 OUT5 K0 K1 K2 K3 K4 DIV0 DIV1 DIV2 DIV3 DIV4 SUMMER
.ends SDM

*****************************************--SDM--*****************************************

*########################################################################################
