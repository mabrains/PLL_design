* Extracted by KLayout with SKY130 LVS runset on : 16/11/2022 12:33

.SUBCKT integer_pll VDD dn ibias_bgr ibias_cp up ibias_vco vn VOP vctrl vp
+ vco_out FB modi P7 P6 P5 P4 modo P0 P1 P2 P3 REF GND
M$1 VDD dn \$3 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$2 \$14 \$52 \$18 VDD sky130_fd_pr__pfet_01v8 L=0.6U W=66.6U AS=19.314P
+ AD=19.314P PS=139U PD=139U
M$5 \$8 \$52 \$121 VDD sky130_fd_pr__pfet_01v8 L=0.6U W=13.32U AS=3.8628P
+ AD=3.8628P PS=27.8U PD=27.8U
M$14 GND \$10 \$280 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$15 \$106 VOP \$280 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$16 ibias_cp ibias_cp VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=40U AS=9.5P
+ AD=9.5P PS=61.9U PD=61.9U
M$18 VDD ibias_cp \$174 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=10U AS=2.9P
+ AD=2.9P PS=20.58U PD=20.58U
M$21 \$10 up \$18 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=10U AS=2.9P AD=2.9P
+ PS=20.58U PD=20.58U
M$22 VOP \$309 \$18 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=10U AS=2.9P AD=2.9P
+ PS=20.58U PD=20.58U
M$23 \$95 \$52 \$282 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=1U AS=0.29P AD=0.29P
+ PS=2.58U PD=2.58U
M$24 \$10 \$52 \$284 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=1U AS=0.29P AD=0.29P
+ PS=2.58U PD=2.58U
M$25 VDD \$121 \$14 VDD sky130_fd_pr__pfet_01v8 L=0.6U W=66.6U AS=19.314P
+ AD=19.314P PS=139U PD=139U
M$28 VDD \$121 \$8 VDD sky130_fd_pr__pfet_01v8 L=0.6U W=13.32U AS=3.8628P
+ AD=3.8628P PS=27.8U PD=27.8U
M$31 VDD \$121 \$280 VDD sky130_fd_pr__pfet_01v8 L=0.6U W=6.66U AS=1.9314P
+ AD=1.9314P PS=13.9U PD=13.9U
M$38 \$282 \$121 VDD VDD sky130_fd_pr__pfet_01v8 L=0.6U W=8U AS=2.32P AD=2.32P
+ PS=17.16U PD=17.16U
M$39 \$284 \$121 VDD VDD sky130_fd_pr__pfet_01v8 L=0.6U W=8U AS=2.32P AD=2.32P
+ PS=17.16U PD=17.16U
M$42 \$330 vn VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=60U AS=10.625P
+ AD=10.625P PS=69.25U PD=69.25U
M$54 vco_out vp VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=60U AS=10.625P
+ AD=10.625P PS=69.25U PD=69.25U
M$66 VDD up \$309 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$67 vn vp \$472 \$472 sky130_fd_pr__pfet_01v8 L=0.15U W=250U AS=48.5P
+ AD=41.25P PS=301.94U PD=251.65U
M$68 \$472 vn vp \$472 sky130_fd_pr__pfet_01v8 L=0.15U W=250U AS=41.25P
+ AD=48.5P PS=251.65U PD=301.94U
M$77 \$501 \$444 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$78 \$502 \$455 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$79 \$349 \$444 \$525 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$80 \$525 \$352 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$81 \$352 \$501 \$528 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$82 \$528 \$428 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$83 \$355 \$444 \$531 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$84 \$531 \$359 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$85 \$359 \$501 \$534 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$86 \$534 \$384 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$87 \$503 \$467 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$88 \$368 \$384 \$566 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$89 \$566 \$371 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$90 \$371 \$500 \$515 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$91 \$515 \$413 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$92 \$373 \$384 \$567 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$93 \$567 \$419 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$94 \$419 \$500 \$520 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$95 \$520 FB VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$96 \$500 \$384 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$97 \$387 \$455 \$570 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$98 \$570 \$389 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$99 \$389 \$502 \$543 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$100 \$543 \$434 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$101 \$392 \$455 \$546 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$102 \$546 \$396 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$103 \$396 \$502 \$549 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$104 \$549 \$444 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$105 \$401 \$467 \$573 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$106 \$573 \$451 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$107 \$451 \$503 \$574 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$108 \$574 \$447 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$109 \$405 \$467 \$558 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$110 \$558 \$410 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$111 \$410 \$503 \$561 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$112 \$561 \$455 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$113 \$472 ibias_vco VDD VDD sky130_fd_pr__pfet_01v8 L=0.5U W=1000U AS=147.9P
+ AD=147.9P PS=1034.79U PD=1034.79U
M$122 VDD ibias_vco ibias_vco VDD sky130_fd_pr__pfet_01v8 L=0.5U W=200U AS=29P
+ AD=29P PS=202.9U PD=202.9U
M$173 \$413 \$417 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$174 VDD FB \$417 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$175 VDD modi \$417 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$176 VDD \$373 FB VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$177 VDD \$427 FB VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$178 VDD \$368 \$427 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$179 VDD \$384 \$427 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$180 VDD P7 \$427 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$181 \$428 \$380 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$182 VDD \$384 \$380 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$183 VDD \$368 \$380 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$184 VDD \$355 \$384 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$185 VDD \$385 \$384 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$186 VDD \$349 \$385 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$187 VDD \$444 \$385 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$188 VDD P6 \$385 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$189 \$434 \$438 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$190 VDD \$444 \$438 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$191 VDD \$349 \$438 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$192 VDD \$392 \$444 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$193 VDD \$399 \$444 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$194 VDD \$387 \$399 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$195 VDD \$455 \$399 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$196 VDD P5 \$399 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$197 \$447 \$450 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$198 VDD \$455 \$450 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$199 VDD \$387 \$450 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$200 VDD \$405 \$455 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$201 VDD \$458 \$455 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$202 VDD \$401 \$458 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$203 VDD \$467 \$458 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$204 VDD P4 \$458 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$205 VDD \$874 \$871 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U AS=1.45P
+ AD=1.45P PS=10.58U PD=10.58U
M$206 \$871 REF \$859 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$207 VDD \$859 \$872 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U AS=1.45P
+ AD=1.45P PS=10.58U PD=10.58U
M$208 \$860 REF \$872 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$209 VDD \$872 \$873 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U AS=1.16P AD=0.58P
+ PS=8.58U PD=4.29U
M$210 \$873 \$875 \$874 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U AS=0.58P
+ AD=1.16P PS=4.29U PD=8.58U
M$211 VDD \$872 up VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U AS=1.45P AD=1.45P
+ PS=10.58U PD=10.58U
M$212 dn \$875 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U AS=1.45P AD=1.45P
+ PS=10.58U PD=10.58U
M$213 \$875 FB \$861 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$214 \$875 \$862 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U AS=1.45P
+ AD=1.45P PS=10.58U PD=10.58U
M$215 \$862 FB \$876 VDD sky130_fd_pr__pfet_01v8 L=0.2U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$216 \$876 \$874 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=5U AS=1.45P
+ AD=1.45P PS=10.58U PD=10.58U
M$217 \$611 P0 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$218 \$611 vco_out VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$219 \$611 modo VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$220 \$739 \$611 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$221 \$739 \$622 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$222 VDD vco_out \$614 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$223 VDD \$739 \$616 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$224 \$616 \$614 \$618 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$225 VDD \$618 \$620 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$226 \$620 vco_out \$622 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$227 VDD \$634 \$624 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$228 \$624 \$614 \$626 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$229 VDD \$626 \$628 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$230 \$628 vco_out modo VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$231 \$632 \$649 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$232 \$632 \$739 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$233 VDD \$632 \$634 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$234 \$635 P1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$235 \$635 \$739 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$236 \$635 \$649 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$237 \$740 \$635 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$238 \$740 \$698 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$239 VDD \$739 \$696 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$240 VDD \$740 \$697 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$241 \$697 \$696 \$640 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$242 VDD \$640 \$642 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$243 \$642 \$739 \$698 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$244 VDD \$653 \$645 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$245 \$645 \$696 \$699 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$246 VDD \$699 \$700 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$247 \$700 \$739 \$649 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$248 \$651 \$670 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$249 \$651 \$740 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$250 VDD \$651 \$653 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$251 \$654 P2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$252 \$654 \$740 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$253 \$654 \$670 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$254 \$741 \$654 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$255 \$741 \$664 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$256 VDD \$740 \$657 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$257 VDD \$741 \$701 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$258 \$701 \$657 \$660 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$259 VDD \$660 \$662 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$260 \$662 \$740 \$664 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$261 VDD \$674 \$702 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$262 \$702 \$657 \$703 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$263 VDD \$703 \$668 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$264 \$668 \$740 \$670 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$265 \$672 \$691 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$266 \$672 \$741 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$267 VDD \$672 \$674 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$268 \$675 P3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$269 \$675 \$741 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$270 \$675 \$691 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$271 \$467 \$675 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$272 \$467 \$684 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$273 VDD \$741 \$704 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$274 VDD \$467 \$679 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$275 \$679 \$704 \$681 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$276 VDD \$681 \$705 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$277 \$705 \$741 \$684 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$278 VDD \$695 \$686 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$279 \$686 \$704 \$706 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$280 VDD \$706 \$689 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$281 \$689 \$741 \$691 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$282 \$693 \$401 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$283 \$693 \$467 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$284 VDD \$693 \$695 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$285 VDD \$17 ibias_bgr VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5U W=200U
+ AS=30.74P AD=30.74P PS=273.48U PD=273.48U
M$317 VDD \$17 \$17 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5U W=44U AS=6.38P
+ AD=6.38P PS=56.76U PD=56.76U
M$357 \$30 \$17 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1U W=40U AS=8.7P AD=8.7P
+ PS=60.87U PD=60.87U
M$359 \$24 \$30 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1U W=40U AS=8.7P AD=8.7P
+ PS=60.87U PD=60.87U
M$361 \$35 \$29 \$33 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5U W=90U AS=15.225P
+ AD=15.225P PS=107.03U PD=107.03U
M$362 \$33 \$24 \$36 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5U W=90U AS=13.05P
+ AD=13.05P PS=91.74U PD=91.74U
M$381 VDD \$17 \$29 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5U W=20U AS=2.9P
+ AD=2.9P PS=25.8U PD=25.8U
M$383 VDD \$17 \$24 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5U W=20U AS=2.9P
+ AD=2.9P PS=25.8U PD=25.8U
M$437 VDD \$17 \$33 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5U W=4U AS=0.58P
+ AD=0.58P PS=5.16U PD=5.16U
M$589 GND dn \$3 GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U AS=0.29P AD=0.29P
+ PS=2.58U PD=2.58U
M$590 \$258 dn VOP GND sky130_fd_pr__nfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$591 \$258 \$3 \$10 GND sky130_fd_pr__nfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$592 GND \$9 \$56 GND sky130_fd_pr__nfet_01v8 L=0.6U W=20U AS=5.8P AD=5.8P
+ PS=45.8U PD=45.8U
M$594 GND \$9 \$57 GND sky130_fd_pr__nfet_01v8 L=0.6U W=4U AS=1.16P AD=1.16P
+ PS=9.16U PD=9.16U
M$596 GND \$9 \$58 GND sky130_fd_pr__nfet_01v8 L=0.6U W=4U AS=1.16P AD=1.16P
+ PS=9.16U PD=9.16U
M$599 GND \$9 \$59 GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$607 \$106 \$95 GND GND sky130_fd_pr__nfet_01v8 L=1U W=1.3U AS=0.377P
+ AD=0.377P PS=3.18U PD=3.18U
M$608 \$95 \$174 \$106 GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U AS=0.29P
+ AD=0.29P PS=2.58U PD=2.58U
M$609 GND \$95 GND GND sky130_fd_pr__nfet_01v8 L=1U W=1.3U AS=0.377P AD=0.377P
+ PS=3.18U PD=3.18U
M$610 \$10 \$174 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U AS=0.29P AD=0.29P
+ PS=2.58U PD=2.58U
M$611 \$56 \$174 \$258 GND sky130_fd_pr__nfet_01v8 L=0.6U W=20U AS=5.8P AD=5.8P
+ PS=45.8U PD=45.8U
M$614 \$58 \$174 \$52 GND sky130_fd_pr__nfet_01v8 L=0.6U W=4U AS=1.16P AD=1.16P
+ PS=9.16U PD=9.16U
M$617 \$59 \$174 \$9 GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$624 \$284 \$10 \$57 GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U AS=0.29P
+ AD=0.29P PS=2.58U PD=2.58U
M$625 \$282 VOP \$57 GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U AS=0.29P AD=0.29P
+ PS=2.58U PD=2.58U
M$626 vn vp GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=100U AS=19.4P AD=16.5P
+ PS=121.94U PD=101.65U
M$627 GND vn vp GND sky130_fd_pr__nfet_01v8 L=0.15U W=100U AS=16.5P AD=19.4P
+ PS=101.65U PD=121.94U
M$636 ibias_vco ibias_bgr GND GND sky130_fd_pr__nfet_01v8 L=1U W=250U
+ AS=39.875P AD=39.875P PS=278.19U PD=278.19U
M$641 GND ibias_bgr ibias_bgr GND sky130_fd_pr__nfet_01v8 L=1U W=50U AS=7.25P
+ AD=7.25P PS=50.58U PD=50.58U
M$648 ibias_cp ibias_bgr GND GND sky130_fd_pr__nfet_01v8 L=1U W=25U AS=7.25P
+ AD=7.25P PS=50.58U PD=50.58U
M$649 GND up \$309 GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U AS=0.29P AD=0.29P
+ PS=2.58U PD=2.58U
M$650 vco_out vp GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=4.2U AS=1.218P
+ AD=1.218P PS=8.98U PD=8.98U
M$651 \$330 vn GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=4.2U AS=1.218P
+ AD=1.218P PS=8.98U PD=8.98U
M$652 \$348 \$413 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$653 \$349 \$501 \$430 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$654 \$430 \$352 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$655 \$352 \$444 \$354 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$656 \$354 \$428 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$657 \$355 \$501 \$357 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$658 \$357 \$359 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$659 \$359 \$444 \$431 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$660 \$431 \$384 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$661 \$387 \$502 \$439 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$662 \$439 \$389 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$663 \$389 \$455 \$440 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$664 \$440 \$434 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$665 \$392 \$502 \$393 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$666 \$393 \$396 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$667 \$396 \$455 \$441 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$668 \$441 \$444 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$669 \$363 \$447 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$670 \$368 \$500 \$369 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$671 \$369 \$371 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$672 \$371 \$384 \$348 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$673 \$373 \$500 \$418 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$674 \$418 \$419 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$675 \$419 \$384 \$420 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$676 \$420 FB GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$677 GND \$444 \$501 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$678 GND \$349 \$432 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$679 \$432 \$444 \$433 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$680 \$433 P6 \$385 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$681 GND \$455 \$502 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$682 \$401 \$503 \$362 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$683 \$362 \$451 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$684 \$451 \$467 \$363 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$685 \$405 \$503 \$407 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$686 \$407 \$410 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$687 \$410 \$467 \$411 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$688 \$411 \$455 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$689 GND \$467 \$503 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$690 \$611 P0 \$766 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$691 GND \$417 \$413 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$692 \$766 vco_out \$767 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$693 GND FB \$415 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$694 \$767 modo GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$695 \$415 modi \$417 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$696 \$739 \$611 \$746 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$697 \$746 \$622 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$698 GND \$384 \$500 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$699 GND \$373 \$422 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$700 \$422 \$427 FB GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$701 \$632 \$649 \$768 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$702 GND \$368 \$425 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$703 \$768 \$739 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$704 \$425 \$384 \$426 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$705 \$426 P7 \$427 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$706 GND \$380 \$428 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$707 GND \$384 \$429 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$708 \$429 \$368 \$380 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$709 \$740 \$635 \$771 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$710 \$771 \$698 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$711 GND \$355 \$382 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$712 \$382 \$385 \$384 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$713 \$651 \$670 \$753 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$714 \$753 \$740 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$715 GND \$438 \$434 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$716 GND \$444 \$436 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$717 \$436 \$349 \$438 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$718 GND \$392 \$398 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$719 \$398 \$399 \$444 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$720 GND \$387 \$445 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$721 \$445 \$455 \$446 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$722 \$446 P5 \$399 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$723 GND \$450 \$447 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$724 GND \$455 \$400 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$725 \$400 \$387 \$450 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$726 GND \$405 \$453 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$727 \$453 \$458 \$455 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$728 GND \$401 \$456 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$729 \$456 \$467 \$457 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$730 \$457 P4 \$458 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$731 \$635 P1 \$769 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$732 \$769 \$739 \$770 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$733 \$770 \$649 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$734 \$741 \$654 \$756 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$735 \$756 \$664 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$736 \$672 \$691 \$774 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$737 \$774 \$741 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$738 \$467 \$675 \$761 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$739 \$761 \$684 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$740 \$693 \$401 \$764 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$741 \$764 \$467 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$742 \$614 vco_out GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$743 GND \$739 \$778 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$744 \$778 vco_out \$618 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$745 GND \$618 \$781 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$746 \$781 \$614 \$622 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$747 \$783 vco_out \$626 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$748 GND \$626 \$786 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$749 \$786 \$614 modo GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$750 \$634 \$632 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$751 \$696 \$739 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$752 GND \$740 \$789 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$753 \$789 \$739 \$640 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$754 GND \$640 \$792 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$755 \$792 \$696 \$698 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$756 \$794 \$739 \$699 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$757 GND \$699 \$797 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$758 \$797 \$696 \$649 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$759 \$653 \$651 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$760 \$654 P2 \$772 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$761 \$772 \$740 \$773 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$762 \$773 \$670 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$763 \$674 \$672 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$764 \$675 P3 \$775 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$765 \$775 \$741 \$776 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$766 \$776 \$691 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$767 \$695 \$693 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$768 GND \$874 \$859 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U AS=0.725P
+ AD=0.725P PS=5.58U PD=5.58U
M$769 \$860 \$859 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U AS=0.725P
+ AD=0.725P PS=5.58U PD=5.58U
M$770 GND \$872 up GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U AS=0.725P
+ AD=0.725P PS=5.58U PD=5.58U
M$771 \$874 \$872 GND GND sky130_fd_pr__nfet_01v8 L=0.2U W=2U AS=0.58P AD=0.29P
+ PS=4.58U PD=2.29U
M$772 GND \$875 \$874 GND sky130_fd_pr__nfet_01v8 L=0.2U W=2U AS=0.29P AD=0.58P
+ PS=2.29U PD=4.58U
M$773 dn \$875 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U AS=0.725P
+ AD=0.725P PS=5.58U PD=5.58U
M$774 GND \$862 \$861 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U AS=0.725P
+ AD=0.725P PS=5.58U PD=5.58U
M$775 \$862 \$874 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2.5U AS=0.725P
+ AD=0.725P PS=5.58U PD=5.58U
M$776 GND \$634 \$783 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$777 GND \$653 \$794 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$778 \$657 \$740 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$779 GND \$741 \$800 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$780 \$800 \$740 \$660 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$781 GND \$660 \$803 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$782 \$803 \$657 \$664 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$783 GND \$674 \$820 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$784 \$820 \$740 \$703 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$785 GND \$703 \$807 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$786 \$807 \$657 \$670 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$787 \$704 \$741 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$788 GND \$467 \$810 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$789 \$810 \$741 \$681 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$790 GND \$681 \$813 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$791 \$813 \$704 \$684 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$792 GND \$695 \$815 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$793 \$815 \$741 \$706 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$794 GND \$706 \$818 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$795 \$818 \$704 \$691 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$796 vctrl vn vctrl GND sky130_fd_pr__nfet_01v8_lvt L=8U W=17U AS=4.93P
+ AD=2.465P PS=34.58U PD=17.29U
M$797 vctrl vp vctrl GND sky130_fd_pr__nfet_01v8_lvt L=8U W=17U AS=2.465P
+ AD=4.93P PS=17.29U PD=34.58U
M$798 GND \$35 \$17 GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5U W=4.2U AS=1.218P
+ AD=1.218P PS=14.2U PD=14.2U
M$808 \$30 \$17 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=20U W=0.42U AS=0.1218P
+ AD=0.1218P PS=1.42U PD=1.42U
M$809 \$35 \$36 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5U W=1.68U AS=0.3654P
+ AD=0.3654P PS=4.26U PD=4.26U
M$810 GND \$36 \$36 GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5U W=1.68U AS=0.3654P
+ AD=0.3654P PS=4.26U PD=4.26U
Q$817 GND GND \$203 GND sky130_fd_pr__pnp_05v5_W0p68L0p68 AE=3.6992P PE=21.76U
+ AB=4.3681P PB=8.36U AC=4.3681P PC=8.36U NE=8
Q$818 GND GND \$24 GND sky130_fd_pr__pnp_05v5_W0p68L0p68 AE=0.4624P PE=2.72U
+ AB=4.3681P PB=8.36U AC=4.3681P PC=8.36U NE=1
R$826 VDD VDD VDD 17264.1509434 sky130_fd_pr__res_iso_pw L=30U W=5.3U
R$827 \$9 \$174 VDD 23018.8679245 sky130_fd_pr__res_iso_pw L=60U W=7.95U
R$828 \$52 \$121 VDD 11509.4339623 sky130_fd_pr__res_iso_pw L=30U W=7.95U
R$837 GND GND GND 1620.94607173 sky130_fd_pr__res_xhigh_po_1p41
+ L=7.07137723794U W=8.725U
R$844 GND \$24 GND 100482.269504 sky130_fd_pr__res_xhigh_po_1p41 L=70.84U
+ W=1.41U
R$846 \$29 \$203 GND 28709.2198582 sky130_fd_pr__res_xhigh_po_1p41 L=20.24U
+ W=1.41U
R$852 GND \$29 GND 100482.269504 sky130_fd_pr__res_xhigh_po_1p41 L=70.84U
+ W=1.41U
R$865 \$15 VOP GND 6468.08510638 sky130_fd_pr__res_xhigh_po_1p41 L=4.56U W=1.41U
R$872 vctrl VOP GND 90553.1914894 sky130_fd_pr__res_xhigh_po_1p41 L=63.84U
+ W=1.41U
C$874 \$15 GND 4.97289984e-10 sky130_fd_pr__model__cap_mim A=248644.992P
+ P=35680U
C$1066 GND VOP 2.5120144e-11 sky130_fd_pr__model__cap_mim A=12560.072P P=2004.8U
C$1076 vn vp 3.64e-13 sky130_fd_pr__model__cap_mim A=182P P=54U
C$1151 vctrl GND 1.74227e-12 sky130_fd_pr__model__cap_mim A=871.135P P=118.06U

.ENDS integer_pll
