** Test bench for BGR

.include ../spice_files/BGR_cir.ckt


.lib /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice ss
.temp -40.00
.options tnom=-40.00

VDD VDD GND 1.62
VTuner out GND 0.80


xvco out GND VDD BGR_Banba

**** begin user architecture code

.control
    set wr_singlescale
    set wr_vecnames
    set appendwrite

    op
    let Iref = i(VTuner)
    print Iref
    print all

   
    
.endc

.GLOBAL GND
.GLOBAL VDD
.end