** divider  cdl

.subckt DIVIDER VDD fout0 GND p2 p7 p1 p6 p5 p4 p3 p0 fin modo

*FIRST CELL
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_2
M_div_0 fout0 2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_1 fout0 1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_2 fout0 2 div_net1 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M_div_3 div_net1 1 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M_div_4 31 fout0 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_5 31 modi0 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_6 31 modi0 div_net2 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_7 div_net2 fout0 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M8 3 31 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M9 3 31 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M_div_10 finb fin vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_11 finb fin gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M_div_12 2 fin vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_13 2 p0 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_14 2 p0 div_net1_nand3 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_15 div_net1_nand3 fin div_net2_nand3 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_16 2 modo vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_17 div_net2_nand3 modo gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M_div_18 div_net1_ff1 fout0 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_19 div_net3_ff1 finb div_net1_ff1 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_20 div_net3_ff1 fin div_net2_ff1 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_21 div_net2_ff1 fout0 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_22 div_net4_ff1 div_net3_ff1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_23 1 fin div_net4_ff1 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_24 1 finb div_net5_ff1 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_25 div_net5_ff1 div_net3_ff1 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M_div_26 div_net1_ff2 3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_27 div_net3_ff2 finb div_net1_ff2 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_28 div_net3_ff2 fin div_net2_ff2 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_29 div_net2_ff2 3 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_30 div_net4_ff2 div_net3_ff2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_31 modo fin div_net4_ff2 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_32 modo finb div_net5_ff2 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_33 div_net5_ff2 div_net3_ff2 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1



*********************************///////////////SECOND CELL\\\\\\\\\\\\\*****************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_2
M_div_100 fout1 201 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_101 fout1 101 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_102 fout1 201 div_net1 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M_div_103 div_net1 101 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M_div_104 3101 fout1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_105 3101 modi1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_106 3101 modi1 div_net201 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_107 div_net201 fout1 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_108 301 3101 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_109 301 3101 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M_div_110 finb01 fout0 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_111 finb01 fout0 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M_div_112 201 fout0 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_113 201 p1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_114 201 p1 div_net1_nand301 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_115 div_net1_nand301 fout0 div_net2_nand301 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_116 291 modi0 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_117 div_net2_nand301 modi0 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M_div_118 div_net1_ff101 fout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_119 div_net3_ff101 finb01 div_net1_ff101 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_120 div_net3_ff101 fout0 div_net2_ff101 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_121 div_net2_ff101 fout1 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_122 div_net4_ff101 div_net3_ff101 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_123 101 fout0 div_net4_ff101 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_124 101 finb01 div_net5_ff101 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_125 div_net5_ff101 div_net3_ff101 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M_div_126 div_net1_ff201 301 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_127 div_net3_ff201 finb01 div_net1_ff201 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_128 div_net3_ff201 fout0 div_net2_ff201 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_129 div_net2_ff201 301 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_130 div_net4_ff201 div_net3_ff201 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_131 modi0 fout0 div_net4_ff201 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_132 modi0 finb01 div_net5_ff201 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_133 div_net5_ff201 div_net3_ff201 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1



*********************************///////////////THIRD CELL\\\\\\\\\\\\\*****************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_2
M_div_200 fout2 202 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_201 fout2 102 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_202 fout2 202 div_net1 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M_div_203 div_net1 102 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M_div_204 3102 fout2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_205 3102 modi2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_206 3102 modi2 div_net202 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_207 div_net202 fout2 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_208 302 3102 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_209 302 3102 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M_div_210 finb02 fout1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_211 finb02 fout1 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M_div_212 202 fout1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_213 202 p2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_214 202 p2 div_net1_nand302 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_215 div_net1_nand302 fout1 div_net2_nand302 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_216 291 modi1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_217 div_net2_nand302 modi1 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M_div_218 div_net1_ff102 fout2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_219 div_net3_ff102 finb02 div_net1_ff102 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_220 div_net3_ff102 fout1 div_net2_ff102 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_221 div_net2_ff102 fout2 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_222 div_net4_ff102 div_net3_ff102 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_223 102 fout1 div_net4_ff102 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_224 102 finb02 div_net5_ff102 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_225 div_net5_ff102 div_net3_ff102 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M_div_226 div_net1_ff202 302 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_227 div_net3_ff202 finb02 div_net1_ff202 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_228 div_net3_ff202 fout1 div_net2_ff202 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_229 div_net2_ff202 302 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_230 div_net4_ff202 div_net3_ff202 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_231 modi1 fout1 div_net4_ff202 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_232 modi1 finb02 div_net5_ff202 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_233 div_net5_ff202 div_net3_ff202 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1



*********************************///////////////FOURTH CELL\\\\\\\\\\\\\*****************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************


** NAND_2
M_div_300 fout3 203 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_301 fout3 103 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_302 fout3 203 div_net1 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M_div_303 div_net1 103 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M_div_304 3103 fout3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_305 3103 modi3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_306 3103 modi3 div_net203 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_307 div_net203 fout3 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_308 303 3103 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_309 303 3103 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M_div_310 finb03 fout2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_311 finb03 fout2 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M_div_312 203 fout2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_313 203 p3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_314 203 p3 div_net1_nand303 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_315 div_net1_nand303 fout2 div_net2_nand303 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_316 291 modi2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_317 div_net2_nand303 modi2 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M_div_318 div_net1_ff103 fout3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_319 div_net3_ff103 finb03 div_net1_ff103 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_320 div_net3_ff103 fout2 div_net2_ff103 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_321 div_net2_ff103 fout3 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_322 div_net4_ff103 div_net3_ff103 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_323 103 fout2 div_net4_ff103 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_324 103 finb03 div_net5_ff103 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_325 div_net5_ff103 div_net3_ff103 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M_div_326 div_net1_ff203 303 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_327 div_net3_ff203 finb03 div_net1_ff203 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_328 div_net3_ff203 fout2 div_net2_ff203 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_329 div_net2_ff203 303 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_330 div_net4_ff203 div_net3_ff203 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_331 modi2 fout2 div_net4_ff203 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_332 modi2 finb03 div_net5_ff203 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_333 div_net5_ff203 div_net3_ff203 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1


*********************************///////////////FIFTH CELL\\\\\\\\\\\\\*****************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_2
M_div_400 fout4 204 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_401 fout4 104 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_402 fout4 204 div_net1 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M_div_403 div_net1 104 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M_div_404 3104 fout4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_405 3104 modi4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_406 3104 modi4 div_net204 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_407 div_net204 fout4 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_408 304 3104 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_409 304 3104 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M_div_410 finb04 fout3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_411 finb04 fout3 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M_div_412 204 fout3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_413 204 p4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_414 204 p4 div_net1_nand304 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_415 div_net1_nand304 fout3 div_net2_nand304 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_416 291 modi3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_417 div_net2_nand304 modi3 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M_div_418 div_net1_ff104 fout4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_419 div_net3_ff104 finb04 div_net1_ff104 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_420 div_net3_ff104 fout3 div_net2_ff104 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_421 div_net2_ff104 fout4 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_422 div_net4_ff104 div_net3_ff104 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_423 104 fout3 div_net4_ff104 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_424 104 finb04 div_net5_ff104 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_425 div_net5_ff104 div_net3_ff104 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M_div_426 div_net1_ff204 304 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_427 div_net3_ff204 finb04 div_net1_ff204 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_428 div_net3_ff204 fout3 div_net2_ff204 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_429 div_net2_ff204 304 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_430 div_net4_ff204 div_net3_ff204 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_431 modi3 fout3 div_net4_ff204 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_432 modi3 finb04 div_net5_ff204 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_433 div_net5_ff204 div_net3_ff204 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*********************************///////////////SIXTHS CELL\\\\\\\\\\\\\*****************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_2
M_div_500 fout5 205 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_501 fout5 105 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_502 fout5 205 div_net1 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M_div_503 div_net1 105 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M_div_504 3105 fout5 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_505 3105 modi5 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_506 3105 modi5 div_net205 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_507 div_net205 fout5 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_508 305 3105 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_509 305 3105 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M_div_510 finb05 fout4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_511 finb05 fout4 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M_div_512 205 fout4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_513 205 p5 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_514 205 p5 div_net1_nand305 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_515 div_net1_nand305 fout4 div_net2_nand305 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_516 291 modi4 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_517 div_net2_nand305 modi4 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M_div_518 div_net1_ff105 fout5 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_519 div_net3_ff105 finb05 div_net1_ff105 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_520 div_net3_ff105 fout4 div_net2_ff105 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_521 div_net2_ff105 fout5 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_522 div_net4_ff105 div_net3_ff105 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_523 105 fout4 div_net4_ff105 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_524 105 finb05 div_net5_ff105 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_525 div_net5_ff105 div_net3_ff105 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M_div_526 div_net1_ff205 305 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_527 div_net3_ff205 finb05 div_net1_ff205 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_528 div_net3_ff205 fout4 div_net2_ff205 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_529 div_net2_ff205 305 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_530 div_net4_ff205 div_net3_ff205 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_531 modi4 fout4 div_net4_ff205 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_532 modi4 finb05 div_net5_ff205 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_533 div_net5_ff205 div_net3_ff205 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*********************************///////////////SEVENTH CELL\\\\\\\\\\\\\*****************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_2
M_div_600 fout6 206 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_601 fout6 106 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_602 fout6 206 div_net1 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M_div_603 div_net1 106 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M_div_604 3106 fout6 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_605 3106 modi6 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_606 3106 modi6 div_net206 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_607 div_net206 fout6 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_608 306 3106 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_609 306 3106 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M_div_610 finb06 fout5 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_611 finb06 fout5 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M_div_612 206 fout5 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_613 206 p6 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_614 206 p6 div_net1_nand306 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_615 div_net1_nand306 fout5 div_net2_nand306 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_616 291 modi5 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_617 div_net2_nand306 modi5 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M_div_618 div_net1_ff106 fout6 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_619 div_net3_ff106 finb06 div_net1_ff106 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_620 div_net3_ff106 fout5 div_net2_ff106 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_621 div_net2_ff106 fout6 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_622 div_net4_ff106 div_net3_ff106 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_623 106 fout5 div_net4_ff106 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_624 106 finb06 div_net5_ff106 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_625 div_net5_ff106 div_net3_ff106 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M_div_626 div_net1_ff206 306 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_627 div_net3_ff206 finb06 div_net1_ff206 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_628 div_net3_ff206 fout5 div_net2_ff206 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_629 div_net2_ff206 306 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_630 div_net4_ff206 div_net3_ff206 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_631 modi5 fout5 div_net4_ff206 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_632 modi5 finb06 div_net5_ff206 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_633 div_net5_ff206 div_net3_ff206 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1



*********************************///////////////EIGHTS CELL\\\\\\\\\\\\\*****************************************
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_2
M_div_700 fout 207 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_701 fout 107 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_702 fout 207 div_net1 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
M_div_703 div_net1 107 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** AND
M_div_704 3107 fout vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_705 3107 modi vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_706 3107 modi div_net207 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_707 div_net207 fout gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_708 307 3107 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_709 307 3107 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** INV
M_div_710 finb07 fout6 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_711 finb07 fout6 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** NAND_3
*M D G S B
M_div_712 207 fout6 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_713 207 p7 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1

M_div_714 207 p7 div_net1_nand307 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_715 div_net1_nand307 fout6 div_net2_nand307 gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

M_div_716 291 modi6 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_717 div_net2_nand307 modi6 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15U W=6U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 1 
M_div_718 div_net1_ff107 fout VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_719 div_net3_ff107 finb07 div_net1_ff107 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_720 div_net3_ff107 fout6 div_net2_ff107 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_721 div_net2_ff107 fout GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_722 div_net4_ff107 div_net3_ff107 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_723 107 fout6 div_net4_ff107 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_724 107 finb07 div_net5_ff107 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_725 div_net5_ff107 div_net3_ff107 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

*****************************************************************************************************************
*****************************************************************************************************************
*****************************************************************************************************************
** FF 2
M_div_726 div_net1_ff207 307 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_727 div_net3_ff207 finb07 div_net1_ff207 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_728 div_net3_ff207 fout6 div_net2_ff207 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_729 div_net2_ff207 307 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1

M_div_730 div_net4_ff207 div_net3_ff207 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_731 modi6 fout6 div_net4_ff207 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_div_732 modi6 finb07 div_net5_ff207 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1
M_div_733 div_net5_ff207 div_net3_ff207 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U nf=1 m=1


.ends