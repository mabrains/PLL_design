** sch_path: /home/ahmed/PLL_Internship/Ahmed Elshahat LC VCO/CMOS_LC_VCO/CMOS_VCO_tb1.sch
**.subckt CMOS_VCO_tb1

.param w1 = 10
.param w2 = 20
.param w3 = 40
.param w4 = 40
.param w5 = 40
.param w6 = 40
.param ISS = 4.5m
.param Rp = 400
.param Rs = 1.6
.param L = 1.6n


VDD VDD GND 1.8



XM1 net2 net2 GND GND sky130_fd_pr__nfet_01v8_lvt L=1 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=20

XM2 net1 net2 GND GND sky130_fd_pr__nfet_01v8_lvt L=1 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=20

XM3 vn vp net1 net1 sky130_fd_pr__nfet_01v8_lvt L=0.35 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1

XM4 vp vn net1 net1 sky130_fd_pr__nfet_01v8_lvt L=0.35 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1

XM5 vn vp VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=4

XM6 vp vn VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=4

I0 VDD net2 dc=ISS
L1 vn net3 1.6n m=1
R2 vp net3 1.6 m=1
R3 vp vn 400 m=1

XCF vp vn sky130_fd_pr__cap_mim_m3_1 W=10 L=2.3 MF=1 m=1
XC3 vn GND sky130_fd_pr__cap_mim_m3_1 W=1 L=1.95 MF=1 m=1
XC2 vp GND sky130_fd_pr__cap_mim_m3_1 W=1 L=1.95 MF=1 m=1
XC_load vp vn sky130_fd_pr__cap_mim_m3_1 W=30 L=38.6 MF=1 m=1



**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD



.tran 0.01ns 75ns
.save all
*.measure tran tperiod TRIG par('(v(vp)-v(vn))') VAL=0.5 RISE=6 TARG par('(v(vp)-v(vn))')
*+ VAL=0.5 RISE=7
*.measure tran ypp PP v(vp) from=30n to=50n

.control


op
save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[id]

let Id1 = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
let Id2 = @m.xm2.msky130_fd_pr__nfet_01v8_lvt[id]
let Id3 = @m.xm3.msky130_fd_pr__nfet_01v8_lvt[id]
let Id4 = @m.xm4.msky130_fd_pr__nfet_01v8_lvt[id]
let Id5 = @m.xm5.msky130_fd_pr__pfet_01v8_lvt[id]
let Id6 = @m.xm6.msky130_fd_pr__pfet_01v8_lvt[id]

let vgs1 = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vgs]
let vgs2 = @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vgs]
let vgs3 = @m.xm3.msky130_fd_pr__nfet_01v8_lvt[vgs]
let vgs4 = @m.xm4.msky130_fd_pr__nfet_01v8_lvt[vgs]
let vgs5 = @m.xm5.msky130_fd_pr__pfet_01v8_lvt[vgs]
let vgs6 = @m.xm6.msky130_fd_pr__pfet_01v8_lvt[vgs]

let vds1 = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vds]
let vds2 = @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vds]
let vds3 = @m.xm3.msky130_fd_pr__nfet_01v8_lvt[vds]
let vds4 = @m.xm4.msky130_fd_pr__nfet_01v8_lvt[vds]
let vds5 = @m.xm5.msky130_fd_pr__pfet_01v8_lvt[vds]
let vds6 = @m.xm6.msky130_fd_pr__pfet_01v8_lvt[vds]

let vth1 = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vth]
let vth2 = @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vth]
let vth3 = @m.xm3.msky130_fd_pr__nfet_01v8_lvt[vth]
let vth4 = @m.xm4.msky130_fd_pr__nfet_01v8_lvt[vth]
let vth5 = @m.xm5.msky130_fd_pr__pfet_01v8_lvt[vth]
let vth6 = @m.xm6.msky130_fd_pr__pfet_01v8_lvt[vth]

let gm1 = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm2 = @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm3 = @m.xm3.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm4 = @m.xm4.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm5 = @m.xm5.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm6 = @m.xm6.msky130_fd_pr__pfet_01v8_lvt[gm]

let gds1 = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gds]
let gds2 = @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gds]
let gds3 = @m.xm3.msky130_fd_pr__nfet_01v8_lvt[gds]
let gds4 = @m.xm4.msky130_fd_pr__nfet_01v8_lvt[gds]
let gds5 = @m.xm5.msky130_fd_pr__pfet_01v8_lvt[gds]
let gds6 = @m.xm6.msky130_fd_pr__pfet_01v8_lvt[gds]

let ro1 = 1/gds1
let ro2 = 1/gds2
let ro3 = 1/gds3
let ro4 = 1/gds4
let ro5 = 1/gds5
let ro6 = 1/gds6


let cgd3 = @m.xm3.msky130_fd_pr__nfet_01v8_lvt[cgd]
let cgd4 = @m.xm4.msky130_fd_pr__nfet_01v8_lvt[cgd] 
let cgd5 = @m.xm5.msky130_fd_pr__pfet_01v8_lvt[cgd] 
let cgd6 = @m.xm6.msky130_fd_pr__pfet_01v8_lvt[cgd] 

let cgs3 = @m.xm3.msky130_fd_pr__nfet_01v8_lvt[cgs]
let cgs4 = @m.xm4.msky130_fd_pr__nfet_01v8_lvt[cgs] 
let cgs5 = @m.xm5.msky130_fd_pr__pfet_01v8_lvt[cgs] 
let cgs6 = @m.xm6.msky130_fd_pr__pfet_01v8_lvt[cgs] 

let cgb3 = @m.xm3.msky130_fd_pr__nfet_01v8_lvt[cgb]
let cgb4 = @m.xm4.msky130_fd_pr__nfet_01v8_lvt[cgb] 
let cgb5 = @m.xm5.msky130_fd_pr__pfet_01v8_lvt[cgb] 
let cgb6 = @m.xm6.msky130_fd_pr__pfet_01v8_lvt[cgb] 

let cdb3 = @m.xm3.msky130_fd_pr__nfet_01v8_lvt[cdb]
let cdb4 = @m.xm4.msky130_fd_pr__nfet_01v8_lvt[cdb] 
let cdb5 = @m.xm5.msky130_fd_pr__pfet_01v8_lvt[cdb] 
let cdb6 = @m.xm6.msky130_fd_pr__pfet_01v8_lvt[cdb] 

let cds3 = @m.xm3.msky130_fd_pr__nfet_01v8_lvt[cds]
let cds4 = @m.xm4.msky130_fd_pr__nfet_01v8_lvt[cds] 
let cds5 = @m.xm5.msky130_fd_pr__pfet_01v8_lvt[cds] 
let cds6 = @m.xm6.msky130_fd_pr__pfet_01v8_lvt[cds] 

let CNMOS1 = 4*cgd3 + cgs3 + cgb3+ cdb3 + cds3
let CNMOS2 = 4*cgd4 + cgs4 + cgb4+ cdb4 + cds4

let CPMOS1 = 4*cgd5 + cgs5 + cgb5+ cdb5 + cds5
let CPMOS2 = 4*cgd6 + cgs6 + cgb6+ cdb6 + cds6

echo ===================Id==================
print Id1 Id2 Id3 Id4 Id5 Id6

echo ===================vds=================
print vds1 vds2 vds3 vds4 vds5 vds6

echo ===================vgs=================
print vgs1 vgs2 vgs3 vgs4 vgs5 vgs6

echo ===================on_check===========
print vgs1-vth1 vgs2-vth2 vgs3-vth3 vgs4-vth4 vgs5-vth5 vgs6-vth6

echo ===================sat_check===========
print vds1-vgs1+vth1 vds2-vgs2+vth2 vds3-vgs3+vth3 vds4-vgs4+vth4 vds5-vgs5+vth5 vds6-vgs6+vth6

echo ===================gm==================
print gm1 gm2 gm3 gm4 gm5 gm6

echo ===================gds=================
print gds1 gds2 gds3 gds4 gds5 gds6

echo ===================ro=================
print ro1 ro2 ro3 ro4 ro5 ro6

echo ===================vout================
print vp vn

echo ===================g_active/tank==================
let gactive = 0.25*(gm3+gm4+gm5+gm6)
let gtank = 0.25*(gds3+gds4+gds5+gds6) + 1/400 
print gactive gtank gactive/gtank 

echo ===================Capacitances==================
let cF = 50e-15
let C1 = 25e-15
let C_tank = -0.25*(CNMOS1+CNMOS2+CPMOS1+CPMOS2)+cF+0.5*c1
let c_load_255G = 1/(1.6e-9*(2*(22/7)*2.55e9)*(2*(22/7)*2.55e9)) - C_tank
let c_load_235G = 1/(1.6e-9*(2*(22/7)*2.35e9)*(2*(22/7)*2.35e9)) - C_tank
let delta_c = c_load_235G - c_load_255G
print CNMOS1 CNMOS2  CPMOS1 CPMOS2 cF c1 C_tank c_load_255G c_load_235G delta_c

echo ===================Transient================================================

*run
tran 0.01ns 250ns
*plot v(vn)  
*plot v(vp)  
*plot v(vp)-v(vn)
*let vp_max =  vecmax(vp)
*let vn_max =  vecmax(vn)
let vdiff_max =  vecmax(vp-vn)
print vdiff_max
*echo ===================swing===============
*print vp_max vn_max vdiff_max

*save @m.xm2.msky130_fd_pr__nfet_01v8_lvt[id]
*plot @m.xm2.msky130_fd_pr__nfet_01v8_lvt[id]




quit
.endc
.end



*=============================sweep ISS===================================
*compose  iss_vector   start=1m          stop=10m          step=0.1m
*let iss_counter = 0
*let swingvec = vector(length(iss_vector))
*let curr_value = iss_vector[0]
*set appendwrite


*while iss_counter < length(iss_vector)
 *   print curr_value
 *   alter I0  $&curr_value
 *   tran 0.01ns 75ns
 *   *plot vp-vn
 *   let max_swing = vecmax(vp-vn)
 *   
 *   setplot op1
 *   let swingvec[iss_counter] = tran.max_swing
 *   wrdata csv_files/swing_vs_ISS.csv swingvec[iss_counter]
 *   reset
 *   let iss_counter = iss_counter + 1
 *   let curr_value = iss_vector[iss_counter]
*end
*print swingvec


*=============================sweep RP===================================
*set appendwrite
*let vdiff_max =  vecmax(vp-vn)
*setplot const
*let swing_value = tran1.vdiff_max
*wrdata csv_files/swing_vs_L.csv swing_value