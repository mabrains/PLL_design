

*########################### 1/2 DIV behave ###############################
.subckt 1_2div VDD gnd MODOa MODIa FIn FOUT Pa

+ TR=1e-15 TF=1e-15

	* Analog to Digital nodes Models
	.model adc_buff adc_bridge(in_low = 0.9 in_high = 0.9)

	* Digital INPUT
	aref [FIn Pa MODIa] [FI P MODI] adc_buff

	*Define the and gate
	a_andGate [MODI FO] 2 and1
	.model and1 d_and(rise_delay = TR fall_delay = TF
	+ input_load = 0 )

	*Define the NAND 
	a_nandGate3 [FI P MODO] 1 nand1
	a_nandGate2 [3 1] FO nand1
	.model nand1 d_nand(rise_delay = TR fall_delay = TF
	+ input_load = 0 )


	* * Define the ff from lateches 2latches 
	XDFF_2latches1 FO FI 3 DFF_2latches
	XDFF_2latches2 2 FI MODO DFF_2latches


	* Digital to Analog nodes Models
	abridge-w1 [FO MODO] [FOUT MODOa] dac1 
	.model dac1 dac_bridge(out_low = 0 out_high = 1.8 out_undef = 0.9
	+ input_load = 0 t_rise = 1e-15
	+ t_fall = 1e-15)

.ends 1_2DIV

*########################### 1/2 DIV behave ###############################
.subckt DFF_2latches DATA_D CLK_D OUT


   ainv232 CLK_D CLK_D_bar invd1
   
   
   aL1 DATA_D CLK_D set reset OUT1 OUT1_bar latch1
   
   aL2 OUT1 CLK_D_bar set reset OUT OUT_bar latch1
   
   
   .model latch1 d_dlatch(data_delay = 1p enable_delay = 0
   + set_delay = 0
   + reset_delay = 0 ic = 0
   + rise_delay = 1p fall_delay = 1p)

.ends DFF_2latches
