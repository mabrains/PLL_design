* Circuit Model for DIVIDER

*########################### 1/2 DIV behave ###############################
.subckt 1_2div VDD gnd MODO MODI FIn FOUT P

+ TR=8.5e-12 TF=8.5e-12

	* Analog to Digital nodes Models
	.model adc_buff adc_bridge(in_low = 0.9 in_high = 0.9)

	* Digital INPUT
	aref [FIn] [FI] adc_buff

	*Define the and gate
	a_andGate [MODI FO] 2 and1

	.model and1 d_and(rise_delay = TR fall_delay = TF
	+ input_load = 0.5e-12 )

	*Define the NAND 
	a_nandGate3 [FI P MODO] 1 nand1
	a_nandGate2 [3 1] FO nand1

	.model nand1 d_nand(rise_delay = TR fall_delay = TF
	+ input_load = 0.5e-12)


	*Define FF D OUT CLK CLKb
	* XSS_FF1 OUT_AND MODO FI FIB SS_FF
	* XSS_FF2 FO OUTFF_IN_NAND FI FIB SS_FF

	*Define FF D CLK SET RESET out out-

	*Define the flip flops
	aF1 FO FI d_d0 d_d0 3 3_ flop1

	aF2 2 FI d_d0 d_d0 MODO MOD0_ flop1

	.model flop1 d_dff(clk_delay = 1e-15 set_delay = 1e-15
	+ reset_delay = 1e-15 ic = 0 rise_delay = TR
	+ fall_delay = TF )
	
	* Digital to Analog nodes Models
	abridge-w1 [FO] [FOUT] dac1 
	.model dac1 dac_bridge(out_low = 0 out_high = 1.8 out_undef = 0.9
	+ input_load = 1e-15 t_rise = 1e-15
	+ t_fall = 1e-15)

.ends 1_2DIV

*########################### 1/2 DIV behave ###############################

*########################### 1/2 DIV ideal ###############################
.param div=2

.subckt 1_2DIV_lib FIn FOUT

	* Analog to Digital nodes Models
	.model adc_buff adc_bridge(in_low = 0.9 in_high = 0.9)

	* Digital INPUT
	aref [FIn] [FI] adc_buff

	adivtest FI FO divider
	* .model divider d_fdiv(div_factor = 'divisor' high_cycles = 'divisor/2'
	* + i_count = 0 rise_delay = 1-e9
	* + fall_delay = 1e-9)
	.model divider d_fdiv(div_factor = 'div' high_cycles = 'div/2'
	+ i_count = 0 rise_delay = 8.5e-12
	+ fall_delay = 8.5e-12)


	* Digital to Analog nodes Models
	* Digital to Analog nodes Models
	abrigediev1 [FO] [FOUT] dac1 

	.model dac1 dac_bridge(out_low = 0 out_high = 1.8 out_undef = 0.9
	+ input_load = 1e-15 t_rise = 1e-15
	+ t_fall = 1e-15)

.ends  1_2div_lib
*########################### 1/2 DIV ideal ###############################

*########################### Static FF ###################################
* .subckt SFF D OUT CLK CLKb

* 	*LATCH
* 	* D CLK SET RESET OUT OUT_
* 	aTG1 D CLK d_d0 d_d0 1 1_ latch1
* 	aTG2 3 CLKb d_d0 d_d0 1 1_ latch1
* 	aTG3 2 CLKb d_d0 d_d0 4 4_ latch1
* 	aTG4 5 CLK d_d0 d_d0 4 4_ latch1

* 	.model latch1 d_dlatch(data_delay = 1e-15 enable_delay = 1e-15
* 	+ set_delay = 1e-15
* 	+ reset_delay = 1e-15 ic = 0
* 	+ rise_delay = 1e-15 fall_delay = 1e-15

* 	*
* 	*Define Inverter

* 	.model invd1 d_inverter(rise_delay = 1e-10 fall_delay = 1e-10)
* 	a_a1 1 2 invd1
* 	a_a2 2 3 invd1
* 	a_a3 4 OUT invd1
* 	a_a4 OUT 5 invd1

* .ends SFF

*########################### Static FF ###################################

*########################### 8 (2to1) DIVIDER ###################################

.subckt divider VDD gnd modo modi Fin Fout P0 P1 P2 P3 P4 P5 P6 P7

	X1_2div1 VDD gnd modo m1 Fin F1 P0 1_2div
	X1_2div2 VDD gnd m1 m2 F1 F2 P1 1_2div
	X1_2div3 VDD gnd m2 m3 F2 F3 P2 1_2div
	X1_2div4 VDD gnd m3 m4 F3 F4 P3 1_2div
	X1_2div5 VDD gnd m4 m5 F4 F5 P4 1_2div
	X1_2div6 VDD gnd m5 m6 F5 F6 P5 1_2div
	X1_2div7 VDD gnd m6 m7 F6 F7 P6 1_2div
	X1_2div8 VDD gnd m7 modid F7 Fout P7 1_2div

.ends divider

*########################### 8 (2to1) DIVIDER ###################################
