** sch_path: /home/tarek/Mabrains/Inv/Crystal.sch
**.subckt Crystal
.include ../xschem/ring_cir.ckt
V1 VDD GND PWL(0 0 1u 1.8 1m 1.8)
xring Vin out VDD GND ring
**** begin user architecture code

** opencircuitdesign pdks install
.lib /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt



.control
tran 5n 1m
plot out
meas tran tperiod TRIG out VAL=0.9 RISE=750 TARG out VAL=0.9 RISE=751
let freq = 1/(tperiod*1000000)
print freq
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
