** sch_path: /home/ahmed/Mabrains_internship/VCO_Try3/VCO_Full_Phase_Noise.sch
**.subckt VCO_Full_Phase_Noise
VDD VDD GND 1.8
XM8 net3 net22 GND GND sky130_fd_pr__nfet_01v8 L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
XM9 net1 net23 GND GND sky130_fd_pr__nfet_01v8 L=1 W=25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
XM11 vp net24 net4 net4 sky130_fd_pr__pfet_01v8 L=0.15 W=50 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
XM1 vn net19 net4 net4 sky130_fd_pr__pfet_01v8 L=0.15 W=50 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
XM2 vp net20 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
L1 vp net37 4n m=1
R1 net35 vn 1182 m=1
R2 net36 vn 3 m=1
XM7 vn net21 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
C1 vp vn 5f m=10
C3 vp GND 5f m=5
C2 vn GND 5f m=5
VTuner net6 GND 0.2
C13 vp vn 10f m=34
XM6 net6 vn net6 GND sky130_fd_pr__nfet_01v8_lvt L=1.8 W=12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
XM3 net6 vp net6 GND sky130_fd_pr__nfet_01v8_lvt L=1.8 W=12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
XM4 net4 net5 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=50 m=50
XM5 net1 net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
XM13 net8 net25 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM14 VBE net26 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XQ10 GND GND VBE sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ2 GND GND net7 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ3 GND GND net7 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ4 GND GND net7 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ5 GND GND net7 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ6 GND GND net7 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ7 GND GND net7 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ8 GND GND net7 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ9 GND GND net7 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XR4 net38 net8 GND sky130_fd_pr__res_xhigh_po_1p41 L=20 mult=1 m=1
XM15 net10 net27 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM16 net11 net28 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=44 m=44
XM17 net12 net29 net10 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6
XM18 net9 net30 net10 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6
XM19 net11 net31 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
XM20 net12 net32 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM21 net9 net33 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM22 net13 net14 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM23 net13 net15 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=20 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM24 VBE net34 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XR3 net16 net8 net16 sky130_fd_pr__res_xhigh_po_1p41 L=70 mult=1 m=1
XR5 net17 VBE net17 sky130_fd_pr__res_xhigh_po_1p41 L=70 mult=1 m=1
XM10 net3 net18 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=40 m=40


V1 net19 vp DC 0 trnoise (0 0 0 0)
V2 net20 vn DC 0 trnoise (0 0 0 0)
V4 net5 net1 DC 0 trnoise (0 0 0 0)
V5 net2 net1 DC 0 trnoise (0 0 0 0)
V7 net21 vp DC 0 trnoise (0 0 0 0)
V8 net22 net3 DC 0 trnoise (0 0 0 0)
V9 net23 net3 DC 0 trnoise (0 0 0 0)
V10 net18 net11 DC 0 trnoise (0 0 0 0)
V11 net24 vn DC 0 trnoise (0 0 0 0)
V13 net25 net11 DC 0 trnoise (0 0 0 0)
V14 net26 net11 DC 0 trnoise (0 0 0 0)
V15 net27 net11 DC 0 trnoise (0 0 0 0)
V16 net28 net11 DC 0 trnoise (0 0 0 0)
V17 net29 net8 DC 0 trnoise (0 0 0 0)
V18 net30 VBE DC 0 trnoise (0 0 0 0)
V19 net31 net12 DC 0 trnoise (0 0 0 0)
V20 net32 net9 DC 0 trnoise (0 0 0 0)
V21 net33 net9 DC 0 trnoise (0 0 0 0)
V22 net14 net11 DC 0 trnoise (0 0 0 0)
V23 net15 net11 DC 0 trnoise (0 0 0 0)
V24 net34 net13 DC 0 trnoise (0 0 0 0)
VR1 net35 vp DC 0 trnoise (0 0 0 0)
VR2 net36 net37 DC 0 trnoise (0 0 0 0)
VR3 net16 GND DC 0 trnoise (0 0 0 0)
VR4 net38 net7 DC 0 trnoise (0 0 0 0)
VR5 net17 GND DC 0 trnoise (0 0 0 0)


**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


.tran 0.01n 0.03u
.save all
.control
op
  save @m.xm1.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm11.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm2.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm4.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm5.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm7.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm8.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm9.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm10.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm13.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm14.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm15.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm16.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm17.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm18.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm19.msky130_fd_pr__nfet_g5v0d10v5[gm]
  save @m.xm20.msky130_fd_pr__nfet_g5v0d10v5[gm]
  save @m.xm21.msky130_fd_pr__nfet_g5v0d10v5[gm]
  save @m.xm23.msky130_fd_pr__nfet_g5v0d10v5[gm]
  save @m.xm22.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm24.msky130_fd_pr__pfet_g5v0d10v5[gm]
  
run
  save @m.xm1.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm11.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm2.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm4.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm5.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm7.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm8.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm9.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm10.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm13.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm14.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm15.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm16.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm17.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm18.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm19.msky130_fd_pr__nfet_g5v0d10v5[gm]
  save @m.xm20.msky130_fd_pr__nfet_g5v0d10v5[gm]
  save @m.xm21.msky130_fd_pr__nfet_g5v0d10v5[gm]
  save @m.xm23.msky130_fd_pr__nfet_g5v0d10v5[gm]
  save @m.xm22.msky130_fd_pr__pfet_g5v0d10v5[gm]
  save @m.xm24.msky130_fd_pr__pfet_g5v0d10v5[gm]
  
  
  let vdiff = v(vp)-v(vn)
  save vdiff
  *plot vdiff
  linearize vdiff
  *save vdiff
  *fft (v(vp)-v(vn))
  fft vdiff
  
  wrdata gm1_no_noise.csv tran1.@m.xm1.msky130_fd_pr__pfet_01v8[gm]
  wrdata gm11_no_noise.csv tran1.@m.xm11.msky130_fd_pr__pfet_01v8[gm]
  wrdata gm2_no_noise.csv tran1.@m.xm2.msky130_fd_pr__nfet_01v8[gm]
  wrdata gm4_no_noise.csv tran1.@m.xm4.msky130_fd_pr__pfet_01v8[gm]
  wrdata gm5_no_noise.csv tran1.@m.xm5.msky130_fd_pr__pfet_01v8[gm]
  wrdata gm7_no_noise.csv tran1.@m.xm7.msky130_fd_pr__nfet_01v8[gm]
  wrdata gm8_no_noise.csv tran1.@m.xm8.msky130_fd_pr__nfet_01v8[gm]
  wrdata gm9_no_noise.csv tran1.@m.xm9.msky130_fd_pr__nfet_01v8[gm]
  wrdata gm10_no_noise.csv tran1.@m.xm10.msky130_fd_pr__pfet_g5v0d10v5[gm]
  wrdata gm13_no_noise.csv tran1.@m.xm13.msky130_fd_pr__pfet_g5v0d10v5[gm]
  wrdata gm14_no_noise.csv tran1.@m.xm14.msky130_fd_pr__pfet_g5v0d10v5[gm]
  wrdata gm15_no_noise.csv tran1.@m.xm15.msky130_fd_pr__pfet_g5v0d10v5[gm]
  wrdata gm16_no_noise.csv tran1.@m.xm16.msky130_fd_pr__pfet_g5v0d10v5[gm]
  wrdata gm17_no_noise.csv tran1.@m.xm17.msky130_fd_pr__pfet_g5v0d10v5[gm]
  wrdata gm18_no_noise.csv tran1.@m.xm18.msky130_fd_pr__pfet_g5v0d10v5[gm]
  wrdata gm19_no_noise.csv tran1.@m.xm19.msky130_fd_pr__nfet_g5v0d10v5[gm]
  wrdata gm20_no_noise.csv tran1.@m.xm20.msky130_fd_pr__nfet_g5v0d10v5[gm]
  wrdata gm21_no_noise.csv tran1.@m.xm21.msky130_fd_pr__nfet_g5v0d10v5[gm]
  wrdata gm23_no_noise.csv tran1.@m.xm23.msky130_fd_pr__nfet_g5v0d10v5[gm]
  wrdata gm22_no_noise.csv tran1.@m.xm22.msky130_fd_pr__pfet_g5v0d10v5[gm]
  wrdata gm24_no_noise.csv tran1.@m.xm24.msky130_fd_pr__pfet_g5v0d10v5[gm]
  
  plot mag(sp2.vdiff)
  
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
