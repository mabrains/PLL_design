* Extracted by KLayout with SKY130 LVS runset on : 20/10/2022 14:31

.SUBCKT CP
X$1 \$429 \$731 via_new$1
X$2 \$429 \$731 via_new
M$1 \$55 \$72 \$56 \$50 sky130_fd_pr__pfet_01v8 L=0.15 W=2 AS=0.58 AD=0.58
+ PS=4.58 PD=4.58
M$2 \$31 \$75 \$91 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314 AD=1.9314
+ PS=13.9 PD=13.9
M$3 \$33 \$75 \$93 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314 AD=1.9314
+ PS=13.9 PD=13.9
M$4 \$34 \$75 \$97 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314 AD=1.9314
+ PS=13.9 PD=13.9
M$5 \$14 \$75 \$102 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$6 \$37 \$75 \$107 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$7 \$38 \$75 \$142 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$8 \$112 \$75 \$115 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$9 \$40 \$75 \$119 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$10 \$43 \$75 \$121 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$11 \$125 \$75 \$126 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$12 \$44 \$75 \$131 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$13 \$46 \$75 \$135 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$14 \$48 \$75 \$143 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$15 \$9 \$313 \$286 \$8 sky130_fd_pr__pfet_01v8 L=0.6 W=4 AS=1.16 AD=1.16
+ PS=8.58 PD=8.58
M$16 \$335 \$365 VON \$8 sky130_fd_pr__pfet_01v8 L=0.15 W=1 AS=0.29 AD=0.29
+ PS=2.58 PD=2.58
M$17 \$9 \$313 \$287 \$8 sky130_fd_pr__pfet_01v8 L=0.6 W=4 AS=1.16 AD=1.16
+ PS=8.58 PD=8.58
M$18 \$326 \$365 VON \$8 sky130_fd_pr__pfet_01v8 L=0.15 W=1 AS=0.29 AD=0.29
+ PS=2.58 PD=2.58
M$19 \$398 \$451 \$430 \$10 sky130_fd_pr__pfet_01v8 L=0.15 W=4 AS=1.16 AD=1.16
+ PS=8.58 PD=8.58
M$20 \$398 \$452 \$431 \$10 sky130_fd_pr__pfet_01v8 L=0.15 W=4 AS=1.16 AD=1.16
+ PS=8.58 PD=8.58
M$21 \$453 \$514 \$592 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$22 \$455 \$514 \$596 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$23 \$458 \$514 \$598 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$24 \$432 \$514 \$602 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$25 \$459 \$514 \$628 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$26 \$461 \$514 \$608 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$27 \$196 \$192 \$199 \$1 sky130_fd_pr__pfet_01v8 L=0.15 W=10 AS=2.9 AD=2.9
+ PS=20.58 PD=20.58
M$28 \$196 \$193 \$203 \$1 sky130_fd_pr__pfet_01v8 L=0.15 W=10 AS=2.9 AD=2.9
+ PS=20.58 PD=20.58
M$29 \$463 \$514 \$611 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$30 \$465 \$514 \$614 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$31 \$434 \$514 \$617 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$32 \$468 \$514 \$621 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$33 \$470 \$514 \$623 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$34 \$471 \$514 \$627 \$1 sky130_fd_pr__pfet_01v8 L=0.6 W=6.66 AS=1.9314
+ AD=1.9314 PS=13.9 PD=13.9
M$35 \$699 \$708 \$695 \$693 sky130_fd_pr__pfet_01v8 L=0.15 W=2 AS=0.58 AD=0.58
+ PS=4.58 PD=4.58
M$36 \$80 \$72 \$82 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 AS=0.29
+ AD=0.29 PS=2.58 PD=2.58
M$37 \$179 \$252 \$211 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$38 \$179 \$252 \$214 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$39 \$179 \$252 \$217 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$40 \$178 \$252 \$220 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$41 \$179 \$252 \$248 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$42 \$179 \$252 \$249 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$43 \$149 \$252 \$228 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$44 \$179 \$252 \$231 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$45 \$179 \$252 \$250 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$46 \$178 \$252 \$237 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$47 \$179 \$252 \$241 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$48 \$179 \$252 \$244 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$49 \$179 \$252 \$247 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$50 \$491 \$449 \$440 sky130_gnd sky130_fd_pr__nfet_01v8 L=1 W=1.3 AS=0.377
+ AD=0.377 PS=3.18 PD=3.18
M$51 \$402 \$391 VON sky130_gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 AS=0.29
+ AD=0.29 PS=2.58 PD=2.58
M$52 \$404 \$391 VON sky130_gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 AS=0.29
+ AD=0.29 PS=2.58 PD=2.58
M$53 \$491 \$449 \$442 sky130_gnd sky130_fd_pr__nfet_01v8 L=1 W=1.3 AS=0.377
+ AD=0.377 PS=3.18 PD=3.18
M$54 \$342 \$290 \$341 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 AS=0.29
+ AD=0.29 PS=2.58 PD=2.58
M$55 \$342 \$316 \$344 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 AS=0.29
+ AD=0.29 PS=2.58 PD=2.58
M$56 \$501 \$568 \$559 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$57 \$501 \$568 \$523 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$58 \$500 \$568 \$526 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$59 \$501 \$568 \$529 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$60 \$488 \$568 \$532 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$61 \$501 \$568 \$535 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$62 \$501 \$568 \$538 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$63 \$436 \$568 \$560 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$64 \$501 \$568 \$543 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$65 \$501 \$568 \$561 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$66 \$488 \$568 \$562 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$67 \$501 \$568 \$563 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$68 \$500 \$568 \$552 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$69 \$501 \$568 \$555 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$70 \$501 \$568 \$558 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.6 W=2 AS=0.58
+ AD=0.58 PS=4.58 PD=4.58
M$71 VON \$665 \$629 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.15 W=4 AS=1.16
+ AD=1.16 PS=8.58 PD=8.58
M$72 \$292 \$669 \$629 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.15 W=4 AS=1.16
+ AD=1.16 PS=8.58 PD=8.58
M$73 \$715 \$708 \$717 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 AS=0.29
+ AD=0.29 PS=2.58 PD=2.58
R$74 \$294 \$294 \$294 sky130_fd_pr__res_iso_pw R=41208.8888889 L=30.4 W=2.25
+ A=79.5 P=65.3
R$75 \$447 \$448 \$294 sky130_fd_pr__res_iso_pw R=41208.8888889 L=30.4 W=2.25
+ A=79.5 P=65.3
R$76 \$447 \$448 \$294 sky130_fd_pr__res_iso_pw R=41208.8888889 L=30.4 W=2.25
+ A=79.5 P=65.3
R$77 \$379 \$157 \$294 sky130_fd_pr__res_iso_pw R=41208.8888889 L=30.4 W=2.25
+ A=79.5 P=65.3
R$78 \$379 \$157 \$294 sky130_fd_pr__res_iso_pw R=41208.8888889 L=30.4 W=2.25
+ A=79.5 P=65.3
R$79 \$21 \$321 \$294 sky130_fd_pr__res_iso_pw R=41208.8888889 L=30.4 W=2.25
+ A=79.5 P=65.3
R$80 \$379 \$157 \$294 sky130_fd_pr__res_iso_pw R=41208.8888889 L=30.4 W=2.25
+ A=79.5 P=65.3
R$81 \$21 \$321 \$294 sky130_fd_pr__res_iso_pw R=41208.8888889 L=30.4 W=2.25
+ A=79.5 P=65.3
R$82 \$447 \$448 \$294 sky130_fd_pr__res_iso_pw R=41208.8888889 L=30.4 W=2.25
+ A=79.5 P=65.3
R$83 \$21 \$321 \$294 sky130_fd_pr__res_iso_pw R=41208.8888889 L=30.4 W=2.25
+ A=79.5 P=65.3
R$84 \$294 \$294 \$294 sky130_fd_pr__res_iso_pw R=41208.8888889 L=30.4 W=2.25
+ A=79.5 P=65.3
.ENDS CP

.SUBCKT via_new$1 \$1 \$2
.ENDS via_new$1

.SUBCKT via_new \$1 \$2
.ENDS via_new
