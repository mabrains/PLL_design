* NGSPICE file created from DIV_CELL.ext - technology: sky130A

.subckt DIV_CELL net1_ff2 fin P modo net1 net1_nand3 net2 net2_nand3 net1_ff1 net2_ff1
+ net4_ff1 net5_ff1 net4_ff2 net2_ff2 net5_ff2 2 1 3 modi fout 31 finb net3_ff1 net3_ff2
+ VDD GND
X0 VDD.t14 2.t4 fout.t1 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1 net1_ff1.t0 fout.t3 VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2 GND.t7 modo.t2 net2_nand3.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X3 net2.t1 modi.t0 31.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X4 net4_ff1.t1 net3_ff1.t2 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X5 net1_nand3.t0 P.t0 2.t2 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X6 net5_ff2.t0 net3_ff2.t2 GND.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X7 GND.t11 31.t3 3.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 net3_ff1.t1 finb.t2 net1_ff1.t1 VDD.t23 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9 VDD.t8 modi.t1 31.t2 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X10 net1.t1 2.t5 fout.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X11 GND.t10 fin.t0 finb.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 VDD.t22 1.t2 fout.t2 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13 net3_ff1.t0 fin.t1 net2_ff1.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 modo.t1 finb.t3 net5_ff2.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X15 VDD.t10 fin.t2 2.t1 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X16 GND.t1 1.t3 net1.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X17 modo.t0 fin.t3 net4_ff2.t1 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X18 net3_ff2.t0 fin.t4 net2_ff2.t1 GND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 1.t0 fin.t5 net4_ff1.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X20 net2_ff1.t1 fout.t4 GND.t9 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X21 GND.t8 fout.t5 net2.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X22 1.t1 finb.t4 net5_ff1.t0 GND.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 net2_nand3.t0 fin.t6 net1_nand3.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X24 net5_ff1.t1 net3_ff1.t3 GND.t4 GND.t3 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X25 net3_ff2.t1 finb.t5 net4_ff2 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.716e+07u w=4e+06u l=150000u
X26 finb.t1 fin.t7 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X27 net4_ff2.t3 net3_ff2.t3 VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X28 VDD.t4 modo.t3 2.t0 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X29 net4_ff2 3.t2 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X30 net2_ff2.t0 3.t3 GND.t6 GND.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X31 VDD.t25 P.t1 2.t3 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X32 VDD.t16 fout.t6 31.t0 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X33 3.t0 31.t4 VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
R0 2.n0 2.t5 1040.28
R1 2.n0 2.t4 794.529
R2 2.n188 2.n187 13.176
R3 2.n336 2.t0 11.614
R4 2.n336 2.t1 11.298
R5 2.n337 2.t3 10.376
R6 2.n8 2.n6 9.3
R7 2.n310 2.n309 9.3
R8 2.n56 2.n55 9.3
R9 2.n58 2.n57 9.3
R10 2.n115 2.n114 9.3
R11 2.n112 2.n111 9.3
R12 2.n70 2.n69 9.3
R13 2.n68 2.n67 9.3
R14 2.n194 2.n193 9.3
R15 2.n93 2.n92 9.3
R16 2.n101 2.n100 9.3
R17 2.n104 2.n103 9.3
R18 2.n224 2.n223 9.3
R19 2.n221 2.n220 9.3
R20 2.n305 2.n304 9.3
R21 2.n303 2.n302 9.3
R22 2.n296 2.n295 8.097
R23 2.n103 2.n102 5.457
R24 2.n223 2.n222 5.08
R25 2.n294 2.n293 4.65
R26 2.n233 2.n232 4.65
R27 2.n315 2.n308 4.5
R28 2.n289 2.n288 4.5
R29 2.n282 2.n281 4.5
R30 2.n213 2.n212 4.5
R31 2.n203 2.n202 4.5
R32 2.n190 2.n189 4.5
R33 2.n166 2.n165 4.5
R34 2.n98 2.n90 4.5
R35 2.n121 2.n120 4.5
R36 2.n66 2.n65 4.5
R37 2.n78 2.n77 4.5
R38 2.n85 2.n84 4.5
R39 2.n129 2.n128 4.5
R40 2.n109 2.n108 4.5
R41 2.n275 2.n274 4.5
R42 2.n54 2.n53 4.5
R43 2.n324 2.n321 4.5
R44 2.n11 2.n10 4.5
R45 2.n77 2.n75 4.314
R46 2.n128 2.n125 3.944
R47 2.n288 2.n287 3.937
R48 2.n274 2.n273 3.567
R49 2.n234 2.n227 3.033
R50 2.n298 2.n297 3.033
R51 2.n295 2.t2 2.9
R52 2.n127 2.n126 2.258
R53 2.n272 2.n271 2.258
R54 2.n83 2.n82 1.882
R55 2.n84 2.n83 1.882
R56 2.n280 2.n279 1.882
R57 2 2.n338 1.829
R58 2 2.n0 1.566
R59 2.n274 2.n272 1.505
R60 2.n281 2.n280 1.505
R61 2.n316 2.n315 1.5
R62 2.n167 2.n166 1.5
R63 2.n204 2.n203 1.5
R64 2.n235 2.n234 1.5
R65 2.n214 2.n213 1.5
R66 2.n325 2.n324 1.5
R67 2.n12 2.n11 1.5
R68 2.n338 2.n335 1.477
R69 2.n53 2.n52 1.129
R70 2.n128 2.n127 1.129
R71 2.n120 2.n119 1.129
R72 2.n130 2.n129 1.042
R73 2.n338 2.n337 1.022
R74 2.n147 2.n146 0.853
R75 2.n237 2.n236 0.853
R76 2.n331 2.n330 0.853
R77 2.n24 2.n23 0.853
R78 2.n10 2.n9 0.752
R79 2.n202 2.n201 0.752
R80 2.n212 2.n211 0.752
R81 2.n288 2.n286 0.752
R82 2.n308 2.n307 0.752
R83 2.n321 2.n320 0.752
R84 2.n14 2.n13 0.717
R85 2.n193 2.n192 0.536
R86 2.n92 2.n91 0.536
R87 2.n114 2.n113 0.475
R88 2.n232 2.n231 0.475
R89 2.n297 2.n296 0.382
R90 2.n64 2.n63 0.382
R91 2.n65 2.n64 0.376
R92 2.n77 2.n76 0.376
R93 2.n108 2.n107 0.376
R94 2.n90 2.n89 0.376
R95 2.n165 2.n164 0.376
R96 2.n189 2.n188 0.376
R97 2.n52 2.n51 0.349
R98 2.n307 2.n306 0.349
R99 2.n337 2.n336 0.316
R100 2.n105 2.n104 0.047
R101 2.n95 2.n94 0.047
R102 2.n184 2.n183 0.047
R103 2.n197 2.n196 0.047
R104 2.n225 2.n224 0.047
R105 2.n312 2.n311 0.047
R106 2.n291 2.n290 0.043
R107 2.n260 2.n259 0.043
R108 2.n74 2.n73 0.041
R109 2.n41 2.n40 0.041
R110 2.n300 2.n299 0.035
R111 2.n168 2.n167 0.035
R112 2.n173 2.n172 0.035
R113 2.n266 2.n265 0.035
R114 2.n61 2.n60 0.034
R115 2.n182 2.n181 0.034
R116 2.n186 2.n185 0.034
R117 2.n303 2.n301 0.034
R118 2.n21 2.n20 0.034
R119 2.n19 2.n18 0.034
R120 2.n137 2.n136 0.034
R121 2.n144 2.n143 0.034
R122 2.n204 2.n180 0.034
R123 2.n206 2.n205 0.034
R124 2.n219 2.n218 0.034
R125 2.n268 2.n267 0.034
R126 2.n59 2.n58 0.032
R127 2.n234 2.n233 0.032
R128 2.n298 2.n294 0.032
R129 2.n142 2.n141 0.032
R130 2.n316 2.n268 0.032
R131 2.n26 2.n25 0.031
R132 2.n37 2.n36 0.031
R133 2.n149 2.n148 0.031
R134 2.n160 2.n159 0.031
R135 2.n239 2.n238 0.031
R136 2.n250 2.n249 0.031
R137 2.n333 2.n332 0.031
R138 2.n68 2.n66 0.03
R139 2.n112 2.n110 0.03
R140 2.n97 2.n96 0.03
R141 2.n199 2.n198 0.03
R142 2.n313 2.n312 0.03
R143 2.n22 2.n21 0.03
R144 2.n16 2.n15 0.03
R145 2.n140 2.n139 0.03
R146 2.n178 2.n177 0.03
R147 2.n207 2.n206 0.03
R148 2.n263 2.n262 0.03
R149 2.n330 2.n329 0.03
R150 2.n11 2.n8 0.028
R151 2.n49 2.n48 0.028
R152 2.n72 2.n71 0.028
R153 2.n87 2.n86 0.028
R154 2.n129 2.n88 0.028
R155 2.n118 2.n117 0.028
R156 2.n234 2.n226 0.028
R157 2.n278 2.n277 0.028
R158 2.n292 2.n291 0.028
R159 2.n315 2.n305 0.028
R160 2.n12 2.n4 0.028
R161 2.n39 2.n38 0.028
R162 2.n46 2.n45 0.028
R163 2.n130 2.n47 0.028
R164 2.n135 2.n134 0.028
R165 2.n145 2.n144 0.028
R166 2.n162 2.n161 0.028
R167 2.n175 2.n174 0.028
R168 2.n236 2.n235 0.028
R169 2.n255 2.n254 0.028
R170 2.n261 2.n260 0.028
R171 2.n326 2.n325 0.028
R172 2.n30 2.n29 0.027
R173 2.n33 2.n32 0.027
R174 2.n153 2.n152 0.027
R175 2.n156 2.n155 0.027
R176 2.n243 2.n242 0.027
R177 2.n246 2.n245 0.027
R178 2.n56 2.n54 0.026
R179 2.n109 2.n106 0.026
R180 2.n229 2.n228 0.026
R181 2.n276 2.n275 0.026
R182 2.n132 2.n131 0.026
R183 2.n146 2.n138 0.026
R184 2.n217 2.n216 0.026
R185 2.n253 2.n252 0.026
R186 2.n258 2.n257 0.026
R187 2.n328 2.n327 0.026
R188 2.n13 2.n12 0.024
R189 2.n116 2.n115 0.024
R190 2.n233 2.n230 0.024
R191 2.n3 2.n2 0.024
R192 2.n43 2.n42 0.024
R193 2.n138 2.n137 0.024
R194 2.n171 2.n170 0.024
R195 2.n214 2.n208 0.024
R196 2.n80 2.n79 0.022
R197 2.n106 2.n105 0.022
R198 2.n194 2.n191 0.022
R199 2.n230 2.n229 0.022
R200 2.n285 2.n284 0.022
R201 2.n2 2.n1 0.022
R202 2.n146 2.n145 0.022
R203 2.n170 2.n169 0.022
R204 2.n235 2.n219 0.022
R205 2.n218 2.n217 0.022
R206 2.n123 2.n122 0.02
R207 2.n121 2.n118 0.02
R208 2.n117 2.n116 0.02
R209 2.n226 2.n225 0.02
R210 2.n210 2.n209 0.02
R211 2.n23 2.n22 0.02
R212 2.n136 2.n135 0.02
R213 2.n236 2.n207 0.02
R214 2.n329 2.n328 0.02
R215 2.n325 2.n319 0.02
R216 2.n24 2.n14 0.019
R217 2.n25 2.n24 0.019
R218 2.n147 2.n37 0.019
R219 2.n148 2.n147 0.019
R220 2.n237 2.n160 0.019
R221 2.n238 2.n237 0.019
R222 2.n331 2.n250 0.019
R223 2.n332 2.n331 0.019
R224 2.n294 2.n292 0.018
R225 2.n44 2.n43 0.018
R226 2.n330 2.n316 0.018
R227 2.n71 2.n70 0.017
R228 2.n99 2.n98 0.017
R229 2.n96 2.n95 0.017
R230 2.n323 2.n322 0.017
R231 2.n131 2.n130 0.017
R232 2.n134 2.n133 0.017
R233 2.n143 2.n142 0.017
R234 2.n141 2.n140 0.017
R235 2.n216 2.n215 0.017
R236 2.n257 2.n256 0.017
R237 2.n262 2.n261 0.017
R238 2.n319 2.n318 0.017
R239 2.n50 2.n49 0.015
R240 2.n60 2.n59 0.015
R241 2.n88 2.n87 0.015
R242 2.n198 2.n197 0.015
R243 2.n203 2.n200 0.015
R244 2.n277 2.n276 0.015
R245 2.n282 2.n278 0.015
R246 2.n314 2.n313 0.015
R247 2.n20 2.n19 0.015
R248 2.n18 2.n17 0.015
R249 2.n47 2.n46 0.015
R250 2.n177 2.n176 0.015
R251 2.n180 2.n179 0.015
R252 2.n205 2.n204 0.015
R253 2.n254 2.n253 0.015
R254 2.n256 2.n255 0.015
R255 2.n62 2.n61 0.013
R256 2.n86 2.n85 0.013
R257 2.n101 2.n99 0.013
R258 2.n299 2.n298 0.013
R259 2.n301 2.n300 0.013
R260 2.n45 2.n44 0.013
R261 2.n265 2.n264 0.013
R262 2.n267 2.n266 0.013
R263 2.n335 2.n334 0.013
R264 2.n31 2.n30 0.012
R265 2.n32 2.n31 0.012
R266 2.n154 2.n153 0.012
R267 2.n155 2.n154 0.012
R268 2.n244 2.n243 0.012
R269 2.n245 2.n244 0.012
R270 2.n124 2.n123 0.011
R271 2.n28 2.n27 0.011
R272 2.n35 2.n34 0.011
R273 2.n151 2.n150 0.011
R274 2.n158 2.n157 0.011
R275 2.n241 2.n240 0.011
R276 2.n248 2.n247 0.011
R277 2.n8 2.n7 0.009
R278 2.n81 2.n80 0.009
R279 2.n85 2.n81 0.009
R280 2.n183 2.n182 0.009
R281 2.n284 2.n283 0.009
R282 2.n4 2.n3 0.009
R283 2.n169 2.n168 0.009
R284 2.n78 2.n74 0.007
R285 2.n166 2.n163 0.007
R286 2.n185 2.n184 0.007
R287 2.n191 2.n190 0.007
R288 2.n283 2.n282 0.007
R289 2.n311 2.n310 0.007
R290 2.n42 2.n41 0.007
R291 2.n167 2.n162 0.007
R292 2.n172 2.n171 0.007
R293 2.n174 2.n173 0.007
R294 2.n327 2.n326 0.007
R295 2.n318 2.n317 0.007
R296 2.n27 2.n26 0.006
R297 2.n29 2.n28 0.006
R298 2.n34 2.n33 0.006
R299 2.n36 2.n35 0.006
R300 2.n150 2.n149 0.006
R301 2.n152 2.n151 0.006
R302 2.n157 2.n156 0.006
R303 2.n159 2.n158 0.006
R304 2.n240 2.n239 0.006
R305 2.n242 2.n241 0.006
R306 2.n247 2.n246 0.006
R307 2.n249 2.n248 0.006
R308 2.n334 2.n333 0.006
R309 2.n54 2.n50 0.005
R310 2.n58 2.n56 0.005
R311 2.n129 2.n124 0.005
R312 2.n122 2.n121 0.005
R313 2.n94 2.n93 0.005
R314 2.n195 2.n194 0.005
R315 2.n270 2.n269 0.005
R316 2.n290 2.n289 0.005
R317 2.n215 2.n214 0.005
R318 2.n259 2.n258 0.005
R319 2.n11 2.n5 0.003
R320 2.n203 2.n199 0.003
R321 2.n224 2.n221 0.003
R322 2.n213 2.n210 0.003
R323 2.n289 2.n285 0.003
R324 2.n305 2.n303 0.003
R325 2.n315 2.n314 0.003
R326 2.n324 2.n323 0.003
R327 2.n133 2.n132 0.003
R328 2.n264 2.n263 0.003
R329 2.n66 2.n62 0.001
R330 2.n70 2.n68 0.001
R331 2.n73 2.n72 0.001
R332 2.n79 2.n78 0.001
R333 2.n115 2.n112 0.001
R334 2.n110 2.n109 0.001
R335 2.n104 2.n101 0.001
R336 2.n98 2.n97 0.001
R337 2.n190 2.n186 0.001
R338 2.n196 2.n195 0.001
R339 2.n275 2.n270 0.001
R340 2.n17 2.n16 0.001
R341 2.n40 2.n39 0.001
R342 2.n176 2.n175 0.001
R343 2.n179 2.n178 0.001
R344 2.n252 2.n251 0.001
R345 fout.n8 fout.t5 1037.29
R346 fout.n9 fout.t6 797.225
R347 fout.n378 fout.t3 732.331
R348 fout.n393 fout.t4 397.315
R349 fout.n218 fout.n217 13.176
R350 fout.n30 fout.t2 11.72
R351 fout.n30 fout.t1 10.993
R352 fout.n38 fout.n36 9.3
R353 fout.n340 fout.n339 9.3
R354 fout.n86 fout.n85 9.3
R355 fout.n88 fout.n87 9.3
R356 fout.n145 fout.n144 9.3
R357 fout.n142 fout.n141 9.3
R358 fout.n100 fout.n99 9.3
R359 fout.n98 fout.n97 9.3
R360 fout.n224 fout.n223 9.3
R361 fout.n123 fout.n122 9.3
R362 fout.n131 fout.n130 9.3
R363 fout.n134 fout.n133 9.3
R364 fout.n249 fout.n248 9.3
R365 fout.n246 fout.n245 9.3
R366 fout.n335 fout.n334 9.3
R367 fout.n333 fout.n332 9.3
R368 fout.n326 fout.n325 8.097
R369 fout.n133 fout.n132 5.457
R370 fout.n248 fout.n247 5.08
R371 fout.n324 fout.n323 4.65
R372 fout.n263 fout.n262 4.65
R373 fout.n345 fout.n338 4.5
R374 fout.n319 fout.n318 4.5
R375 fout.n312 fout.n311 4.5
R376 fout.n257 fout.n256 4.5
R377 fout.n233 fout.n232 4.5
R378 fout.n220 fout.n219 4.5
R379 fout.n196 fout.n195 4.5
R380 fout.n128 fout.n120 4.5
R381 fout.n151 fout.n150 4.5
R382 fout.n96 fout.n95 4.5
R383 fout.n108 fout.n107 4.5
R384 fout.n115 fout.n114 4.5
R385 fout.n159 fout.n158 4.5
R386 fout.n139 fout.n138 4.5
R387 fout.n305 fout.n304 4.5
R388 fout.n84 fout.n83 4.5
R389 fout.n354 fout.n351 4.5
R390 fout.n41 fout.n40 4.5
R391 fout.n107 fout.n105 4.314
R392 fout.n158 fout.n155 3.944
R393 fout.n318 fout.n317 3.937
R394 fout.n304 fout.n303 3.567
R395 fout.n264 fout.n252 3.033
R396 fout.n328 fout.n327 3.033
R397 fout.n325 fout.t0 2.9
R398 fout.n157 fout.n156 2.258
R399 fout.n302 fout.n301 2.258
R400 fout.n113 fout.n112 1.882
R401 fout.n114 fout.n113 1.882
R402 fout.n310 fout.n309 1.882
R403 fout.n366 fout.n30 1.516
R404 fout.n304 fout.n302 1.505
R405 fout.n311 fout.n310 1.505
R406 fout.n346 fout.n345 1.5
R407 fout.n197 fout.n196 1.5
R408 fout.n234 fout.n233 1.5
R409 fout.n265 fout.n264 1.5
R410 fout.n355 fout.n354 1.5
R411 fout.n42 fout.n41 1.5
R412 fout.n22 fout.n8 1.388
R413 fout.n10 fout.n9 1.354
R414 fout.n395 fout.n393 1.354
R415 fout.n379 fout.n378 1.354
R416 fout.n396 fout.n395 1.142
R417 fout.n397 fout.n396 1.138
R418 fout.n380 fout.n379 1.137
R419 fout.n406 fout.n405 1.137
R420 fout.n371 fout.n370 1.137
R421 fout.n402 fout.n401 1.137
R422 fout.n386 fout.n385 1.137
R423 fout.n408 fout.n407 1.136
R424 fout.n382 fout.n381 1.136
R425 fout.n83 fout.n82 1.129
R426 fout.n158 fout.n157 1.129
R427 fout.n150 fout.n149 1.129
R428 fout.n160 fout.n159 1.042
R429 fout.n177 fout.n176 0.853
R430 fout.n267 fout.n266 0.853
R431 fout.n361 fout.n360 0.853
R432 fout.n54 fout.n53 0.853
R433 fout.n410 fout.n29 0.827
R434 fout.n40 fout.n39 0.752
R435 fout.n232 fout.n231 0.752
R436 fout.n256 fout.n255 0.752
R437 fout.n318 fout.n316 0.752
R438 fout.n338 fout.n337 0.752
R439 fout.n351 fout.n350 0.752
R440 fout.n44 fout.n43 0.717
R441 fout.n366 fout.n365 0.69
R442 fout.n367 fout.n366 0.68
R443 fout.n223 fout.n222 0.536
R444 fout.n122 fout.n121 0.536
R445 fout.n144 fout.n143 0.475
R446 fout.n262 fout.n261 0.475
R447 fout.n410 fout.n409 0.471
R448 fout.n23 fout.n22 0.44
R449 fout.n327 fout.n326 0.382
R450 fout.n94 fout.n93 0.382
R451 fout.n95 fout.n94 0.376
R452 fout.n107 fout.n106 0.376
R453 fout.n138 fout.n137 0.376
R454 fout.n120 fout.n119 0.376
R455 fout.n195 fout.n194 0.376
R456 fout.n219 fout.n218 0.376
R457 fout.n82 fout.n81 0.349
R458 fout.n337 fout.n336 0.349
R459 fout fout.n410 0.124
R460 fout.n393 fout.n392 0.083
R461 fout.n378 fout.n377 0.083
R462 fout.n8 fout.n7 0.076
R463 fout.n4 fout.n3 0.059
R464 fout.n135 fout.n134 0.047
R465 fout.n125 fout.n124 0.047
R466 fout.n214 fout.n213 0.047
R467 fout.n227 fout.n226 0.047
R468 fout.n250 fout.n249 0.047
R469 fout.n342 fout.n341 0.047
R470 fout.n321 fout.n320 0.043
R471 fout.n290 fout.n289 0.043
R472 fout.n104 fout.n103 0.041
R473 fout.n71 fout.n70 0.041
R474 fout.n330 fout.n329 0.035
R475 fout.n198 fout.n197 0.035
R476 fout.n203 fout.n202 0.035
R477 fout.n296 fout.n295 0.035
R478 fout.n91 fout.n90 0.034
R479 fout.n212 fout.n211 0.034
R480 fout.n216 fout.n215 0.034
R481 fout.n333 fout.n331 0.034
R482 fout.n51 fout.n50 0.034
R483 fout.n49 fout.n48 0.034
R484 fout.n167 fout.n166 0.034
R485 fout.n174 fout.n173 0.034
R486 fout.n234 fout.n210 0.034
R487 fout.n236 fout.n235 0.034
R488 fout.n244 fout.n243 0.034
R489 fout.n298 fout.n297 0.034
R490 fout.n401 fout.n400 0.032
R491 fout.n18 fout.n17 0.032
R492 fout.n17 fout.n16 0.032
R493 fout.n89 fout.n88 0.032
R494 fout.n264 fout.n263 0.032
R495 fout.n328 fout.n324 0.032
R496 fout.n172 fout.n171 0.032
R497 fout.n346 fout.n298 0.032
R498 fout.n22 fout.n21 0.032
R499 fout.n56 fout.n55 0.031
R500 fout.n67 fout.n66 0.031
R501 fout.n179 fout.n178 0.031
R502 fout.n190 fout.n189 0.031
R503 fout.n269 fout.n268 0.031
R504 fout.n280 fout.n279 0.031
R505 fout.n363 fout.n362 0.031
R506 fout.n12 fout.n11 0.03
R507 fout.n98 fout.n96 0.03
R508 fout.n142 fout.n140 0.03
R509 fout.n127 fout.n126 0.03
R510 fout.n229 fout.n228 0.03
R511 fout.n343 fout.n342 0.03
R512 fout.n52 fout.n51 0.03
R513 fout.n46 fout.n45 0.03
R514 fout.n170 fout.n169 0.03
R515 fout.n208 fout.n207 0.03
R516 fout.n237 fout.n236 0.03
R517 fout.n293 fout.n292 0.03
R518 fout.n360 fout.n359 0.03
R519 fout.n392 fout.n391 0.028
R520 fout.n390 fout.n389 0.028
R521 fout.n375 fout.n374 0.028
R522 fout.n377 fout.n376 0.028
R523 fout.n385 fout.n384 0.028
R524 fout.n401 fout.n399 0.028
R525 fout.n405 fout.n404 0.028
R526 fout.n370 fout.n368 0.028
R527 fout.n21 fout.n20 0.028
R528 fout.n19 fout.n18 0.028
R529 fout.n16 fout.n15 0.028
R530 fout.n14 fout.n13 0.028
R531 fout.n41 fout.n38 0.028
R532 fout.n79 fout.n78 0.028
R533 fout.n102 fout.n101 0.028
R534 fout.n117 fout.n116 0.028
R535 fout.n159 fout.n118 0.028
R536 fout.n148 fout.n147 0.028
R537 fout.n264 fout.n251 0.028
R538 fout.n308 fout.n307 0.028
R539 fout.n322 fout.n321 0.028
R540 fout.n345 fout.n335 0.028
R541 fout.n42 fout.n34 0.028
R542 fout.n69 fout.n68 0.028
R543 fout.n76 fout.n75 0.028
R544 fout.n160 fout.n77 0.028
R545 fout.n165 fout.n164 0.028
R546 fout.n175 fout.n174 0.028
R547 fout.n192 fout.n191 0.028
R548 fout.n205 fout.n204 0.028
R549 fout.n266 fout.n265 0.028
R550 fout.n285 fout.n284 0.028
R551 fout.n291 fout.n290 0.028
R552 fout.n356 fout.n355 0.028
R553 fout.n60 fout.n59 0.027
R554 fout.n63 fout.n62 0.027
R555 fout.n183 fout.n182 0.027
R556 fout.n186 fout.n185 0.027
R557 fout.n273 fout.n272 0.027
R558 fout.n276 fout.n275 0.027
R559 fout.n7 fout.n6 0.026
R560 fout.n5 fout.n4 0.026
R561 fout.n3 fout.n2 0.026
R562 fout.n1 fout.n0 0.026
R563 fout.n86 fout.n84 0.026
R564 fout.n139 fout.n136 0.026
R565 fout.n259 fout.n258 0.026
R566 fout.n306 fout.n305 0.026
R567 fout.n162 fout.n161 0.026
R568 fout.n176 fout.n168 0.026
R569 fout.n242 fout.n241 0.026
R570 fout.n283 fout.n282 0.026
R571 fout.n288 fout.n287 0.026
R572 fout.n358 fout.n357 0.026
R573 fout.n43 fout.n42 0.024
R574 fout.n146 fout.n145 0.024
R575 fout.n263 fout.n260 0.024
R576 fout.n33 fout.n32 0.024
R577 fout.n73 fout.n72 0.024
R578 fout.n168 fout.n167 0.024
R579 fout.n201 fout.n200 0.024
R580 fout.n239 fout.n238 0.024
R581 fout.n26 fout.n25 0.023
R582 fout.n110 fout.n109 0.022
R583 fout.n136 fout.n135 0.022
R584 fout.n224 fout.n221 0.022
R585 fout.n260 fout.n259 0.022
R586 fout.n258 fout.n257 0.022
R587 fout.n315 fout.n314 0.022
R588 fout.n32 fout.n31 0.022
R589 fout.n176 fout.n175 0.022
R590 fout.n200 fout.n199 0.022
R591 fout.n265 fout.n244 0.022
R592 fout.n243 fout.n242 0.022
R593 fout.n153 fout.n152 0.02
R594 fout.n151 fout.n148 0.02
R595 fout.n147 fout.n146 0.02
R596 fout.n251 fout.n250 0.02
R597 fout.n254 fout.n253 0.02
R598 fout.n53 fout.n52 0.02
R599 fout.n166 fout.n165 0.02
R600 fout.n266 fout.n237 0.02
R601 fout.n359 fout.n358 0.02
R602 fout.n355 fout.n349 0.02
R603 fout.n54 fout.n44 0.019
R604 fout.n55 fout.n54 0.019
R605 fout.n177 fout.n67 0.019
R606 fout.n178 fout.n177 0.019
R607 fout.n267 fout.n190 0.019
R608 fout.n268 fout.n267 0.019
R609 fout.n361 fout.n280 0.019
R610 fout.n362 fout.n361 0.019
R611 fout.n324 fout.n322 0.018
R612 fout.n74 fout.n73 0.018
R613 fout.n360 fout.n346 0.018
R614 fout.n395 fout.n394 0.017
R615 fout.n385 fout.n383 0.017
R616 fout.n370 fout.n369 0.017
R617 fout.n379 fout.n373 0.017
R618 fout.n13 fout.n12 0.017
R619 fout.n11 fout.n10 0.017
R620 fout.n101 fout.n100 0.017
R621 fout.n129 fout.n128 0.017
R622 fout.n126 fout.n125 0.017
R623 fout.n353 fout.n352 0.017
R624 fout.n161 fout.n160 0.017
R625 fout.n164 fout.n163 0.017
R626 fout.n173 fout.n172 0.017
R627 fout.n171 fout.n170 0.017
R628 fout.n241 fout.n240 0.017
R629 fout.n287 fout.n286 0.017
R630 fout.n292 fout.n291 0.017
R631 fout.n349 fout.n348 0.017
R632 fout.n402 fout.n398 0.016
R633 fout.n406 fout.n403 0.016
R634 fout.n391 fout.n390 0.015
R635 fout.n376 fout.n375 0.015
R636 fout.n20 fout.n19 0.015
R637 fout.n15 fout.n14 0.015
R638 fout.n80 fout.n79 0.015
R639 fout.n90 fout.n89 0.015
R640 fout.n118 fout.n117 0.015
R641 fout.n228 fout.n227 0.015
R642 fout.n233 fout.n230 0.015
R643 fout.n307 fout.n306 0.015
R644 fout.n312 fout.n308 0.015
R645 fout.n344 fout.n343 0.015
R646 fout.n50 fout.n49 0.015
R647 fout.n48 fout.n47 0.015
R648 fout.n77 fout.n76 0.015
R649 fout.n207 fout.n206 0.015
R650 fout.n210 fout.n209 0.015
R651 fout.n235 fout.n234 0.015
R652 fout.n284 fout.n283 0.015
R653 fout.n286 fout.n285 0.015
R654 fout.n6 fout.n5 0.013
R655 fout.n2 fout.n1 0.013
R656 fout.n92 fout.n91 0.013
R657 fout.n116 fout.n115 0.013
R658 fout.n131 fout.n129 0.013
R659 fout.n329 fout.n328 0.013
R660 fout.n331 fout.n330 0.013
R661 fout.n75 fout.n74 0.013
R662 fout.n295 fout.n294 0.013
R663 fout.n297 fout.n296 0.013
R664 fout.n365 fout.n364 0.013
R665 fout.n407 fout.n402 0.012
R666 fout.n407 fout.n406 0.012
R667 fout.n61 fout.n60 0.012
R668 fout.n62 fout.n61 0.012
R669 fout.n184 fout.n183 0.012
R670 fout.n185 fout.n184 0.012
R671 fout.n274 fout.n273 0.012
R672 fout.n275 fout.n274 0.012
R673 fout.n388 fout.n387 0.011
R674 fout.n381 fout.n372 0.011
R675 fout.n154 fout.n153 0.011
R676 fout.n58 fout.n57 0.011
R677 fout.n65 fout.n64 0.011
R678 fout.n181 fout.n180 0.011
R679 fout.n188 fout.n187 0.011
R680 fout.n271 fout.n270 0.011
R681 fout.n278 fout.n277 0.011
R682 fout.n24 fout.n23 0.01
R683 fout.n25 fout.n24 0.01
R684 fout.n28 fout.n27 0.009
R685 fout.n38 fout.n37 0.009
R686 fout.n111 fout.n110 0.009
R687 fout.n115 fout.n111 0.009
R688 fout.n213 fout.n212 0.009
R689 fout.n314 fout.n313 0.009
R690 fout.n34 fout.n33 0.009
R691 fout.n199 fout.n198 0.009
R692 fout.n108 fout.n104 0.007
R693 fout.n196 fout.n193 0.007
R694 fout.n215 fout.n214 0.007
R695 fout.n221 fout.n220 0.007
R696 fout.n313 fout.n312 0.007
R697 fout.n341 fout.n340 0.007
R698 fout.n72 fout.n71 0.007
R699 fout.n197 fout.n192 0.007
R700 fout.n202 fout.n201 0.007
R701 fout.n204 fout.n203 0.007
R702 fout.n357 fout.n356 0.007
R703 fout.n348 fout.n347 0.007
R704 fout.n387 fout.n386 0.006
R705 fout.n372 fout.n371 0.006
R706 fout.n381 fout.n380 0.006
R707 fout.n57 fout.n56 0.006
R708 fout.n59 fout.n58 0.006
R709 fout.n64 fout.n63 0.006
R710 fout.n66 fout.n65 0.006
R711 fout.n180 fout.n179 0.006
R712 fout.n182 fout.n181 0.006
R713 fout.n187 fout.n186 0.006
R714 fout.n189 fout.n188 0.006
R715 fout.n270 fout.n269 0.006
R716 fout.n272 fout.n271 0.006
R717 fout.n277 fout.n276 0.006
R718 fout.n279 fout.n278 0.006
R719 fout.n364 fout.n363 0.006
R720 fout.n27 fout.n26 0.005
R721 fout.n29 fout.n28 0.005
R722 fout.n84 fout.n80 0.005
R723 fout.n88 fout.n86 0.005
R724 fout.n159 fout.n154 0.005
R725 fout.n152 fout.n151 0.005
R726 fout.n124 fout.n123 0.005
R727 fout.n225 fout.n224 0.005
R728 fout.n300 fout.n299 0.005
R729 fout.n320 fout.n319 0.005
R730 fout.n240 fout.n239 0.005
R731 fout.n289 fout.n288 0.005
R732 fout.n409 fout.n408 0.004
R733 fout.n382 fout.n367 0.003
R734 fout.n41 fout.n35 0.003
R735 fout.n233 fout.n229 0.003
R736 fout.n249 fout.n246 0.003
R737 fout.n257 fout.n254 0.003
R738 fout.n319 fout.n315 0.003
R739 fout.n335 fout.n333 0.003
R740 fout.n345 fout.n344 0.003
R741 fout.n354 fout.n353 0.003
R742 fout.n163 fout.n162 0.003
R743 fout.n294 fout.n293 0.003
R744 fout.n396 fout.n388 0.003
R745 fout.n408 fout.n397 0.002
R746 fout.n397 fout.n382 0.002
R747 fout.n96 fout.n92 0.001
R748 fout.n100 fout.n98 0.001
R749 fout.n103 fout.n102 0.001
R750 fout.n109 fout.n108 0.001
R751 fout.n145 fout.n142 0.001
R752 fout.n140 fout.n139 0.001
R753 fout.n134 fout.n131 0.001
R754 fout.n128 fout.n127 0.001
R755 fout.n220 fout.n216 0.001
R756 fout.n226 fout.n225 0.001
R757 fout.n305 fout.n300 0.001
R758 fout.n47 fout.n46 0.001
R759 fout.n70 fout.n69 0.001
R760 fout.n206 fout.n205 0.001
R761 fout.n209 fout.n208 0.001
R762 fout.n282 fout.n281 0.001
R763 VDD.t5 VDD.t7 282.282
R764 VDD.t11 VDD.t23 244.603
R765 VDD.t6 VDD.t1 243.985
R766 VDD.t21 VDD.t26 192.1
R767 VDD.n13 VDD.t0 180.981
R768 VDD.t1 VDD.t5 176.657
R769 VDD.t28 VDD.t6 176.657
R770 VDD.t0 VDD.t11 176.04
R771 VDD.t23 VDD.t17 176.04
R772 VDD.t15 VDD.t19 174.187
R773 VDD.t7 VDD.t15 160.598
R774 VDD.t13 VDD.t21 160.598
R775 VDD.n180 VDD.t24 158.127
R776 VDD.t3 VDD.t13 150.097
R777 VDD.t9 VDD.t3 123.537
R778 VDD.t24 VDD.t9 123.537
R779 VDD.n13 VDD.t28 109.947
R780 VDD.n101 VDD.n100 56.47
R781 VDD.n85 VDD.n84 56.47
R782 VDD.n252 VDD.n251 56.47
R783 VDD.n268 VDD.n267 56.47
R784 VDD.n112 VDD.n111 49.411
R785 VDD.n74 VDD.n73 49.411
R786 VDD.n241 VDD.n240 49.411
R787 VDD.n279 VDD.n278 49.411
R788 VDD.n18 VDD.n17 45.882
R789 VDD.n123 VDD.n122 42.352
R790 VDD.n63 VDD.n62 42.352
R791 VDD.n230 VDD.n229 42.352
R792 VDD.n290 VDD.n289 42.352
R793 VDD.n134 VDD.n133 35.294
R794 VDD.n52 VDD.n51 35.294
R795 VDD.n219 VDD.n218 35.294
R796 VDD.n301 VDD.n300 35.294
R797 VDD.n145 VDD.n144 28.235
R798 VDD.n41 VDD.n40 28.235
R799 VDD.n208 VDD.n207 28.235
R800 VDD.n312 VDD.n311 28.235
R801 VDD.n156 VDD.n155 21.176
R802 VDD.n30 VDD.n29 21.176
R803 VDD.n197 VDD.n196 21.176
R804 VDD.n323 VDD.n322 21.176
R805 VDD.n185 VDD.n184 20.411
R806 VDD.n333 VDD.n332 20.411
R807 VDD.n166 VDD.n165 20.411
R808 VDD.n182 VDD.n180 17.939
R809 VDD.n15 VDD.n13 17.939
R810 VDD.n196 VDD.n195 17.569
R811 VDD.n322 VDD.n321 17.569
R812 VDD.n29 VDD.n28 17.569
R813 VDD.n155 VDD.n154 17.569
R814 VDD.n207 VDD.n206 14.627
R815 VDD.n311 VDD.n310 14.627
R816 VDD.n40 VDD.n39 14.627
R817 VDD.n144 VDD.n143 14.627
R818 VDD.n167 VDD.n166 14.117
R819 VDD.n186 VDD.n185 14.117
R820 VDD.n334 VDD.n333 14.117
R821 VDD.n19 VDD.n18 12.531
R822 VDD.n218 VDD.n217 11.58
R823 VDD.n300 VDD.n299 11.58
R824 VDD.n51 VDD.n50 11.58
R825 VDD.n133 VDD.n132 11.58
R826 VDD.n20 VDD.n19 9.93
R827 VDD.n354 VDD.t12 9.536
R828 VDD.n0 VDD.t2 9.53
R829 VDD.n5 VDD.t8 9.51
R830 VDD.n176 VDD.t29 9.407
R831 VDD.n348 VDD.t27 9.393
R832 VDD.n347 VDD.t18 9.38
R833 VDD.n2 VDD.t20 9.363
R834 VDD.n2 VDD.t16 9.358
R835 VDD.n349 VDD.t22 9.358
R836 VDD.n350 VDD.t14 9.358
R837 VDD.n346 VDD.t4 9.358
R838 VDD.n345 VDD.t10 9.358
R839 VDD.n344 VDD.t25 9.358
R840 VDD.n190 VDD.n189 9.3
R841 VDD.n201 VDD.n200 9.3
R842 VDD.n212 VDD.n211 9.3
R843 VDD.n223 VDD.n222 9.3
R844 VDD.n234 VDD.n233 9.3
R845 VDD.n245 VDD.n244 9.3
R846 VDD.n256 VDD.n255 9.3
R847 VDD.n263 VDD.n262 9.3
R848 VDD.n274 VDD.n273 9.3
R849 VDD.n285 VDD.n284 9.3
R850 VDD.n296 VDD.n295 9.3
R851 VDD.n307 VDD.n306 9.3
R852 VDD.n318 VDD.n317 9.3
R853 VDD.n329 VDD.n328 9.3
R854 VDD.n338 VDD.n337 9.3
R855 VDD.n258 VDD.n257 9.3
R856 VDD.n247 VDD.n246 9.3
R857 VDD.n236 VDD.n235 9.3
R858 VDD.n225 VDD.n224 9.3
R859 VDD.n214 VDD.n213 9.3
R860 VDD.n203 VDD.n202 9.3
R861 VDD.n192 VDD.n191 9.3
R862 VDD.n261 VDD.n260 9.3
R863 VDD.n272 VDD.n271 9.3
R864 VDD.n283 VDD.n282 9.3
R865 VDD.n294 VDD.n293 9.3
R866 VDD.n305 VDD.n304 9.3
R867 VDD.n316 VDD.n315 9.3
R868 VDD.n327 VDD.n326 9.3
R869 VDD.n340 VDD.n339 9.3
R870 VDD.n188 VDD.n187 9.3
R871 VDD.n187 VDD.n186 9.3
R872 VDD.n199 VDD.n198 9.3
R873 VDD.n198 VDD.n197 9.3
R874 VDD.n210 VDD.n209 9.3
R875 VDD.n209 VDD.n208 9.3
R876 VDD.n221 VDD.n220 9.3
R877 VDD.n220 VDD.n219 9.3
R878 VDD.n232 VDD.n231 9.3
R879 VDD.n231 VDD.n230 9.3
R880 VDD.n243 VDD.n242 9.3
R881 VDD.n242 VDD.n241 9.3
R882 VDD.n254 VDD.n253 9.3
R883 VDD.n253 VDD.n252 9.3
R884 VDD.n270 VDD.n269 9.3
R885 VDD.n269 VDD.n268 9.3
R886 VDD.n281 VDD.n280 9.3
R887 VDD.n280 VDD.n279 9.3
R888 VDD.n292 VDD.n291 9.3
R889 VDD.n291 VDD.n290 9.3
R890 VDD.n303 VDD.n302 9.3
R891 VDD.n302 VDD.n301 9.3
R892 VDD.n314 VDD.n313 9.3
R893 VDD.n313 VDD.n312 9.3
R894 VDD.n325 VDD.n324 9.3
R895 VDD.n324 VDD.n323 9.3
R896 VDD.n336 VDD.n335 9.3
R897 VDD.n335 VDD.n334 9.3
R898 VDD.n342 VDD.n341 9.3
R899 VDD.n173 VDD.n172 9.3
R900 VDD.n162 VDD.n161 9.3
R901 VDD.n151 VDD.n150 9.3
R902 VDD.n140 VDD.n139 9.3
R903 VDD.n129 VDD.n128 9.3
R904 VDD.n118 VDD.n117 9.3
R905 VDD.n107 VDD.n106 9.3
R906 VDD.n96 VDD.n95 9.3
R907 VDD.n89 VDD.n88 9.3
R908 VDD.n78 VDD.n77 9.3
R909 VDD.n67 VDD.n66 9.3
R910 VDD.n56 VDD.n55 9.3
R911 VDD.n45 VDD.n44 9.3
R912 VDD.n34 VDD.n33 9.3
R913 VDD.n23 VDD.n22 9.3
R914 VDD.n25 VDD.n24 9.3
R915 VDD.n21 VDD.n20 9.3
R916 VDD.n36 VDD.n35 9.3
R917 VDD.n32 VDD.n31 9.3
R918 VDD.n31 VDD.n30 9.3
R919 VDD.n47 VDD.n46 9.3
R920 VDD.n43 VDD.n42 9.3
R921 VDD.n42 VDD.n41 9.3
R922 VDD.n58 VDD.n57 9.3
R923 VDD.n54 VDD.n53 9.3
R924 VDD.n53 VDD.n52 9.3
R925 VDD.n69 VDD.n68 9.3
R926 VDD.n65 VDD.n64 9.3
R927 VDD.n64 VDD.n63 9.3
R928 VDD.n80 VDD.n79 9.3
R929 VDD.n76 VDD.n75 9.3
R930 VDD.n75 VDD.n74 9.3
R931 VDD.n91 VDD.n90 9.3
R932 VDD.n87 VDD.n86 9.3
R933 VDD.n86 VDD.n85 9.3
R934 VDD.n94 VDD.n93 9.3
R935 VDD.n103 VDD.n102 9.3
R936 VDD.n102 VDD.n101 9.3
R937 VDD.n105 VDD.n104 9.3
R938 VDD.n114 VDD.n113 9.3
R939 VDD.n113 VDD.n112 9.3
R940 VDD.n116 VDD.n115 9.3
R941 VDD.n125 VDD.n124 9.3
R942 VDD.n124 VDD.n123 9.3
R943 VDD.n127 VDD.n126 9.3
R944 VDD.n136 VDD.n135 9.3
R945 VDD.n135 VDD.n134 9.3
R946 VDD.n138 VDD.n137 9.3
R947 VDD.n147 VDD.n146 9.3
R948 VDD.n146 VDD.n145 9.3
R949 VDD.n149 VDD.n148 9.3
R950 VDD.n158 VDD.n157 9.3
R951 VDD.n157 VDD.n156 9.3
R952 VDD.n160 VDD.n159 9.3
R953 VDD.n169 VDD.n168 9.3
R954 VDD.n168 VDD.n167 9.3
R955 VDD.n171 VDD.n170 9.3
R956 VDD.n175 VDD.n174 9.3
R957 VDD.n182 VDD.n181 8.679
R958 VDD.n15 VDD.n14 8.679
R959 VDD.n229 VDD.n228 8.422
R960 VDD.n289 VDD.n288 8.422
R961 VDD.n62 VDD.n61 8.422
R962 VDD.n122 VDD.n121 8.422
R963 VDD.n260 VDD.n259 6.787
R964 VDD.n93 VDD.n92 6.787
R965 VDD.n240 VDD.n239 5.147
R966 VDD.n278 VDD.n277 5.147
R967 VDD.n73 VDD.n72 5.147
R968 VDD.n111 VDD.n110 5.147
R969 VDD.n253 VDD.n249 3.103
R970 VDD.n269 VDD.n265 3.103
R971 VDD.n86 VDD.n82 3.103
R972 VDD.n102 VDD.n98 3.103
R973 VDD.n242 VDD.n238 2.715
R974 VDD.n280 VDD.n276 2.715
R975 VDD.n75 VDD.n71 2.715
R976 VDD.n113 VDD.n109 2.715
R977 VDD.n188 VDD.n182 2.611
R978 VDD.n21 VDD.n15 2.611
R979 VDD.n331 VDD.n330 2.521
R980 VDD.n164 VDD.n163 2.521
R981 VDD.n231 VDD.n227 2.327
R982 VDD.n291 VDD.n287 2.327
R983 VDD.n64 VDD.n60 2.327
R984 VDD.n124 VDD.n120 2.327
R985 VDD.n194 VDD.n193 2.133
R986 VDD.n320 VDD.n319 2.133
R987 VDD.n27 VDD.n26 2.133
R988 VDD.n153 VDD.n152 2.133
R989 VDD.n220 VDD.n216 1.939
R990 VDD.n302 VDD.n298 1.939
R991 VDD.n53 VDD.n49 1.939
R992 VDD.n135 VDD.n131 1.939
R993 VDD.n251 VDD.n250 1.748
R994 VDD.n267 VDD.n266 1.748
R995 VDD.n84 VDD.n83 1.748
R996 VDD.n100 VDD.n99 1.748
R997 VDD.n205 VDD.n204 1.745
R998 VDD.n309 VDD.n308 1.745
R999 VDD.n38 VDD.n37 1.745
R1000 VDD.n142 VDD.n141 1.745
R1001 VDD.n209 VDD.n205 1.551
R1002 VDD.n313 VDD.n309 1.551
R1003 VDD.n42 VDD.n38 1.551
R1004 VDD.n146 VDD.n142 1.551
R1005 VDD.n216 VDD.n215 1.357
R1006 VDD.n298 VDD.n297 1.357
R1007 VDD.n49 VDD.n48 1.357
R1008 VDD.n131 VDD.n130 1.357
R1009 VDD.n198 VDD.n194 1.163
R1010 VDD.n324 VDD.n320 1.163
R1011 VDD.n31 VDD.n27 1.163
R1012 VDD.n157 VDD.n153 1.163
R1013 VDD.n227 VDD.n226 0.969
R1014 VDD.n287 VDD.n286 0.969
R1015 VDD.n60 VDD.n59 0.969
R1016 VDD.n120 VDD.n119 0.969
R1017 VDD.n187 VDD.n183 0.775
R1018 VDD.n335 VDD.n331 0.775
R1019 VDD.n20 VDD.n16 0.775
R1020 VDD.n168 VDD.n164 0.775
R1021 VDD.n238 VDD.n237 0.581
R1022 VDD.n276 VDD.n275 0.581
R1023 VDD.n71 VDD.n70 0.581
R1024 VDD.n109 VDD.n108 0.581
R1025 VDD.n176 VDD.n175 0.38
R1026 VDD.n343 VDD.n342 0.361
R1027 VDD.n249 VDD.n248 0.193
R1028 VDD.n265 VDD.n264 0.193
R1029 VDD.n82 VDD.n81 0.193
R1030 VDD.n98 VDD.n97 0.193
R1031 VDD.n261 VDD.n258 0.132
R1032 VDD.n94 VDD.n91 0.132
R1033 VDD.n177 VDD.n176 0.121
R1034 VDD.n199 VDD.n192 0.1
R1035 VDD.n210 VDD.n203 0.1
R1036 VDD.n221 VDD.n214 0.1
R1037 VDD.n232 VDD.n225 0.1
R1038 VDD.n243 VDD.n236 0.1
R1039 VDD.n254 VDD.n247 0.1
R1040 VDD.n272 VDD.n270 0.1
R1041 VDD.n283 VDD.n281 0.1
R1042 VDD.n294 VDD.n292 0.1
R1043 VDD.n305 VDD.n303 0.1
R1044 VDD.n316 VDD.n314 0.1
R1045 VDD.n327 VDD.n325 0.1
R1046 VDD.n338 VDD.n336 0.1
R1047 VDD.n32 VDD.n25 0.1
R1048 VDD.n43 VDD.n36 0.1
R1049 VDD.n54 VDD.n47 0.1
R1050 VDD.n65 VDD.n58 0.1
R1051 VDD.n76 VDD.n69 0.1
R1052 VDD.n87 VDD.n80 0.1
R1053 VDD.n105 VDD.n103 0.1
R1054 VDD.n116 VDD.n114 0.1
R1055 VDD.n127 VDD.n125 0.1
R1056 VDD.n138 VDD.n136 0.1
R1057 VDD.n149 VDD.n147 0.1
R1058 VDD.n160 VDD.n158 0.1
R1059 VDD.n171 VDD.n169 0.1
R1060 VDD.n4 VDD.n2 0.089
R1061 VDD.n352 VDD.n351 0.068
R1062 VDD.n348 VDD.n347 0.06
R1063 VDD.n344 VDD.n343 0.058
R1064 VDD.n350 VDD.n349 0.05
R1065 VDD.n349 VDD.n348 0.043
R1066 VDD.n346 VDD.n345 0.039
R1067 VDD.n345 VDD.n344 0.039
R1068 VDD.n351 VDD.n346 0.03
R1069 VDD.n256 VDD.n254 0.03
R1070 VDD.n270 VDD.n263 0.03
R1071 VDD.n89 VDD.n87 0.03
R1072 VDD.n103 VDD.n96 0.03
R1073 VDD.n8 VDD.n7 0.029
R1074 VDD.n12 VDD.n10 0.029
R1075 VDD.n340 VDD.n338 0.028
R1076 VDD.n173 VDD.n171 0.028
R1077 VDD.n245 VDD.n243 0.026
R1078 VDD.n281 VDD.n274 0.026
R1079 VDD.n78 VDD.n76 0.026
R1080 VDD.n114 VDD.n107 0.026
R1081 VDD.n192 VDD.n190 0.024
R1082 VDD.n329 VDD.n327 0.024
R1083 VDD.n25 VDD.n23 0.024
R1084 VDD.n162 VDD.n160 0.024
R1085 VDD.n234 VDD.n232 0.022
R1086 VDD.n292 VDD.n285 0.022
R1087 VDD.n67 VDD.n65 0.022
R1088 VDD.n125 VDD.n118 0.022
R1089 VDD.n203 VDD.n201 0.02
R1090 VDD.n318 VDD.n316 0.02
R1091 VDD.n36 VDD.n34 0.02
R1092 VDD.n151 VDD.n149 0.02
R1093 VDD VDD.n179 0.019
R1094 VDD.n223 VDD.n221 0.018
R1095 VDD.n303 VDD.n296 0.018
R1096 VDD.n56 VDD.n54 0.018
R1097 VDD.n136 VDD.n129 0.018
R1098 VDD.n214 VDD.n212 0.017
R1099 VDD.n307 VDD.n305 0.017
R1100 VDD.n47 VDD.n45 0.017
R1101 VDD.n140 VDD.n138 0.017
R1102 VDD.n351 VDD.n350 0.016
R1103 VDD.n212 VDD.n210 0.015
R1104 VDD.n314 VDD.n307 0.015
R1105 VDD.n45 VDD.n43 0.015
R1106 VDD.n147 VDD.n140 0.015
R1107 VDD.n1 VDD.n0 0.014
R1108 VDD.n355 VDD.n354 0.014
R1109 VDD.n225 VDD.n223 0.013
R1110 VDD.n296 VDD.n294 0.013
R1111 VDD.n58 VDD.n56 0.013
R1112 VDD.n129 VDD.n127 0.013
R1113 VDD.n178 VDD.n177 0.012
R1114 VDD.n6 VDD.n5 0.012
R1115 VDD.n201 VDD.n199 0.011
R1116 VDD.n325 VDD.n318 0.011
R1117 VDD.n34 VDD.n32 0.011
R1118 VDD.n158 VDD.n151 0.011
R1119 VDD VDD.n356 0.009
R1120 VDD.n236 VDD.n234 0.009
R1121 VDD.n285 VDD.n283 0.009
R1122 VDD.n69 VDD.n67 0.009
R1123 VDD.n118 VDD.n116 0.009
R1124 VDD.n190 VDD.n188 0.007
R1125 VDD.n336 VDD.n329 0.007
R1126 VDD.n23 VDD.n21 0.007
R1127 VDD.n169 VDD.n162 0.007
R1128 VDD.n247 VDD.n245 0.005
R1129 VDD.n274 VDD.n272 0.005
R1130 VDD.n80 VDD.n78 0.005
R1131 VDD.n107 VDD.n105 0.005
R1132 VDD.n179 VDD.n178 0.005
R1133 VDD.n7 VDD.n6 0.005
R1134 VDD.n342 VDD.n340 0.003
R1135 VDD.n175 VDD.n173 0.003
R1136 VDD.n10 VDD.n9 0.003
R1137 VDD.n353 VDD.n352 0.003
R1138 VDD.n4 VDD.n3 0.001
R1139 VDD.n12 VDD.n11 0.001
R1140 VDD.n258 VDD.n256 0.001
R1141 VDD.n263 VDD.n261 0.001
R1142 VDD.n91 VDD.n89 0.001
R1143 VDD.n96 VDD.n94 0.001
R1144 VDD.n178 VDD.n12 0.001
R1145 VDD.n6 VDD.n4 0.001
R1146 VDD.n356 VDD.n355 0.001
R1147 VDD.n356 VDD.n353 0.001
R1148 VDD.n8 VDD.n1 0.001
R1149 VDD.n9 VDD.n8 0.001
R1150 net1_ff1.n13 net1_ff1.n10 9.3
R1151 net1_ff1.n5 net1_ff1.n3 9.3
R1152 net1_ff1.n24 net1_ff1.n21 9.3
R1153 net1_ff1.n16 net1_ff1.n14 9.3
R1154 net1_ff1.n35 net1_ff1.n32 9.3
R1155 net1_ff1.n30 net1_ff1.n28 9.3
R1156 net1_ff1.n41 net1_ff1.n39 9.3
R1157 net1_ff1.n41 net1_ff1.n40 9.3
R1158 net1_ff1.n59 net1_ff1.n57 9.3
R1159 net1_ff1.n59 net1_ff1.n58 9.3
R1160 net1_ff1.n70 net1_ff1.n68 9.3
R1161 net1_ff1.n70 net1_ff1.n69 9.3
R1162 net1_ff1.n81 net1_ff1.n79 9.3
R1163 net1_ff1.n81 net1_ff1.n80 9.3
R1164 net1_ff1.n27 net1_ff1.n25 9.3
R1165 net1_ff1.n35 net1_ff1.n34 9.3
R1166 net1_ff1.n38 net1_ff1.n36 9.3
R1167 net1_ff1.n44 net1_ff1.n42 9.3
R1168 net1_ff1.n56 net1_ff1.n53 9.3
R1169 net1_ff1.n62 net1_ff1.n60 9.3
R1170 net1_ff1.n67 net1_ff1.n64 9.3
R1171 net1_ff1.n73 net1_ff1.n71 9.3
R1172 net1_ff1.n78 net1_ff1.n75 9.3
R1173 net1_ff1.n84 net1_ff1.n82 9.3
R1174 net1_ff1.n89 net1_ff1.n86 9.3
R1175 net1_ff1.n95 net1_ff1.n93 9.3
R1176 net1_ff1.n92 net1_ff1.n90 9.3
R1177 net1_ff1.n38 net1_ff1.n37 9.3
R1178 net1_ff1.n44 net1_ff1.n43 9.3
R1179 net1_ff1.n56 net1_ff1.n55 9.3
R1180 net1_ff1.n62 net1_ff1.n61 9.3
R1181 net1_ff1.n67 net1_ff1.n66 9.3
R1182 net1_ff1.n73 net1_ff1.n72 9.3
R1183 net1_ff1.n78 net1_ff1.n77 9.3
R1184 net1_ff1.n84 net1_ff1.n83 9.3
R1185 net1_ff1.n89 net1_ff1.n88 9.3
R1186 net1_ff1.n95 net1_ff1.n94 9.3
R1187 net1_ff1.n92 net1_ff1.n91 9.3
R1188 net1_ff1.n30 net1_ff1.n29 9.3
R1189 net1_ff1.n27 net1_ff1.n26 9.3
R1190 net1_ff1.n24 net1_ff1.n23 9.3
R1191 net1_ff1.n19 net1_ff1.n17 9.3
R1192 net1_ff1.n19 net1_ff1.n18 9.3
R1193 net1_ff1.n16 net1_ff1.n15 9.3
R1194 net1_ff1.n13 net1_ff1.n12 9.3
R1195 net1_ff1.n8 net1_ff1.n6 9.3
R1196 net1_ff1.n8 net1_ff1.n7 9.3
R1197 net1_ff1.n5 net1_ff1.n4 9.3
R1198 net1_ff1.n48 net1_ff1.t1 7.141
R1199 net1_ff1.n45 net1_ff1.t0 7.141
R1200 net1_ff1.n47 net1_ff1.n46 5.418
R1201 net1_ff1.n50 net1_ff1.n49 5.418
R1202 net1_ff1.n2 net1_ff1.n0 4.728
R1203 net1_ff1.n98 net1_ff1.n96 4.728
R1204 net1_ff1.n98 net1_ff1.n97 4.728
R1205 net1_ff1.n2 net1_ff1.n1 4.727
R1206 net1_ff1.n51 net1_ff1.n47 4.65
R1207 net1_ff1.n51 net1_ff1.n50 4.65
R1208 net1_ff1.n46 net1_ff1.n45 1.844
R1209 net1_ff1.n49 net1_ff1.n48 1.844
R1210 net1_ff1.n12 net1_ff1.n11 0.144
R1211 net1_ff1.n10 net1_ff1.n9 0.144
R1212 net1_ff1.n86 net1_ff1.n85 0.144
R1213 net1_ff1.n88 net1_ff1.n87 0.144
R1214 net1_ff1.n23 net1_ff1.n22 0.133
R1215 net1_ff1.n77 net1_ff1.n76 0.133
R1216 net1_ff1.n21 net1_ff1.n20 0.133
R1217 net1_ff1.n75 net1_ff1.n74 0.132
R1218 net1_ff1.n34 net1_ff1.n33 0.121
R1219 net1_ff1.n32 net1_ff1.n31 0.121
R1220 net1_ff1.n64 net1_ff1.n63 0.121
R1221 net1_ff1.n66 net1_ff1.n65 0.121
R1222 net1_ff1.n55 net1_ff1.n54 0.11
R1223 net1_ff1.n53 net1_ff1.n52 0.109
R1224 net1_ff1.n51 net1_ff1.n44 0.036
R1225 net1_ff1.n56 net1_ff1.n51 0.036
R1226 net1_ff1.n5 net1_ff1.n2 0.029
R1227 net1_ff1 net1_ff1.n98 0.028
R1228 net1_ff1.n16 net1_ff1.n13 0.027
R1229 net1_ff1.n27 net1_ff1.n24 0.027
R1230 net1_ff1.n38 net1_ff1.n35 0.027
R1231 net1_ff1.n67 net1_ff1.n62 0.027
R1232 net1_ff1.n78 net1_ff1.n73 0.027
R1233 net1_ff1.n89 net1_ff1.n84 0.027
R1234 net1_ff1.n41 net1_ff1.n38 0.007
R1235 net1_ff1.n62 net1_ff1.n59 0.007
R1236 net1_ff1.n30 net1_ff1.n27 0.006
R1237 net1_ff1.n73 net1_ff1.n70 0.006
R1238 net1_ff1.n19 net1_ff1.n16 0.005
R1239 net1_ff1.n84 net1_ff1.n81 0.005
R1240 net1_ff1.n8 net1_ff1.n5 0.004
R1241 net1_ff1.n13 net1_ff1.n8 0.004
R1242 net1_ff1.n92 net1_ff1.n89 0.004
R1243 net1_ff1.n95 net1_ff1.n92 0.004
R1244 net1_ff1.n24 net1_ff1.n19 0.003
R1245 net1_ff1.n81 net1_ff1.n78 0.003
R1246 net1_ff1.n35 net1_ff1.n30 0.002
R1247 net1_ff1.n70 net1_ff1.n67 0.002
R1248 net1_ff1.n44 net1_ff1.n41 0.001
R1249 net1_ff1.n59 net1_ff1.n56 0.001
R1250 net1_ff1 net1_ff1.n95 0.001
R1251 modo.n257 modo.t2 1037.29
R1252 modo modo.t3 796.318
R1253 modo.n30 modo.n29 92.5
R1254 modo.n46 modo.n45 92.5
R1255 modo.n45 modo.t1 70.344
R1256 modo.n8 modo.n7 31.034
R1257 modo.n65 modo.n64 31.034
R1258 modo.n113 modo.n112 9.3
R1259 modo.n190 modo.n189 9.3
R1260 modo.n15 modo.n14 9.3
R1261 modo.n66 modo.n65 9.3
R1262 modo.n9 modo.n8 9.3
R1263 modo.n77 modo.n76 9.3
R1264 modo.n229 modo.n228 9.154
R1265 modo.n257 modo.n256 8.715
R1266 modo.n31 modo.n30 8.282
R1267 modo.n47 modo.n46 8.282
R1268 modo.n228 modo.t0 7.141
R1269 modo.n149 modo.n148 7.033
R1270 modo.n92 modo.n91 7.033
R1271 modo.n9 modo.n5 5.647
R1272 modo.n66 modo.n62 5.647
R1273 modo.n230 modo.n229 4.65
R1274 modo.n44 modo.n43 4.65
R1275 modo.n176 modo.n175 4.5
R1276 modo.n196 modo.n195 4.5
R1277 modo.n209 modo.n208 4.5
R1278 modo.n216 modo.n213 4.5
R1279 modo.n225 modo.n224 4.5
R1280 modo.n231 modo.n227 4.5
R1281 modo.n100 modo.n97 4.5
R1282 modo.n107 modo.n106 4.5
R1283 modo.n119 modo.n118 4.5
R1284 modo.n129 modo.n128 4.5
R1285 modo.n139 modo.n138 4.5
R1286 modo.n163 modo.n162 4.5
R1287 modo.n83 modo.n81 4.5
R1288 modo.n70 modo.n67 4.5
R1289 modo.n57 modo.n55 4.5
R1290 modo.n32 modo.n31 4.5
R1291 modo.n39 modo.n38 4.5
R1292 modo.n48 modo.n47 4.5
R1293 modo.n12 modo.n11 4.5
R1294 modo.n20 modo.n19 4.5
R1295 modo.n128 modo.n125 4.141
R1296 modo.n162 modo.n161 4.141
R1297 modo.n7 modo.n6 4.137
R1298 modo.n64 modo.n63 4.137
R1299 modo.n118 modo.n115 3.764
R1300 modo.n208 modo.n206 3.764
R1301 modo.n19 modo.n17 3.764
R1302 modo.n67 modo.n60 3.764
R1303 modo.n138 modo.n135 3.388
R1304 modo.n106 modo.n105 3.388
R1305 modo.n195 modo.n194 3.388
R1306 modo.n175 modo.n174 3.388
R1307 modo.n11 modo.n10 3.388
R1308 modo.n81 modo.n80 3.388
R1309 modo.n138 modo.n137 3.011
R1310 modo.n106 modo.n103 3.011
R1311 modo.n97 modo.n95 3.011
R1312 modo.n189 modo.n188 3.011
R1313 modo.n195 modo.n193 3.011
R1314 modo.n175 modo.n173 3.011
R1315 modo.n11 modo.n9 3.011
R1316 modo.n31 modo.n28 3.011
R1317 modo.n81 modo.n79 3.011
R1318 modo.n118 modo.n117 2.635
R1319 modo.n112 modo.n111 2.635
R1320 modo.n213 modo.n212 2.635
R1321 modo.n208 modo.n207 2.635
R1322 modo.n19 modo.n18 2.635
R1323 modo.n55 modo.n54 2.635
R1324 modo.n67 modo.n66 2.635
R1325 modo.n128 modo.n127 2.258
R1326 modo.n162 modo.n160 2.258
R1327 modo.n25 modo.n0 1.754
R1328 modo.n179 modo.n150 1.754
R1329 modo.n25 modo.n24 1.705
R1330 modo.n42 modo.n41 1.705
R1331 modo.n72 modo.n71 1.705
R1332 modo.n86 modo.n85 1.705
R1333 modo.n255 modo.n144 1.705
R1334 modo.n199 modo.n198 1.705
R1335 modo.n219 modo.n218 1.705
R1336 modo.n248 modo.n247 1.705
R1337 modo.n254 modo.n253 1.705
R1338 modo.n242 modo.n241 1.705
R1339 modo.n236 modo.n235 1.705
R1340 modo.n185 modo.n184 1.705
R1341 modo.n179 modo.n178 1.705
R1342 modo.n213 modo.n211 1.505
R1343 modo.n197 modo.n196 1.5
R1344 modo.n210 modo.n209 1.5
R1345 modo.n217 modo.n216 1.5
R1346 modo.n226 modo.n225 1.5
R1347 modo.n232 modo.n231 1.5
R1348 modo.n84 modo.n83 1.5
R1349 modo.n71 modo.n70 1.5
R1350 modo.n33 modo.n32 1.5
R1351 modo.n58 modo.n57 1.5
R1352 modo.n40 modo.n39 1.5
R1353 modo.n49 modo.n48 1.5
R1354 modo.n24 modo.n12 1.5
R1355 modo.n21 modo.n20 1.5
R1356 modo.n256 modo.n255 1.268
R1357 modo modo.n257 1.256
R1358 modo.n97 modo.n96 1.129
R1359 modo.n150 modo.n149 1.127
R1360 modo.n144 modo.n92 1.127
R1361 modo.n140 modo.n139 1.125
R1362 modo.n177 modo.n176 1.125
R1363 modo.n5 modo.n4 0.752
R1364 modo.n62 modo.n61 0.752
R1365 modo.n256 modo.n86 0.709
R1366 modo.n91 modo.n90 0.155
R1367 modo.n148 modo.n147 0.155
R1368 modo.n137 modo.n136 0.144
R1369 modo.n173 modo.n172 0.144
R1370 modo.n127 modo.n126 0.133
R1371 modo.n160 modo.n159 0.132
R1372 modo.n133 modo.n132 0.053
R1373 modo.n123 modo.n122 0.053
R1374 modo.n113 modo.n110 0.053
R1375 modo.n157 modo.n156 0.053
R1376 modo.n167 modo.n166 0.053
R1377 modo.n170 modo.n169 0.053
R1378 modo.n77 modo.n75 0.053
R1379 modo.n42 modo.n25 0.049
R1380 modo.n72 modo.n42 0.049
R1381 modo.n86 modo.n72 0.049
R1382 modo.n255 modo.n254 0.049
R1383 modo.n254 modo.n248 0.049
R1384 modo.n248 modo.n242 0.049
R1385 modo.n242 modo.n236 0.049
R1386 modo.n236 modo.n219 0.049
R1387 modo.n219 modo.n199 0.049
R1388 modo.n199 modo.n185 0.049
R1389 modo.n185 modo.n179 0.049
R1390 modo.n39 modo.n37 0.045
R1391 modo.n57 modo.n53 0.045
R1392 modo.n100 modo.n99 0.043
R1393 modo.n225 modo.n223 0.043
R1394 modo.n88 modo.n87 0.034
R1395 modo.n166 modo.n165 0.032
R1396 modo.n134 modo.n133 0.03
R1397 modo.n132 modo.n131 0.03
R1398 modo.n156 modo.n155 0.03
R1399 modo.n22 modo.n21 0.03
R1400 modo.n84 modo.n74 0.03
R1401 modo.n122 modo.n121 0.028
R1402 modo.n168 modo.n167 0.028
R1403 modo.n171 modo.n170 0.028
R1404 modo.n94 modo.n93 0.025
R1405 modo.n124 modo.n123 0.025
R1406 modo.n48 modo.n44 0.025
R1407 modo.n117 modo.n116 0.024
R1408 modo.n193 modo.n192 0.024
R1409 modo.n231 modo.n230 0.023
R1410 modo.n158 modo.n157 0.023
R1411 modo.n120 modo.n119 0.021
R1412 modo.n114 modo.n113 0.021
R1413 modo.n203 modo.n202 0.021
R1414 modo.n20 modo.n13 0.021
R1415 modo.n16 modo.n15 0.021
R1416 modo.n70 modo.n59 0.021
R1417 modo.n139 modo.n94 0.019
R1418 modo.n110 modo.n109 0.019
R1419 modo.n109 modo.n108 0.019
R1420 modo.n107 modo.n102 0.019
R1421 modo.n204 modo.n203 0.019
R1422 modo.n191 modo.n190 0.019
R1423 modo.n176 modo.n171 0.019
R1424 modo.n2 modo.n1 0.019
R1425 modo.n3 modo.n2 0.019
R1426 modo.n69 modo.n68 0.019
R1427 modo.n78 modo.n77 0.019
R1428 modo.n83 modo.n82 0.019
R1429 modo.n92 modo.n89 0.019
R1430 modo.n149 modo.n146 0.019
R1431 modo.n198 modo.n197 0.018
R1432 modo.n139 modo.n134 0.017
R1433 modo.n130 modo.n129 0.017
R1434 modo.n108 modo.n107 0.017
R1435 modo.n101 modo.n100 0.017
R1436 modo.n196 modo.n191 0.017
R1437 modo.n164 modo.n163 0.017
R1438 modo.n176 modo.n168 0.017
R1439 modo.n12 modo.n3 0.017
R1440 modo.n32 modo.n27 0.017
R1441 modo.n83 modo.n78 0.017
R1442 modo.n142 modo.n141 0.016
R1443 modo.n252 modo.n251 0.016
R1444 modo.n246 modo.n245 0.016
R1445 modo.n181 modo.n180 0.016
R1446 modo.n153 modo.n152 0.016
R1447 modo.n71 modo.n58 0.016
R1448 modo.n119 modo.n114 0.015
R1449 modo.n216 modo.n215 0.015
R1450 modo.n209 modo.n204 0.015
R1451 modo.n238 modo.n237 0.015
R1452 modo.n232 modo.n226 0.015
R1453 modo.n217 modo.n210 0.015
R1454 modo.n20 modo.n16 0.015
R1455 modo.n57 modo.n56 0.015
R1456 modo.n70 modo.n69 0.015
R1457 modo.n40 modo.n35 0.015
R1458 modo.n58 modo.n51 0.015
R1459 modo.n177 modo.n153 0.014
R1460 modo.n34 modo.n33 0.014
R1461 modo.n50 modo.n49 0.014
R1462 modo.n141 modo.n140 0.013
R1463 modo.n233 modo.n232 0.013
R1464 modo.n226 modo.n221 0.013
R1465 modo.n105 modo.n104 0.012
R1466 modo.n206 modo.n205 0.012
R1467 modo.n129 modo.n124 0.012
R1468 modo.n102 modo.n101 0.012
R1469 modo.n215 modo.n214 0.012
R1470 modo.n163 modo.n158 0.012
R1471 modo.n27 modo.n26 0.012
R1472 modo.n143 modo.n142 0.011
R1473 modo.n251 modo.n250 0.011
R1474 modo.n239 modo.n238 0.011
R1475 modo.n218 modo.n217 0.011
R1476 modo.n182 modo.n181 0.011
R1477 modo.n152 modo.n151 0.011
R1478 modo.n24 modo.n23 0.011
R1479 modo.n210 modo.n201 0.01
R1480 modo.n184 modo.n183 0.01
R1481 modo.n253 modo.n252 0.009
R1482 modo.n241 modo.n240 0.009
R1483 modo.n187 modo.n186 0.009
R1484 modo.n99 modo.n98 0.008
R1485 modo.n223 modo.n222 0.008
R1486 modo.n245 modo.n244 0.008
R1487 modo.n244 modo.n243 0.008
R1488 modo.n37 modo.n36 0.008
R1489 modo.n53 modo.n52 0.008
R1490 modo.n85 modo.n84 0.008
R1491 modo.n197 modo.n187 0.007
R1492 modo.n41 modo.n40 0.007
R1493 modo.n74 modo.n73 0.007
R1494 modo.n131 modo.n130 0.006
R1495 modo.n121 modo.n120 0.006
R1496 modo.n155 modo.n154 0.006
R1497 modo.n165 modo.n164 0.006
R1498 modo.n201 modo.n200 0.006
R1499 modo.n23 modo.n22 0.006
R1500 modo.n144 modo.n143 0.005
R1501 modo.n250 modo.n249 0.005
R1502 modo.n240 modo.n239 0.005
R1503 modo.n183 modo.n182 0.005
R1504 modo.n178 modo.n177 0.005
R1505 modo.n89 modo.n88 0.004
R1506 modo.n146 modo.n145 0.004
R1507 modo.n235 modo.n234 0.002
R1508 modo.n234 modo.n233 0.002
R1509 modo.n221 modo.n220 0.002
R1510 modo.n35 modo.n34 0.002
R1511 modo.n51 modo.n50 0.002
R1512 modo.n247 modo.n246 0.001
R1513 net2_nand3.n1 net2_nand3.n0 13.361
R1514 net2_nand3.n86 net2_nand3.n85 13.361
R1515 net2_nand3.n11 net2_nand3.n9 9.3
R1516 net2_nand3.n5 net2_nand3.n3 9.3
R1517 net2_nand3.n16 net2_nand3.n13 9.3
R1518 net2_nand3.n140 net2_nand3.n132 9.3
R1519 net2_nand3.n140 net2_nand3.n139 9.3
R1520 net2_nand3.n22 net2_nand3.n20 9.3
R1521 net2_nand3.n33 net2_nand3.n31 9.3
R1522 net2_nand3.n30 net2_nand3.n28 9.3
R1523 net2_nand3.n41 net2_nand3.n39 9.3
R1524 net2_nand3.n41 net2_nand3.n40 9.3
R1525 net2_nand3.n52 net2_nand3.n50 9.3
R1526 net2_nand3.n52 net2_nand3.n51 9.3
R1527 net2_nand3.n63 net2_nand3.n61 9.3
R1528 net2_nand3.n63 net2_nand3.n62 9.3
R1529 net2_nand3.n74 net2_nand3.n72 9.3
R1530 net2_nand3.n74 net2_nand3.n73 9.3
R1531 net2_nand3.n98 net2_nand3.n96 9.3
R1532 net2_nand3.n98 net2_nand3.n97 9.3
R1533 net2_nand3.n109 net2_nand3.n107 9.3
R1534 net2_nand3.n109 net2_nand3.n108 9.3
R1535 net2_nand3.n167 net2_nand3.n116 9.3
R1536 net2_nand3.n167 net2_nand3.n166 9.3
R1537 net2_nand3.n159 net2_nand3.n121 9.3
R1538 net2_nand3.n159 net2_nand3.n158 9.3
R1539 net2_nand3.n152 net2_nand3.n125 9.3
R1540 net2_nand3.n152 net2_nand3.n151 9.3
R1541 net2_nand3.n27 net2_nand3.n24 9.3
R1542 net2_nand3.n33 net2_nand3.n32 9.3
R1543 net2_nand3.n38 net2_nand3.n35 9.3
R1544 net2_nand3.n44 net2_nand3.n42 9.3
R1545 net2_nand3.n49 net2_nand3.n46 9.3
R1546 net2_nand3.n55 net2_nand3.n53 9.3
R1547 net2_nand3.n60 net2_nand3.n57 9.3
R1548 net2_nand3.n66 net2_nand3.n64 9.3
R1549 net2_nand3.n71 net2_nand3.n68 9.3
R1550 net2_nand3.n77 net2_nand3.n75 9.3
R1551 net2_nand3.n82 net2_nand3.n79 9.3
R1552 net2_nand3.n92 net2_nand3.n89 9.3
R1553 net2_nand3.n95 net2_nand3.n93 9.3
R1554 net2_nand3.n103 net2_nand3.n100 9.3
R1555 net2_nand3.n106 net2_nand3.n104 9.3
R1556 net2_nand3.n114 net2_nand3.n111 9.3
R1557 net2_nand3 net2_nand3.n168 9.3
R1558 net2_nand3.n165 net2_nand3.n119 9.3
R1559 net2_nand3.n161 net2_nand3.n120 9.3
R1560 net2_nand3.n157 net2_nand3.n123 9.3
R1561 net2_nand3.n154 net2_nand3.n124 9.3
R1562 net2_nand3.n150 net2_nand3.n127 9.3
R1563 net2_nand3.n147 net2_nand3.n128 9.3
R1564 net2_nand3.n143 net2_nand3.n131 9.3
R1565 net2_nand3.n145 net2_nand3.n129 9.3
R1566 net2_nand3.n38 net2_nand3.n37 9.3
R1567 net2_nand3.n44 net2_nand3.n43 9.3
R1568 net2_nand3.n49 net2_nand3.n48 9.3
R1569 net2_nand3.n55 net2_nand3.n54 9.3
R1570 net2_nand3.n60 net2_nand3.n59 9.3
R1571 net2_nand3.n66 net2_nand3.n65 9.3
R1572 net2_nand3.n71 net2_nand3.n70 9.3
R1573 net2_nand3.n77 net2_nand3.n76 9.3
R1574 net2_nand3.n82 net2_nand3.n81 9.3
R1575 net2_nand3.n92 net2_nand3.n91 9.3
R1576 net2_nand3.n95 net2_nand3.n94 9.3
R1577 net2_nand3.n103 net2_nand3.n102 9.3
R1578 net2_nand3.n106 net2_nand3.n105 9.3
R1579 net2_nand3.n114 net2_nand3.n113 9.3
R1580 net2_nand3 net2_nand3.n115 9.3
R1581 net2_nand3.n165 net2_nand3.n164 9.3
R1582 net2_nand3.n161 net2_nand3.n160 9.3
R1583 net2_nand3.n157 net2_nand3.n156 9.3
R1584 net2_nand3.n154 net2_nand3.n153 9.3
R1585 net2_nand3.n150 net2_nand3.n149 9.3
R1586 net2_nand3.n147 net2_nand3.n146 9.3
R1587 net2_nand3.n143 net2_nand3.n142 9.3
R1588 net2_nand3.n145 net2_nand3.n144 9.3
R1589 net2_nand3.n30 net2_nand3.n29 9.3
R1590 net2_nand3.n27 net2_nand3.n26 9.3
R1591 net2_nand3.n22 net2_nand3.n21 9.3
R1592 net2_nand3.n19 net2_nand3.n17 9.3
R1593 net2_nand3.n19 net2_nand3.n18 9.3
R1594 net2_nand3.n16 net2_nand3.n15 9.3
R1595 net2_nand3.n136 net2_nand3.n134 9.3
R1596 net2_nand3.n138 net2_nand3.n133 9.3
R1597 net2_nand3.n138 net2_nand3.n137 9.3
R1598 net2_nand3.n136 net2_nand3.n135 9.3
R1599 net2_nand3.n11 net2_nand3.n10 9.3
R1600 net2_nand3.n8 net2_nand3.n6 9.3
R1601 net2_nand3.n8 net2_nand3.n7 9.3
R1602 net2_nand3.n5 net2_nand3.n4 9.3
R1603 net2_nand3.n118 net2_nand3.n117 8.043
R1604 net2_nand3.n163 net2_nand3.n162 8.043
R1605 net2_nand3.n84 net2_nand3.n2 4.558
R1606 net2_nand3.n87 net2_nand3.n1 4.558
R1607 net2_nand3.n84 net2_nand3.n83 4.558
R1608 net2_nand3.n87 net2_nand3.n86 4.558
R1609 net2_nand3.n162 net2_nand3.t1 2.9
R1610 net2_nand3.n117 net2_nand3.t0 2.9
R1611 net2_nand3.n79 net2_nand3.n78 0.536
R1612 net2_nand3.n89 net2_nand3.n88 0.536
R1613 net2_nand3.n81 net2_nand3.n80 0.536
R1614 net2_nand3.n91 net2_nand3.n90 0.536
R1615 net2_nand3.n70 net2_nand3.n69 0.506
R1616 net2_nand3.n102 net2_nand3.n101 0.506
R1617 net2_nand3.n68 net2_nand3.n67 0.506
R1618 net2_nand3.n100 net2_nand3.n99 0.506
R1619 net2_nand3.n57 net2_nand3.n56 0.475
R1620 net2_nand3.n111 net2_nand3.n110 0.475
R1621 net2_nand3.n59 net2_nand3.n58 0.475
R1622 net2_nand3.n113 net2_nand3.n112 0.475
R1623 net2_nand3.n164 net2_nand3.n163 0.445
R1624 net2_nand3.n46 net2_nand3.n45 0.445
R1625 net2_nand3.n119 net2_nand3.n118 0.445
R1626 net2_nand3.n48 net2_nand3.n47 0.445
R1627 net2_nand3.n35 net2_nand3.n34 0.413
R1628 net2_nand3.n123 net2_nand3.n122 0.413
R1629 net2_nand3.n37 net2_nand3.n36 0.413
R1630 net2_nand3.n156 net2_nand3.n155 0.413
R1631 net2_nand3.n26 net2_nand3.n25 0.382
R1632 net2_nand3.n149 net2_nand3.n148 0.382
R1633 net2_nand3.n127 net2_nand3.n126 0.382
R1634 net2_nand3.n24 net2_nand3.n23 0.382
R1635 net2_nand3.n13 net2_nand3.n12 0.349
R1636 net2_nand3.n15 net2_nand3.n14 0.349
R1637 net2_nand3.n131 net2_nand3.n130 0.349
R1638 net2_nand3.n142 net2_nand3.n141 0.349
R1639 net2_nand3.n87 net2_nand3.n84 0.055
R1640 net2_nand3.n16 net2_nand3.n11 0.041
R1641 net2_nand3.n27 net2_nand3.n22 0.041
R1642 net2_nand3.n38 net2_nand3.n33 0.041
R1643 net2_nand3.n49 net2_nand3.n44 0.041
R1644 net2_nand3.n60 net2_nand3.n55 0.041
R1645 net2_nand3.n71 net2_nand3.n66 0.041
R1646 net2_nand3.n82 net2_nand3.n77 0.041
R1647 net2_nand3.n95 net2_nand3.n92 0.041
R1648 net2_nand3.n106 net2_nand3.n103 0.041
R1649 net2_nand3 net2_nand3.n114 0.041
R1650 net2_nand3.n165 net2_nand3.n161 0.041
R1651 net2_nand3.n157 net2_nand3.n154 0.041
R1652 net2_nand3.n150 net2_nand3.n147 0.041
R1653 net2_nand3.n143 net2_nand3.n140 0.041
R1654 net2_nand3.n84 net2_nand3.n82 0.012
R1655 net2_nand3.n92 net2_nand3.n87 0.012
R1656 net2_nand3.n11 net2_nand3.n8 0.011
R1657 net2_nand3.n74 net2_nand3.n71 0.011
R1658 net2_nand3.n103 net2_nand3.n98 0.011
R1659 net2_nand3.n140 net2_nand3.n138 0.011
R1660 net2_nand3.n22 net2_nand3.n19 0.01
R1661 net2_nand3.n147 net2_nand3.n145 0.01
R1662 net2_nand3.n63 net2_nand3.n60 0.009
R1663 net2_nand3.n114 net2_nand3.n109 0.009
R1664 net2_nand3.n33 net2_nand3.n30 0.008
R1665 net2_nand3.n154 net2_nand3.n152 0.008
R1666 net2_nand3.n44 net2_nand3.n41 0.007
R1667 net2_nand3.n52 net2_nand3.n49 0.007
R1668 net2_nand3.n167 net2_nand3.n165 0.007
R1669 net2_nand3.n161 net2_nand3.n159 0.007
R1670 net2_nand3.n41 net2_nand3.n38 0.006
R1671 net2_nand3.n159 net2_nand3.n157 0.006
R1672 net2_nand3.n55 net2_nand3.n52 0.005
R1673 net2_nand3 net2_nand3.n167 0.005
R1674 net2_nand3.n30 net2_nand3.n27 0.004
R1675 net2_nand3.n152 net2_nand3.n150 0.004
R1676 net2_nand3.n19 net2_nand3.n16 0.003
R1677 net2_nand3.n66 net2_nand3.n63 0.003
R1678 net2_nand3.n109 net2_nand3.n106 0.003
R1679 net2_nand3.n145 net2_nand3.n143 0.003
R1680 net2_nand3.n77 net2_nand3.n74 0.002
R1681 net2_nand3.n98 net2_nand3.n95 0.002
R1682 net2_nand3.n8 net2_nand3.n5 0.001
R1683 net2_nand3.n138 net2_nand3.n136 0.001
R1684 GND.t5 GND.t2 3022.52
R1685 GND.t12 GND.t3 3007.96
R1686 GND.n48 GND.t12 2686.73
R1687 GND.n48 GND.t5 1696.78
R1688 GND.n188 GND.n187 589.285
R1689 GND.n164 GND.n163 589.285
R1690 GND.n199 GND.n198 585
R1691 GND.n183 GND.n182 585
R1692 GND.n161 GND.n160 585
R1693 GND.n145 GND.n144 585
R1694 GND.n131 GND.n130 585
R1695 GND.n117 GND.n116 585
R1696 GND.n103 GND.n102 585
R1697 GND.n89 GND.n88 585
R1698 GND.n75 GND.n74 585
R1699 GND.n61 GND.n60 585
R1700 GND.n54 GND.n53 585
R1701 GND.n202 GND.n201 510.714
R1702 GND.n148 GND.n147 510.714
R1703 GND.n134 GND.n133 432.142
R1704 GND.n120 GND.n119 353.571
R1705 GND.n186 GND.n185 292.5
R1706 GND.n159 GND.n158 292.5
R1707 GND.n106 GND.n105 275
R1708 GND.n47 GND.n46 235.714
R1709 GND.n92 GND.n91 196.428
R1710 GND.n189 GND.n186 174.016
R1711 GND.n165 GND.n159 174.016
R1712 GND.n347 GND.t4 124.695
R1713 GND.n284 GND.t0 124.695
R1714 GND.n2 GND.t11 124.695
R1715 GND.n304 GND.t10 124.695
R1716 GND.n324 GND.t9 124.695
R1717 GND.n23 GND.t6 124.688
R1718 GND.n78 GND.n77 117.857
R1719 GND.n346 GND.n345 92.5
R1720 GND.n22 GND.n21 92.5
R1721 GND.n283 GND.n282 92.5
R1722 GND.n1 GND.n0 92.5
R1723 GND.n303 GND.n302 92.5
R1724 GND.n323 GND.n322 92.5
R1725 GND.n48 GND.n47 78.571
R1726 GND.n44 GND.n43 53.678
R1727 GND.n45 GND.n44 52.533
R1728 GND.n275 GND.n274 52.533
R1729 GND.n62 GND.n61 52.533
R1730 GND.n55 GND.n54 52.533
R1731 GND.n189 GND.n184 49.25
R1732 GND.n165 GND.n162 49.25
R1733 GND.n76 GND.n75 45.966
R1734 GND.n203 GND.n200 42.683
R1735 GND.n149 GND.n146 42.683
R1736 GND.n250 GND.n249 39.4
R1737 GND.n90 GND.n89 39.4
R1738 GND.n64 GND.n63 39.285
R1739 GND.n215 GND.n213 36.116
R1740 GND.n135 GND.n132 36.116
R1741 GND.n104 GND.n103 32.833
R1742 GND.n356 GND.n355 31.034
R1743 GND.n32 GND.n31 31.034
R1744 GND.n293 GND.n292 31.034
R1745 GND.n11 GND.n10 31.034
R1746 GND.n313 GND.n312 31.034
R1747 GND.n333 GND.n332 31.034
R1748 GND.n121 GND.n118 29.55
R1749 GND.n226 GND.n225 27.71
R1750 GND.n225 GND.n224 26.266
R1751 GND.n118 GND.n117 26.266
R1752 GND.n240 GND.n238 22.983
R1753 GND.n107 GND.n104 22.983
R1754 GND.n262 GND.n261 22.115
R1755 GND.n263 GND.n262 22.115
R1756 GND.n213 GND.n212 19.7
R1757 GND.n132 GND.n131 19.7
R1758 GND.n93 GND.n90 16.416
R1759 GND.n237 GND.n236 15.969
R1760 GND.n238 GND.n237 15.969
R1761 GND.n251 GND.n250 15.725
R1762 GND.n23 GND.n22 15.433
R1763 GND.n347 GND.n346 15.431
R1764 GND.n284 GND.n283 15.431
R1765 GND.n2 GND.n1 15.431
R1766 GND.n304 GND.n303 15.431
R1767 GND.n324 GND.n323 15.431
R1768 GND.n200 GND.n199 13.133
R1769 GND.n146 GND.n145 13.133
R1770 GND.n265 GND.n263 9.85
R1771 GND.n79 GND.n76 9.85
R1772 GND.n57 GND.n56 9.551
R1773 GND.n50 GND.n49 9.352
R1774 GND.n362 GND.n361 9.3
R1775 GND.n351 GND.n350 9.3
R1776 GND.n349 GND.n348 9.3
R1777 GND.n358 GND.n357 9.3
R1778 GND.n357 GND.n356 9.3
R1779 GND.n360 GND.n359 9.3
R1780 GND.n364 GND.n363 9.3
R1781 GND.n271 GND.n270 9.3
R1782 GND.n258 GND.n257 9.3
R1783 GND.n246 GND.n245 9.3
R1784 GND.n233 GND.n232 9.3
R1785 GND.n221 GND.n220 9.3
R1786 GND.n209 GND.n208 9.3
R1787 GND.n195 GND.n194 9.3
R1788 GND.n179 GND.n178 9.3
R1789 GND.n169 GND.n168 9.3
R1790 GND.n153 GND.n152 9.3
R1791 GND.n139 GND.n138 9.3
R1792 GND.n125 GND.n124 9.3
R1793 GND.n111 GND.n110 9.3
R1794 GND.n97 GND.n96 9.3
R1795 GND.n83 GND.n82 9.3
R1796 GND.n69 GND.n68 9.3
R1797 GND.n269 GND.n268 9.3
R1798 GND.n279 GND.n278 9.3
R1799 GND.n278 GND.n277 9.3
R1800 GND.n256 GND.n255 9.3
R1801 GND.n267 GND.n266 9.3
R1802 GND.n266 GND.n265 9.3
R1803 GND.n244 GND.n243 9.3
R1804 GND.n254 GND.n253 9.3
R1805 GND.n253 GND.n252 9.3
R1806 GND.n231 GND.n230 9.3
R1807 GND.n242 GND.n241 9.3
R1808 GND.n241 GND.n240 9.3
R1809 GND.n219 GND.n218 9.3
R1810 GND.n229 GND.n228 9.3
R1811 GND.n228 GND.n227 9.3
R1812 GND.n207 GND.n206 9.3
R1813 GND.n217 GND.n216 9.3
R1814 GND.n216 GND.n215 9.3
R1815 GND.n215 GND.n214 9.3
R1816 GND.n193 GND.n192 9.3
R1817 GND.n205 GND.n204 9.3
R1818 GND.n204 GND.n203 9.3
R1819 GND.n203 GND.n202 9.3
R1820 GND.n177 GND.n176 9.3
R1821 GND.n191 GND.n190 9.3
R1822 GND.n190 GND.n189 9.3
R1823 GND.n189 GND.n188 9.3
R1824 GND.n171 GND.n170 9.3
R1825 GND.n167 GND.n166 9.3
R1826 GND.n166 GND.n165 9.3
R1827 GND.n165 GND.n164 9.3
R1828 GND.n155 GND.n154 9.3
R1829 GND.n151 GND.n150 9.3
R1830 GND.n150 GND.n149 9.3
R1831 GND.n149 GND.n148 9.3
R1832 GND.n141 GND.n140 9.3
R1833 GND.n137 GND.n136 9.3
R1834 GND.n136 GND.n135 9.3
R1835 GND.n135 GND.n134 9.3
R1836 GND.n127 GND.n126 9.3
R1837 GND.n123 GND.n122 9.3
R1838 GND.n122 GND.n121 9.3
R1839 GND.n121 GND.n120 9.3
R1840 GND.n113 GND.n112 9.3
R1841 GND.n109 GND.n108 9.3
R1842 GND.n108 GND.n107 9.3
R1843 GND.n107 GND.n106 9.3
R1844 GND.n99 GND.n98 9.3
R1845 GND.n95 GND.n94 9.3
R1846 GND.n94 GND.n93 9.3
R1847 GND.n93 GND.n92 9.3
R1848 GND.n85 GND.n84 9.3
R1849 GND.n81 GND.n80 9.3
R1850 GND.n80 GND.n79 9.3
R1851 GND.n79 GND.n78 9.3
R1852 GND.n71 GND.n70 9.3
R1853 GND.n67 GND.n66 9.3
R1854 GND.n66 GND.n65 9.3
R1855 GND.n65 GND.n64 9.3
R1856 GND.n38 GND.n37 9.3
R1857 GND.n27 GND.n26 9.3
R1858 GND.n25 GND.n24 9.3
R1859 GND.n34 GND.n33 9.3
R1860 GND.n33 GND.n32 9.3
R1861 GND.n36 GND.n35 9.3
R1862 GND.n40 GND.n39 9.3
R1863 GND.n299 GND.n298 9.3
R1864 GND.n288 GND.n287 9.3
R1865 GND.n286 GND.n285 9.3
R1866 GND.n295 GND.n294 9.3
R1867 GND.n294 GND.n293 9.3
R1868 GND.n297 GND.n296 9.3
R1869 GND.n301 GND.n300 9.3
R1870 GND.n17 GND.n16 9.3
R1871 GND.n6 GND.n5 9.3
R1872 GND.n4 GND.n3 9.3
R1873 GND.n13 GND.n12 9.3
R1874 GND.n12 GND.n11 9.3
R1875 GND.n15 GND.n14 9.3
R1876 GND.n19 GND.n18 9.3
R1877 GND.n319 GND.n318 9.3
R1878 GND.n308 GND.n307 9.3
R1879 GND.n306 GND.n305 9.3
R1880 GND.n315 GND.n314 9.3
R1881 GND.n314 GND.n313 9.3
R1882 GND.n317 GND.n316 9.3
R1883 GND.n321 GND.n320 9.3
R1884 GND.n339 GND.n338 9.3
R1885 GND.n328 GND.n327 9.3
R1886 GND.n326 GND.n325 9.3
R1887 GND.n335 GND.n334 9.3
R1888 GND.n334 GND.n333 9.3
R1889 GND.n337 GND.n336 9.3
R1890 GND.n341 GND.n340 9.3
R1891 GND.n49 GND.n48 9.105
R1892 GND.n174 GND.n172 7.253
R1893 GND.n174 GND.n173 7.253
R1894 GND.n184 GND.n183 6.566
R1895 GND.n162 GND.n161 6.566
R1896 GND.n357 GND.n353 5.647
R1897 GND.n33 GND.n29 5.647
R1898 GND.n294 GND.n290 5.647
R1899 GND.n12 GND.n8 5.647
R1900 GND.n314 GND.n310 5.647
R1901 GND.n334 GND.n330 5.647
R1902 GND.n343 GND.t7 4.905
R1903 GND.n20 GND.t8 4.829
R1904 GND.n343 GND.t1 4.81
R1905 GND.n175 GND.n174 4.65
R1906 GND.n355 GND.n354 4.137
R1907 GND.n31 GND.n30 4.137
R1908 GND.n292 GND.n291 4.137
R1909 GND.n10 GND.n9 4.137
R1910 GND.n312 GND.n311 4.137
R1911 GND.n332 GND.n331 4.137
R1912 GND.n67 GND.n57 3.638
R1913 GND.n280 GND.n50 3.483
R1914 GND.n42 GND.n41 3.413
R1915 GND.n273 GND.n272 3.413
R1916 GND.n59 GND.n58 3.413
R1917 GND.n52 GND.n51 3.413
R1918 GND.n65 GND.n62 3.283
R1919 GND.n276 GND.n275 3.214
R1920 GND.n49 GND.n45 3.214
R1921 GND.n190 GND.n181 3.2
R1922 GND.n166 GND.n157 3.2
R1923 GND.n56 GND.n55 3.016
R1924 GND.n260 GND.n259 2.986
R1925 GND.n73 GND.n72 2.986
R1926 GND.n204 GND.n197 2.773
R1927 GND.n150 GND.n143 2.773
R1928 GND.n248 GND.n247 2.56
R1929 GND.n87 GND.n86 2.56
R1930 GND.n216 GND.n211 2.346
R1931 GND.n136 GND.n129 2.346
R1932 GND.n235 GND.n234 2.133
R1933 GND.n101 GND.n100 2.133
R1934 GND.n265 GND.n264 2.107
R1935 GND.n240 GND.n239 2.107
R1936 GND.n228 GND.n223 1.92
R1937 GND.n122 GND.n115 1.92
R1938 GND.n223 GND.n222 1.706
R1939 GND.n115 GND.n114 1.706
R1940 GND.n349 GND.n347 1.57
R1941 GND.n286 GND.n284 1.57
R1942 GND.n4 GND.n2 1.57
R1943 GND.n306 GND.n304 1.57
R1944 GND.n326 GND.n324 1.57
R1945 GND.n25 GND.n23 1.553
R1946 GND.n241 GND.n235 1.493
R1947 GND.n108 GND.n101 1.493
R1948 GND.n211 GND.n210 1.28
R1949 GND.n129 GND.n128 1.28
R1950 GND.n253 GND.n248 1.066
R1951 GND.n94 GND.n87 1.066
R1952 GND.n197 GND.n196 0.853
R1953 GND.n143 GND.n142 0.853
R1954 GND.n353 GND.n352 0.752
R1955 GND.n29 GND.n28 0.752
R1956 GND.n290 GND.n289 0.752
R1957 GND.n8 GND.n7 0.752
R1958 GND.n310 GND.n309 0.752
R1959 GND.n330 GND.n329 0.752
R1960 GND.n266 GND.n260 0.64
R1961 GND.n80 GND.n73 0.64
R1962 GND.n366 GND.n301 0.446
R1963 GND.n227 GND.n226 0.441
R1964 GND.n181 GND.n180 0.426
R1965 GND.n157 GND.n156 0.426
R1966 GND.n365 GND.n364 0.42
R1967 GND.n342 GND.n341 0.363
R1968 GND.n20 GND.n19 0.361
R1969 GND.n342 GND.n321 0.323
R1970 GND.n281 GND.n40 0.318
R1971 GND.n281 GND.n280 0.259
R1972 GND.n252 GND.n251 0.25
R1973 GND.n50 GND.n42 0.213
R1974 GND.n278 GND.n273 0.213
R1975 GND.n66 GND.n59 0.213
R1976 GND.n57 GND.n52 0.213
R1977 GND.n280 GND.n279 0.156
R1978 GND.n177 GND.n175 0.145
R1979 GND.n175 GND.n171 0.145
R1980 GND.n360 GND.n358 0.144
R1981 GND.n297 GND.n295 0.144
R1982 GND.n15 GND.n13 0.144
R1983 GND.n317 GND.n315 0.144
R1984 GND.n337 GND.n335 0.144
R1985 GND.n36 GND.n34 0.132
R1986 GND.n269 GND.n267 0.11
R1987 GND.n256 GND.n254 0.11
R1988 GND.n244 GND.n242 0.11
R1989 GND.n231 GND.n229 0.11
R1990 GND.n219 GND.n217 0.11
R1991 GND.n207 GND.n205 0.11
R1992 GND.n193 GND.n191 0.11
R1993 GND.n167 GND.n155 0.11
R1994 GND.n151 GND.n141 0.11
R1995 GND.n137 GND.n127 0.11
R1996 GND.n123 GND.n113 0.11
R1997 GND.n109 GND.n99 0.11
R1998 GND.n95 GND.n85 0.11
R1999 GND.n81 GND.n71 0.11
R2000 GND GND.n20 0.108
R2001 GND.n277 GND.n276 0.052
R2002 GND.n366 GND.n281 0.051
R2003 GND.n365 GND.n344 0.05
R2004 GND.n344 GND.n342 0.048
R2005 GND.n366 GND.n365 0.045
R2006 GND.n358 GND.n351 0.04
R2007 GND.n295 GND.n288 0.04
R2008 GND.n13 GND.n6 0.04
R2009 GND.n315 GND.n308 0.04
R2010 GND.n335 GND.n328 0.04
R2011 GND.n34 GND.n27 0.037
R2012 GND.n364 GND.n362 0.035
R2013 GND.n301 GND.n299 0.035
R2014 GND.n19 GND.n17 0.035
R2015 GND.n321 GND.n319 0.035
R2016 GND.n341 GND.n339 0.035
R2017 GND.n271 GND.n269 0.033
R2018 GND.n71 GND.n69 0.033
R2019 GND.n40 GND.n38 0.032
R2020 GND.n191 GND.n179 0.031
R2021 GND.n169 GND.n167 0.031
R2022 GND.n258 GND.n256 0.029
R2023 GND.n85 GND.n83 0.029
R2024 GND.n205 GND.n195 0.027
R2025 GND.n153 GND.n151 0.027
R2026 GND GND.n366 0.027
R2027 GND.n246 GND.n244 0.025
R2028 GND.n99 GND.n97 0.025
R2029 GND.n217 GND.n209 0.022
R2030 GND.n139 GND.n137 0.022
R2031 GND.n233 GND.n231 0.02
R2032 GND.n113 GND.n111 0.02
R2033 GND.n229 GND.n221 0.018
R2034 GND.n125 GND.n123 0.018
R2035 GND.n221 GND.n219 0.016
R2036 GND.n127 GND.n125 0.016
R2037 GND.n242 GND.n233 0.014
R2038 GND.n111 GND.n109 0.014
R2039 GND.n209 GND.n207 0.012
R2040 GND.n141 GND.n139 0.012
R2041 GND.n362 GND.n360 0.01
R2042 GND.n254 GND.n246 0.01
R2043 GND.n97 GND.n95 0.01
R2044 GND.n38 GND.n36 0.01
R2045 GND.n299 GND.n297 0.01
R2046 GND.n17 GND.n15 0.01
R2047 GND.n319 GND.n317 0.01
R2048 GND.n339 GND.n337 0.01
R2049 GND.n195 GND.n193 0.008
R2050 GND.n155 GND.n153 0.008
R2051 GND.n344 GND.n343 0.007
R2052 GND.n267 GND.n258 0.006
R2053 GND.n83 GND.n81 0.006
R2054 GND.n351 GND.n349 0.005
R2055 GND.n27 GND.n25 0.005
R2056 GND.n288 GND.n286 0.005
R2057 GND.n6 GND.n4 0.005
R2058 GND.n308 GND.n306 0.005
R2059 GND.n328 GND.n326 0.005
R2060 GND.n179 GND.n177 0.004
R2061 GND.n171 GND.n169 0.004
R2062 GND.n279 GND.n271 0.002
R2063 GND.n69 GND.n67 0.002
R2064 modi.n0 modi.t0 1037.95
R2065 modi.n0 modi.t1 796.858
R2066 modi modi.n0 3.352
R2067 31.n0 31.t4 730.676
R2068 31.n0 31.t3 395.824
R2069 31.n323 31.n28 92.5
R2070 31.n323 31.n16 92.219
R2071 31.n323 31.n20 92.219
R2072 31.n323 31.n14 91.846
R2073 31.n323 31.n23 91.846
R2074 31.n323 31.n24 91.661
R2075 31.n323 31.n12 91.661
R2076 31.n34 31.n11 19.393
R2077 31.n26 31.n10 19.393
R2078 31.n92 31.n17 19.059
R2079 31.n131 31.n18 19.059
R2080 31.n182 31.n25 18.597
R2081 31.n148 31.n21 18.438
R2082 31.n48 31.n31 18.22
R2083 31.n277 31.n15 18.061
R2084 31.n176 31.n24 15.231
R2085 31.n300 31.n12 14.855
R2086 31.n138 31.n20 14.115
R2087 31.n265 31.n16 13.739
R2088 31.n164 31.n23 13.356
R2089 31.n106 31.n28 13.176
R2090 31.n115 31.n28 13.176
R2091 31.n287 31.n14 12.979
R2092 31.n1 31.t0 11.728
R2093 31.n1 31.t2 10.985
R2094 31.n35 31.n34 9.3
R2095 31.n327 31.n10 9.3
R2096 31.n47 31.n42 9.3
R2097 31.n49 31.n48 9.3
R2098 31.n153 31.n147 9.3
R2099 31.n155 31.n154 9.3
R2100 31.n131 31.n130 9.3
R2101 31.n261 31.n259 9.3
R2102 31.n263 31.n262 9.3
R2103 31.n275 31.n274 9.3
R2104 31.n291 31.n13 9.3
R2105 31.n323 31.n13 9.3
R2106 31.n290 31.n289 9.3
R2107 31.n300 31.n299 9.3
R2108 31.n52 31.n50 9.3
R2109 31.n302 31.n301 9.3
R2110 31.n288 31.n65 9.3
R2111 31.n276 31.n75 9.3
R2112 31.n273 31.n30 9.3
R2113 31.n323 31.n30 9.3
R2114 31.n264 31.n82 9.3
R2115 31.n120 31.n119 9.3
R2116 31.n116 31.n115 9.3
R2117 31.n107 31.n106 9.3
R2118 31.n104 31.n103 9.3
R2119 31.n93 31.n92 9.3
R2120 31.n88 31.n29 9.3
R2121 31.n323 31.n29 9.3
R2122 31.n84 31.n83 9.3
R2123 31.n137 31.n136 9.3
R2124 31.n135 31.n19 9.3
R2125 31.n323 31.n19 9.3
R2126 31.n156 31.n22 9.3
R2127 31.n323 31.n22 9.3
R2128 31.n210 31.n209 9.3
R2129 31.n206 31.n27 9.3
R2130 31.n323 31.n27 9.3
R2131 31.n208 31.n207 9.3
R2132 31.n187 31.n186 9.3
R2133 31.n183 31.n181 9.3
R2134 31.n182 31.n179 9.3
R2135 31.n44 31.n43 9.3
R2136 31.n324 31.n4 9.3
R2137 31.n322 31.n321 9.3
R2138 31.n324 31.n323 8.47
R2139 31.n323 31.n322 8.469
R2140 31.n323 31.n26 8.124
R2141 31.n323 31.n11 8.124
R2142 31.n323 31.n31 8.097
R2143 31.n323 31.n25 8.097
R2144 31.n323 31.n21 8.016
R2145 31.n323 31.n15 8.016
R2146 31.n323 31.n18 7.964
R2147 31.n323 31.n17 7.964
R2148 31.n139 31.n138 6.4
R2149 31.n177 31.n176 6.4
R2150 31.n301 31.n53 6.023
R2151 31.n264 31.n263 6.023
R2152 31.n91 31.n29 6.023
R2153 31.n105 31.n104 6.023
R2154 31.n119 31.n118 6.023
R2155 31.n34 31.n32 5.647
R2156 31.n132 31.n19 5.647
R2157 31.n184 31.n183 5.647
R2158 31.n325 31.n10 5.647
R2159 31.n83 31.n16 5.457
R2160 31.n47 31.n46 5.27
R2161 31.n136 31.n20 5.08
R2162 31.n176 31.n175 4.65
R2163 31.n140 31.n139 4.65
R2164 31.n335 31.n334 4.524
R2165 31.n289 31.n13 4.517
R2166 31.n208 31.n27 4.517
R2167 31.n317 31.n316 4.5
R2168 31.n329 31.n328 4.5
R2169 31.n315 31.n314 4.5
R2170 31.n309 31.n308 4.5
R2171 31.n56 31.n54 4.5
R2172 31.n71 31.n69 4.5
R2173 31.n260 31.n80 4.5
R2174 31.n89 31.n85 4.5
R2175 31.n102 31.n101 4.5
R2176 31.n114 31.n113 4.5
R2177 31.n134 31.n128 4.5
R2178 31.n145 31.n141 4.5
R2179 31.n162 31.n161 4.5
R2180 31.n192 31.n191 4.5
R2181 31.n188 31.n184 4.5
R2182 31.n193 31.n174 4.5
R2183 31.n205 31.n165 4.5
R2184 31.n211 31.n164 4.5
R2185 31.n163 31.n151 4.5
R2186 31.n146 31.n143 4.5
R2187 31.n219 31.n148 4.5
R2188 31.n133 31.n132 4.5
R2189 31.n118 31.n117 4.5
R2190 31.n105 31.n99 4.5
R2191 31.n91 31.n90 4.5
R2192 31.n257 31.n256 4.5
R2193 31.n77 31.n76 4.5
R2194 31.n278 31.n277 4.5
R2195 31.n70 31.n67 4.5
R2196 31.n61 31.n60 4.5
R2197 31.n303 31.n53 4.5
R2198 31.n307 31.n41 4.5
R2199 31.n292 31.n64 4.5
R2200 31.n287 31.n286 4.5
R2201 31.n73 31.n72 4.5
R2202 31.n266 31.n265 4.5
R2203 31.n251 31.n95 4.5
R2204 31.n245 31.n244 4.5
R2205 31.n243 31.n242 4.5
R2206 31.n237 31.n236 4.5
R2207 31.n235 31.n234 4.5
R2208 31.n229 31.n228 4.5
R2209 31.n159 31.n158 4.5
R2210 31.n9 31.n7 4.5
R2211 31.n46 31.n45 4.5
R2212 31.n326 31.n325 4.5
R2213 31.n327 31.n8 4.5
R2214 31.n318 31.n35 4.5
R2215 31.n320 31.n32 4.5
R2216 31.n64 31.n12 4.314
R2217 31.n276 31.n275 4.141
R2218 31.n154 31.n153 4.141
R2219 31.n72 31.n14 3.944
R2220 31.n165 31.n24 3.937
R2221 31.n158 31.n23 3.567
R2222 31.n336 31.n335 3.438
R2223 31.n57 31.n51 3.41
R2224 31.n78 31.n74 3.41
R2225 31.n39 31.n36 3.41
R2226 31.n311 31.n310 3.41
R2227 31.n58 31.n55 3.41
R2228 31.n280 31.n68 3.41
R2229 31.n269 31.n268 3.41
R2230 31.n298 31.n297 3.41
R2231 31.n306 31.n305 3.41
R2232 31.n294 31.n62 3.41
R2233 31.n284 31.n66 3.41
R2234 31.n272 31.n271 3.41
R2235 31.n313 31.n37 3.41
R2236 31.n251 31.n86 3.41
R2237 31.n126 31.n124 3.41
R2238 31.n144 31.n142 3.41
R2239 31.n255 31.n254 3.41
R2240 31.n250 31.n249 3.41
R2241 31.n122 31.n112 3.41
R2242 31.n231 31.n230 3.41
R2243 31.n224 31.n223 3.41
R2244 31.n217 31.n216 3.41
R2245 31.n258 31.n81 3.41
R2246 31.n252 31.n94 3.41
R2247 31.n246 31.n108 3.41
R2248 31.n241 31.n110 3.41
R2249 31.n238 31.n121 3.41
R2250 31.n233 31.n123 3.41
R2251 31.n227 31.n129 3.41
R2252 31.n157 31.n149 3.41
R2253 31.n203 31.n166 3.41
R2254 31.n213 31.n212 3.41
R2255 31.n221 31.n220 3.41
R2256 31.n198 31.n197 3.41
R2257 31.n334 31.n333 3.41
R2258 31.n199 31.n169 3.41
R2259 31.n190 31.n173 3.41
R2260 31.n331 31.n330 3.41
R2261 31.n200 31.n171 3.41
R2262 31.n195 31.n194 3.41
R2263 31.n185 31.n180 3.41
R2264 31.n3 31.n2 3.41
R2265 31.n226 31.n138 3.033
R2266 31.n178 31.n177 3.033
R2267 31.n323 31.t1 2.9
R2268 31.n275 31.n30 2.258
R2269 31.n154 31.n22 2.258
R2270 31.n170 31.n168 2.25
R2271 31.n321 31.n33 1.962
R2272 31.n100 31.n96 1.94
R2273 31.n289 31.n288 1.882
R2274 31.n288 31.n287 1.882
R2275 31.n209 31.n208 1.882
R2276 31.n63 31.n59 1.705
R2277 31.n109 31.n97 1.705
R2278 31.n167 31.n150 1.705
R2279 31.n158 31.n22 1.505
R2280 31.n209 31.n164 1.505
R2281 31.n189 31.n188 1.5
R2282 31.n205 31.n204 1.5
R2283 31.n117 31.n111 1.5
R2284 31.n99 31.n98 1.5
R2285 31.n90 31.n87 1.5
R2286 31.n304 31.n303 1.5
R2287 31.n293 31.n292 1.5
R2288 31.n286 31.n285 1.5
R2289 31.n279 31.n278 1.5
R2290 31.n267 31.n266 1.5
R2291 31.n133 31.n125 1.5
R2292 31.n226 31.n225 1.5
R2293 31.n211 31.n152 1.5
R2294 31.n219 31.n218 1.5
R2295 31.n160 31.n159 1.5
R2296 31.n178 31.n172 1.5
R2297 31.n45 31.n38 1.5
R2298 31.n326 31.n5 1.5
R2299 31.n320 31.n319 1.5
R2300 31.n337 31.n1 1.345
R2301 31.n297 31.n296 1.137
R2302 31.n305 31.n40 1.137
R2303 31.n295 31.n294 1.137
R2304 31.n284 31.n283 1.137
R2305 31.n282 31.n281 1.137
R2306 31.n271 31.n270 1.137
R2307 31.n253 31.n252 1.137
R2308 31.n248 31.n96 1.137
R2309 31.n247 31.n246 1.137
R2310 31.n241 31.n240 1.137
R2311 31.n239 31.n238 1.137
R2312 31.n233 31.n232 1.137
R2313 31.n215 31.n149 1.137
R2314 31.n203 31.n202 1.137
R2315 31.n214 31.n213 1.137
R2316 31.n222 31.n221 1.137
R2317 31.n333 31.n332 1.137
R2318 31.n201 31.n200 1.137
R2319 31.n196 31.n195 1.137
R2320 31.n46 31.n43 1.129
R2321 31.n48 31.n47 1.129
R2322 31.n72 31.n30 1.129
R2323 31.n277 31.n276 1.129
R2324 31.n281 31.n73 1.042
R2325 31.n337 31.n336 0.983
R2326 31.n313 31.n312 0.853
R2327 31.n81 31.n79 0.853
R2328 31.n129 31.n127 0.853
R2329 31.n180 31.n6 0.853
R2330 31.n322 31.n32 0.752
R2331 31.n132 31.n131 0.752
R2332 31.n136 31.n19 0.752
R2333 31.n153 31.n148 0.752
R2334 31.n165 31.n27 0.752
R2335 31.n183 31.n182 0.752
R2336 31.n186 31.n184 0.752
R2337 31.n325 31.n324 0.752
R2338 31.n39 31.n33 0.717
R2339 31 31.n337 0.566
R2340 31.n119 31.n18 0.536
R2341 31.n104 31.n17 0.536
R2342 31.n259 31.n15 0.475
R2343 31.n139 31.n21 0.475
R2344 31.n177 31.n25 0.382
R2345 31.n52 31.n31 0.382
R2346 31.n53 31.n52 0.376
R2347 31.n301 31.n300 0.376
R2348 31.n64 31.n13 0.376
R2349 31.n263 31.n259 0.376
R2350 31.n265 31.n264 0.376
R2351 31.n83 31.n29 0.376
R2352 31.n92 31.n91 0.376
R2353 31.n106 31.n105 0.376
R2354 31.n118 31.n115 0.376
R2355 31.n43 31.n11 0.349
R2356 31.n186 31.n26 0.349
R2357 31 31.n338 0.137
R2358 31.n338 31.n0 0.063
R2359 31.n316 31.n315 0.047
R2360 31.n257 31.n84 0.047
R2361 31.n100 31.n95 0.047
R2362 31.n244 31.n243 0.047
R2363 31.n236 31.n235 0.047
R2364 31.n228 31.n137 0.047
R2365 31.n328 31.n9 0.047
R2366 31.n170 31.n166 0.043
R2367 31.n203 31.n168 0.043
R2368 31.n62 31.n61 0.041
R2369 31.n294 31.n60 0.041
R2370 31.n194 31.n193 0.035
R2371 31.n246 31.n98 0.035
R2372 31.n241 31.n111 0.035
R2373 31.n195 31.n174 0.035
R2374 31.n307 31.n306 0.034
R2375 31.n108 31.n107 0.034
R2376 31.n116 31.n110 0.034
R2377 31.n192 31.n179 0.034
R2378 31.n310 31.n309 0.034
R2379 31.n305 31.n41 0.034
R2380 31.n268 31.n80 0.034
R2381 31.n255 31.n85 0.034
R2382 31.n233 31.n125 0.034
R2383 31.n230 31.n128 0.034
R2384 31.n224 31.n141 0.034
R2385 31.n191 31.n190 0.034
R2386 31.n308 31.n49 0.032
R2387 31.n226 31.n140 0.032
R2388 31.n178 31.n175 0.032
R2389 31.n252 31.n87 0.032
R2390 31.n190 31.n189 0.032
R2391 31.n311 31.n40 0.031
R2392 31.n270 31.n269 0.031
R2393 31.n196 31.n173 0.031
R2394 31.n332 31.n331 0.031
R2395 31.n303 31.n302 0.03
R2396 31.n262 31.n82 0.03
R2397 31.n94 31.n93 0.03
R2398 31.n130 31.n123 0.03
R2399 31.n185 31.n9 0.03
R2400 31.n310 31.n38 0.03
R2401 31.n55 31.n51 0.03
R2402 31.n251 31.n250 0.03
R2403 31.n124 31.n122 0.03
R2404 31.n230 31.n229 0.03
R2405 31.n199 31.n198 0.03
R2406 31.n180 31.n7 0.03
R2407 31.n254 31.n253 0.03
R2408 31.n232 31.n231 0.03
R2409 31.n223 31.n222 0.03
R2410 31.n320 31.n35 0.028
R2411 31.n315 31.n37 0.028
R2412 31.n298 31.n54 0.028
R2413 31.n70 31.n66 0.028
R2414 31.n73 31.n71 0.028
R2415 31.n272 31.n76 0.028
R2416 31.n227 31.n226 0.028
R2417 31.n212 31.n163 0.028
R2418 31.n171 31.n170 0.028
R2419 31.n188 31.n181 0.028
R2420 31.n327 31.n326 0.028
R2421 31.n319 31.n318 0.028
R2422 31.n314 31.n313 0.028
R2423 31.n297 31.n56 0.028
R2424 31.n284 31.n67 0.028
R2425 31.n281 31.n69 0.028
R2426 31.n271 31.n77 0.028
R2427 31.n256 31.n255 0.028
R2428 31.n101 31.n96 0.028
R2429 31.n238 31.n113 0.028
R2430 31.n225 31.n129 0.028
R2431 31.n213 31.n151 0.028
R2432 31.n200 31.n168 0.028
R2433 31.n8 31.n5 0.028
R2434 31.n296 31.n295 0.027
R2435 31.n283 31.n282 0.027
R2436 31.n45 31.n42 0.026
R2437 31.n266 31.n258 0.026
R2438 31.n220 31.n146 0.026
R2439 31.n162 31.n159 0.026
R2440 31.n280 31.n279 0.026
R2441 31.n267 31.n81 0.026
R2442 31.n221 31.n143 0.026
R2443 31.n161 31.n160 0.026
R2444 31.n204 31.n167 0.026
R2445 31.n330 31.n329 0.026
R2446 31.n248 31.n247 0.026
R2447 31.n240 31.n239 0.026
R2448 31.n215 31.n214 0.026
R2449 31.n202 31.n201 0.026
R2450 31.n319 31.n33 0.024
R2451 31.n261 31.n260 0.024
R2452 31.n145 31.n140 0.024
R2453 31.n317 31.n36 0.024
R2454 31.n293 31.n63 0.024
R2455 31.n268 31.n267 0.024
R2456 31.n242 31.n109 0.024
R2457 31.n218 31.n217 0.024
R2458 31.n291 31.n290 0.022
R2459 31.n258 31.n257 0.022
R2460 31.n103 31.n102 0.022
R2461 31.n120 31.n114 0.022
R2462 31.n146 31.n145 0.022
R2463 31.n220 31.n219 0.022
R2464 31.n207 31.n206 0.022
R2465 31.n314 31.n36 0.022
R2466 31.n256 31.n81 0.022
R2467 31.n245 31.n109 0.022
R2468 31.n225 31.n224 0.022
R2469 31.n143 31.n141 0.022
R2470 31.n274 31.n75 0.02
R2471 31.n278 31.n272 0.02
R2472 31.n260 31.n76 0.02
R2473 31.n228 31.n227 0.02
R2474 31.n155 31.n147 0.02
R2475 31.n313 31.n38 0.02
R2476 31.n80 31.n77 0.02
R2477 31.n229 31.n129 0.02
R2478 31.n330 31.n7 0.02
R2479 31.n333 31.n5 0.02
R2480 31.n312 31.n39 0.019
R2481 31.n312 31.n311 0.019
R2482 31.n173 31.n6 0.019
R2483 31.n331 31.n6 0.019
R2484 31.n175 31.n171 0.018
R2485 31.n285 31.n63 0.018
R2486 31.n189 31.n180 0.018
R2487 31.n269 31.n79 0.018
R2488 31.n254 31.n79 0.018
R2489 31.n231 31.n127 0.018
R2490 31.n223 31.n127 0.018
R2491 31.n299 31.n298 0.017
R2492 31.n90 31.n89 0.017
R2493 31.n95 31.n94 0.017
R2494 31.n334 31.n4 0.017
R2495 31.n297 31.n55 0.017
R2496 31.n281 31.n280 0.017
R2497 31.n271 31.n74 0.017
R2498 31.n87 31.n85 0.017
R2499 31.n252 31.n251 0.017
R2500 31.n250 31.n96 0.017
R2501 31.n221 31.n144 0.017
R2502 31.n217 31.n149 0.017
R2503 31.n167 31.n152 0.017
R2504 31.n200 31.n199 0.017
R2505 31.n333 31.n3 0.017
R2506 31.n44 31.n37 0.015
R2507 31.n308 31.n307 0.015
R2508 31.n71 31.n70 0.015
R2509 31.n235 31.n123 0.015
R2510 31.n134 31.n133 0.015
R2511 31.n163 31.n162 0.015
R2512 31.n212 31.n211 0.015
R2513 31.n187 31.n185 0.015
R2514 31.n309 31.n41 0.015
R2515 31.n305 31.n304 0.015
R2516 31.n69 31.n67 0.015
R2517 31.n237 31.n122 0.015
R2518 31.n234 31.n233 0.015
R2519 31.n128 31.n125 0.015
R2520 31.n161 31.n151 0.015
R2521 31.n213 31.n152 0.015
R2522 31.n306 31.n50 0.013
R2523 31.n286 31.n66 0.013
R2524 31.n89 31.n88 0.013
R2525 31.n135 31.n134 0.013
R2526 31.n194 31.n178 0.013
R2527 31.n193 31.n192 0.013
R2528 31.n285 31.n284 0.013
R2529 31.n195 31.n172 0.013
R2530 31.n191 31.n174 0.013
R2531 31.n336 31.n2 0.013
R2532 31.n295 31.n59 0.012
R2533 31.n283 31.n59 0.012
R2534 31.n274 31.n273 0.011
R2535 31.n156 31.n155 0.011
R2536 31.n58 31.n57 0.011
R2537 31.n78 31.n68 0.011
R2538 31.n249 31.n86 0.011
R2539 31.n247 31.n97 0.011
R2540 31.n240 31.n97 0.011
R2541 31.n126 31.n112 0.011
R2542 31.n216 31.n142 0.011
R2543 31.n214 31.n150 0.011
R2544 31.n202 31.n150 0.011
R2545 31.n197 31.n169 0.011
R2546 31.n316 31.n35 0.009
R2547 31.n290 31.n65 0.009
R2548 31.n286 31.n65 0.009
R2549 31.n244 31.n108 0.009
R2550 31.n210 31.n207 0.009
R2551 31.n318 31.n317 0.009
R2552 31.n246 31.n245 0.009
R2553 31.n292 31.n62 0.007
R2554 31.n102 31.n99 0.007
R2555 31.n243 31.n110 0.007
R2556 31.n117 31.n114 0.007
R2557 31.n211 31.n210 0.007
R2558 31.n328 31.n327 0.007
R2559 31.n294 31.n293 0.007
R2560 31.n101 31.n98 0.007
R2561 31.n242 31.n241 0.007
R2562 31.n113 31.n111 0.007
R2563 31.n329 31.n8 0.007
R2564 31.n335 31.n3 0.007
R2565 31.n338 31 0.007
R2566 31.n57 31.n40 0.006
R2567 31.n296 31.n58 0.006
R2568 31.n282 31.n68 0.006
R2569 31.n270 31.n78 0.006
R2570 31.n253 31.n86 0.006
R2571 31.n249 31.n248 0.006
R2572 31.n239 31.n112 0.006
R2573 31.n232 31.n126 0.006
R2574 31.n222 31.n142 0.006
R2575 31.n216 31.n215 0.006
R2576 31.n201 31.n169 0.006
R2577 31.n197 31.n196 0.006
R2578 31.n332 31.n2 0.006
R2579 31.n45 31.n44 0.005
R2580 31.n49 31.n42 0.005
R2581 31.n273 31.n73 0.005
R2582 31.n278 31.n75 0.005
R2583 31.n103 31.n100 0.005
R2584 31.n121 31.n120 0.005
R2585 31.n157 31.n156 0.005
R2586 31.n205 31.n166 0.005
R2587 31.n218 31.n144 0.005
R2588 31.n204 31.n203 0.005
R2589 31.n321 31.n320 0.003
R2590 31.n133 31.n130 0.003
R2591 31.n137 31.n135 0.003
R2592 31.n219 31.n147 0.003
R2593 31.n206 31.n205 0.003
R2594 31.n181 31.n179 0.003
R2595 31.n188 31.n187 0.003
R2596 31.n326 31.n4 0.003
R2597 31.n279 31.n74 0.003
R2598 31.n198 31.n172 0.003
R2599 31.n303 31.n50 0.001
R2600 31.n302 31.n299 0.001
R2601 31.n61 31.n54 0.001
R2602 31.n292 31.n291 0.001
R2603 31.n262 31.n261 0.001
R2604 31.n266 31.n82 0.001
R2605 31.n88 31.n84 0.001
R2606 31.n93 31.n90 0.001
R2607 31.n107 31.n99 0.001
R2608 31.n117 31.n116 0.001
R2609 31.n236 31.n121 0.001
R2610 31.n159 31.n157 0.001
R2611 31.n304 31.n51 0.001
R2612 31.n60 31.n56 0.001
R2613 31.n238 31.n237 0.001
R2614 31.n234 31.n124 0.001
R2615 31.n160 31.n149 0.001
R2616 net2.n1 net2.n0 13.361
R2617 net2.n86 net2.n85 13.361
R2618 net2.n11 net2.n9 9.3
R2619 net2.n5 net2.n3 9.3
R2620 net2.n16 net2.n13 9.3
R2621 net2.n141 net2.n133 9.3
R2622 net2.n141 net2.n140 9.3
R2623 net2.n22 net2.n20 9.3
R2624 net2.n33 net2.n31 9.3
R2625 net2.n30 net2.n28 9.3
R2626 net2.n41 net2.n39 9.3
R2627 net2.n41 net2.n40 9.3
R2628 net2.n52 net2.n50 9.3
R2629 net2.n52 net2.n51 9.3
R2630 net2.n63 net2.n61 9.3
R2631 net2.n63 net2.n62 9.3
R2632 net2.n74 net2.n72 9.3
R2633 net2.n74 net2.n73 9.3
R2634 net2.n98 net2.n96 9.3
R2635 net2.n98 net2.n97 9.3
R2636 net2.n109 net2.n107 9.3
R2637 net2.n109 net2.n108 9.3
R2638 net2.n167 net2.n118 9.3
R2639 net2.n167 net2.n166 9.3
R2640 net2.n160 net2.n122 9.3
R2641 net2.n160 net2.n159 9.3
R2642 net2.n153 net2.n126 9.3
R2643 net2.n153 net2.n152 9.3
R2644 net2.n27 net2.n24 9.3
R2645 net2.n33 net2.n32 9.3
R2646 net2.n38 net2.n35 9.3
R2647 net2.n44 net2.n42 9.3
R2648 net2.n49 net2.n46 9.3
R2649 net2.n55 net2.n53 9.3
R2650 net2.n60 net2.n57 9.3
R2651 net2.n66 net2.n64 9.3
R2652 net2.n71 net2.n68 9.3
R2653 net2.n77 net2.n75 9.3
R2654 net2.n82 net2.n79 9.3
R2655 net2.n92 net2.n89 9.3
R2656 net2.n95 net2.n93 9.3
R2657 net2.n103 net2.n100 9.3
R2658 net2.n106 net2.n104 9.3
R2659 net2.n116 net2.n112 9.3
R2660 net2.n169 net2.n117 9.3
R2661 net2.n165 net2.n120 9.3
R2662 net2.n162 net2.n121 9.3
R2663 net2.n158 net2.n124 9.3
R2664 net2.n155 net2.n125 9.3
R2665 net2.n151 net2.n128 9.3
R2666 net2.n148 net2.n129 9.3
R2667 net2.n144 net2.n132 9.3
R2668 net2.n146 net2.n130 9.3
R2669 net2.n38 net2.n37 9.3
R2670 net2.n44 net2.n43 9.3
R2671 net2.n49 net2.n48 9.3
R2672 net2.n55 net2.n54 9.3
R2673 net2.n60 net2.n59 9.3
R2674 net2.n66 net2.n65 9.3
R2675 net2.n71 net2.n70 9.3
R2676 net2.n77 net2.n76 9.3
R2677 net2.n82 net2.n81 9.3
R2678 net2.n92 net2.n91 9.3
R2679 net2.n95 net2.n94 9.3
R2680 net2.n103 net2.n102 9.3
R2681 net2.n106 net2.n105 9.3
R2682 net2.n116 net2.n115 9.3
R2683 net2.n169 net2.n168 9.3
R2684 net2.n165 net2.n164 9.3
R2685 net2.n162 net2.n161 9.3
R2686 net2.n158 net2.n157 9.3
R2687 net2.n155 net2.n154 9.3
R2688 net2.n151 net2.n150 9.3
R2689 net2.n148 net2.n147 9.3
R2690 net2.n144 net2.n143 9.3
R2691 net2.n146 net2.n145 9.3
R2692 net2.n30 net2.n29 9.3
R2693 net2.n27 net2.n26 9.3
R2694 net2.n22 net2.n21 9.3
R2695 net2.n19 net2.n17 9.3
R2696 net2.n19 net2.n18 9.3
R2697 net2.n16 net2.n15 9.3
R2698 net2.n137 net2.n135 9.3
R2699 net2.n139 net2.n134 9.3
R2700 net2.n139 net2.n138 9.3
R2701 net2.n137 net2.n136 9.3
R2702 net2.n11 net2.n10 9.3
R2703 net2.n8 net2.n6 9.3
R2704 net2.n8 net2.n7 9.3
R2705 net2.n5 net2.n4 9.3
R2706 net2.n114 net2.n113 8.016
R2707 net2.n111 net2.n110 8.016
R2708 net2.n84 net2.n2 4.558
R2709 net2.n87 net2.n1 4.558
R2710 net2.n84 net2.n83 4.558
R2711 net2.n87 net2.n86 4.558
R2712 net2.n113 net2.t0 2.9
R2713 net2.n110 net2.t1 2.9
R2714 net2.n79 net2.n78 0.536
R2715 net2.n89 net2.n88 0.536
R2716 net2.n81 net2.n80 0.536
R2717 net2.n91 net2.n90 0.536
R2718 net2.n70 net2.n69 0.506
R2719 net2.n102 net2.n101 0.506
R2720 net2.n68 net2.n67 0.506
R2721 net2.n100 net2.n99 0.506
R2722 net2.n57 net2.n56 0.475
R2723 net2.n112 net2.n111 0.475
R2724 net2.n59 net2.n58 0.475
R2725 net2.n115 net2.n114 0.475
R2726 net2.n164 net2.n163 0.445
R2727 net2.n46 net2.n45 0.445
R2728 net2.n120 net2.n119 0.445
R2729 net2.n48 net2.n47 0.445
R2730 net2.n35 net2.n34 0.413
R2731 net2.n124 net2.n123 0.413
R2732 net2.n37 net2.n36 0.413
R2733 net2.n157 net2.n156 0.413
R2734 net2.n26 net2.n25 0.382
R2735 net2.n150 net2.n149 0.382
R2736 net2.n128 net2.n127 0.382
R2737 net2.n24 net2.n23 0.382
R2738 net2.n13 net2.n12 0.349
R2739 net2.n15 net2.n14 0.349
R2740 net2.n132 net2.n131 0.349
R2741 net2.n143 net2.n142 0.349
R2742 net2.n87 net2.n84 0.039
R2743 net2.n16 net2.n11 0.03
R2744 net2.n27 net2.n22 0.03
R2745 net2.n38 net2.n33 0.03
R2746 net2.n49 net2.n44 0.03
R2747 net2.n60 net2.n55 0.03
R2748 net2.n71 net2.n66 0.03
R2749 net2.n82 net2.n77 0.03
R2750 net2.n95 net2.n92 0.03
R2751 net2.n106 net2.n103 0.03
R2752 net2.n165 net2.n162 0.03
R2753 net2.n158 net2.n155 0.03
R2754 net2.n151 net2.n148 0.03
R2755 net2.n144 net2.n141 0.03
R2756 net2 net2.n169 0.018
R2757 net2 net2.n116 0.011
R2758 net2.n84 net2.n82 0.009
R2759 net2.n92 net2.n87 0.009
R2760 net2.n11 net2.n8 0.008
R2761 net2.n141 net2.n139 0.008
R2762 net2.n22 net2.n19 0.007
R2763 net2.n74 net2.n71 0.007
R2764 net2.n103 net2.n98 0.007
R2765 net2.n148 net2.n146 0.007
R2766 net2.n33 net2.n30 0.006
R2767 net2.n63 net2.n60 0.006
R2768 net2.n116 net2.n109 0.006
R2769 net2.n155 net2.n153 0.006
R2770 net2.n44 net2.n41 0.005
R2771 net2.n52 net2.n49 0.005
R2772 net2.n167 net2.n165 0.005
R2773 net2.n162 net2.n160 0.005
R2774 net2.n41 net2.n38 0.004
R2775 net2.n160 net2.n158 0.004
R2776 net2.n30 net2.n27 0.003
R2777 net2.n55 net2.n52 0.003
R2778 net2.n169 net2.n167 0.003
R2779 net2.n153 net2.n151 0.003
R2780 net2.n19 net2.n16 0.002
R2781 net2.n66 net2.n63 0.002
R2782 net2.n109 net2.n106 0.002
R2783 net2.n146 net2.n144 0.002
R2784 net2.n8 net2.n5 0.001
R2785 net2.n77 net2.n74 0.001
R2786 net2.n98 net2.n95 0.001
R2787 net2.n139 net2.n137 0.001
R2788 net3_ff1.n257 net3_ff1.t2 735.052
R2789 net3_ff1.n87 net3_ff1.t3 399.297
R2790 net3_ff1.n32 net3_ff1.n31 92.5
R2791 net3_ff1.n47 net3_ff1.n46 92.5
R2792 net3_ff1.n46 net3_ff1.t0 70.344
R2793 net3_ff1.n10 net3_ff1.n9 31.034
R2794 net3_ff1.n66 net3_ff1.n65 31.034
R2795 net3_ff1.n216 net3_ff1.n215 9.3
R2796 net3_ff1.n106 net3_ff1.n105 9.3
R2797 net3_ff1.n18 net3_ff1.n17 9.3
R2798 net3_ff1.n67 net3_ff1.n66 9.3
R2799 net3_ff1.n11 net3_ff1.n10 9.3
R2800 net3_ff1.n77 net3_ff1.n76 9.3
R2801 net3_ff1.n174 net3_ff1.n173 9.154
R2802 net3_ff1.n33 net3_ff1.n32 8.282
R2803 net3_ff1.n48 net3_ff1.n47 8.282
R2804 net3_ff1.n173 net3_ff1.t1 7.141
R2805 net3_ff1.n99 net3_ff1.n98 7.033
R2806 net3_ff1.n93 net3_ff1.n92 7.033
R2807 net3_ff1.n11 net3_ff1.n7 5.647
R2808 net3_ff1.n67 net3_ff1.n63 5.647
R2809 net3_ff1.n175 net3_ff1.n174 4.65
R2810 net3_ff1.n45 net3_ff1.n44 4.65
R2811 net3_ff1.n134 net3_ff1.n133 4.5
R2812 net3_ff1.n112 net3_ff1.n111 4.5
R2813 net3_ff1.n155 net3_ff1.n154 4.5
R2814 net3_ff1.n162 net3_ff1.n159 4.5
R2815 net3_ff1.n170 net3_ff1.n169 4.5
R2816 net3_ff1.n176 net3_ff1.n172 4.5
R2817 net3_ff1.n203 net3_ff1.n200 4.5
R2818 net3_ff1.n210 net3_ff1.n209 4.5
R2819 net3_ff1.n222 net3_ff1.n221 4.5
R2820 net3_ff1.n232 net3_ff1.n231 4.5
R2821 net3_ff1.n242 net3_ff1.n241 4.5
R2822 net3_ff1.n122 net3_ff1.n121 4.5
R2823 net3_ff1.n83 net3_ff1.n81 4.5
R2824 net3_ff1.n71 net3_ff1.n68 4.5
R2825 net3_ff1.n58 net3_ff1.n56 4.5
R2826 net3_ff1.n34 net3_ff1.n33 4.5
R2827 net3_ff1.n41 net3_ff1.n40 4.5
R2828 net3_ff1.n49 net3_ff1.n48 4.5
R2829 net3_ff1.n14 net3_ff1.n13 4.5
R2830 net3_ff1.n23 net3_ff1.n22 4.5
R2831 net3_ff1.n231 net3_ff1.n228 4.141
R2832 net3_ff1.n121 net3_ff1.n120 4.141
R2833 net3_ff1.n9 net3_ff1.n8 4.137
R2834 net3_ff1.n65 net3_ff1.n64 4.137
R2835 net3_ff1.n221 net3_ff1.n218 3.764
R2836 net3_ff1.n154 net3_ff1.n152 3.764
R2837 net3_ff1.n22 net3_ff1.n20 3.764
R2838 net3_ff1.n68 net3_ff1.n61 3.764
R2839 net3_ff1.n241 net3_ff1.n238 3.388
R2840 net3_ff1.n209 net3_ff1.n208 3.388
R2841 net3_ff1.n111 net3_ff1.n110 3.388
R2842 net3_ff1.n133 net3_ff1.n132 3.388
R2843 net3_ff1.n13 net3_ff1.n12 3.388
R2844 net3_ff1.n81 net3_ff1.n80 3.388
R2845 net3_ff1.n241 net3_ff1.n240 3.011
R2846 net3_ff1.n209 net3_ff1.n206 3.011
R2847 net3_ff1.n200 net3_ff1.n198 3.011
R2848 net3_ff1.n105 net3_ff1.n104 3.011
R2849 net3_ff1.n111 net3_ff1.n109 3.011
R2850 net3_ff1.n133 net3_ff1.n131 3.011
R2851 net3_ff1.n13 net3_ff1.n11 3.011
R2852 net3_ff1.n33 net3_ff1.n30 3.011
R2853 net3_ff1.n81 net3_ff1.n79 3.011
R2854 net3_ff1.n221 net3_ff1.n220 2.635
R2855 net3_ff1.n215 net3_ff1.n214 2.635
R2856 net3_ff1.n159 net3_ff1.n158 2.635
R2857 net3_ff1.n154 net3_ff1.n153 2.635
R2858 net3_ff1.n22 net3_ff1.n21 2.635
R2859 net3_ff1.n56 net3_ff1.n55 2.635
R2860 net3_ff1.n68 net3_ff1.n67 2.635
R2861 net3_ff1.n231 net3_ff1.n230 2.258
R2862 net3_ff1.n121 net3_ff1.n119 2.258
R2863 net3_ff1.n86 net3_ff1.n85 1.705
R2864 net3_ff1.n256 net3_ff1.n247 1.705
R2865 net3_ff1 net3_ff1.n87 1.685
R2866 net3_ff1.n159 net3_ff1.n157 1.505
R2867 net3_ff1.n156 net3_ff1.n155 1.5
R2868 net3_ff1.n163 net3_ff1.n162 1.5
R2869 net3_ff1.n171 net3_ff1.n170 1.5
R2870 net3_ff1.n177 net3_ff1.n176 1.5
R2871 net3_ff1.n84 net3_ff1.n83 1.5
R2872 net3_ff1.n72 net3_ff1.n71 1.5
R2873 net3_ff1.n35 net3_ff1.n34 1.5
R2874 net3_ff1.n59 net3_ff1.n58 1.5
R2875 net3_ff1.n42 net3_ff1.n41 1.5
R2876 net3_ff1.n50 net3_ff1.n49 1.5
R2877 net3_ff1.n27 net3_ff1.n14 1.5
R2878 net3_ff1.n24 net3_ff1.n23 1.5
R2879 net3_ff1.n200 net3_ff1.n199 1.129
R2880 net3_ff1.n100 net3_ff1.n99 1.127
R2881 net3_ff1.n247 net3_ff1.n93 1.127
R2882 net3_ff1.n243 net3_ff1.n242 1.125
R2883 net3_ff1.n135 net3_ff1.n134 1.125
R2884 net3_ff1.n7 net3_ff1.n6 0.752
R2885 net3_ff1.n63 net3_ff1.n62 0.752
R2886 net3_ff1.n92 net3_ff1.n91 0.155
R2887 net3_ff1.n98 net3_ff1.n97 0.155
R2888 net3_ff1.n240 net3_ff1.n239 0.144
R2889 net3_ff1.n131 net3_ff1.n130 0.144
R2890 net3_ff1.n230 net3_ff1.n229 0.133
R2891 net3_ff1.n119 net3_ff1.n118 0.132
R2892 net3_ff1.n87 net3_ff1.n86 0.117
R2893 net3_ff1.n257 net3_ff1.n256 0.112
R2894 net3_ff1 net3_ff1.n257 0.089
R2895 net3_ff1.n236 net3_ff1.n235 0.053
R2896 net3_ff1.n226 net3_ff1.n225 0.053
R2897 net3_ff1.n216 net3_ff1.n213 0.053
R2898 net3_ff1.n116 net3_ff1.n115 0.053
R2899 net3_ff1.n126 net3_ff1.n125 0.053
R2900 net3_ff1.n77 net3_ff1.n75 0.053
R2901 net3_ff1.n1 net3_ff1.n0 0.05
R2902 net3_ff1.n2 net3_ff1.n1 0.05
R2903 net3_ff1.n86 net3_ff1.n2 0.05
R2904 net3_ff1.n256 net3_ff1.n255 0.05
R2905 net3_ff1.n255 net3_ff1.n254 0.05
R2906 net3_ff1.n254 net3_ff1.n253 0.05
R2907 net3_ff1.n253 net3_ff1.n252 0.05
R2908 net3_ff1.n252 net3_ff1.n251 0.05
R2909 net3_ff1.n251 net3_ff1.n250 0.05
R2910 net3_ff1.n250 net3_ff1.n249 0.05
R2911 net3_ff1.n249 net3_ff1.n248 0.05
R2912 net3_ff1.n41 net3_ff1.n39 0.045
R2913 net3_ff1.n58 net3_ff1.n54 0.045
R2914 net3_ff1.n203 net3_ff1.n202 0.043
R2915 net3_ff1.n170 net3_ff1.n168 0.043
R2916 net3_ff1.n89 net3_ff1.n88 0.034
R2917 net3_ff1.n125 net3_ff1.n124 0.032
R2918 net3_ff1.n95 net3_ff1.n94 0.032
R2919 net3_ff1.n237 net3_ff1.n236 0.03
R2920 net3_ff1.n235 net3_ff1.n234 0.03
R2921 net3_ff1.n115 net3_ff1.n114 0.03
R2922 net3_ff1.n225 net3_ff1.n224 0.028
R2923 net3_ff1.n127 net3_ff1.n126 0.028
R2924 net3_ff1.n129 net3_ff1.n128 0.028
R2925 net3_ff1.n25 net3_ff1.n24 0.027
R2926 net3_ff1.n84 net3_ff1.n74 0.027
R2927 net3_ff1.n197 net3_ff1.n196 0.025
R2928 net3_ff1.n227 net3_ff1.n226 0.025
R2929 net3_ff1.n49 net3_ff1.n45 0.025
R2930 net3_ff1.n220 net3_ff1.n219 0.024
R2931 net3_ff1.n109 net3_ff1.n108 0.024
R2932 net3_ff1.n176 net3_ff1.n175 0.023
R2933 net3_ff1.n117 net3_ff1.n116 0.023
R2934 net3_ff1.n223 net3_ff1.n222 0.021
R2935 net3_ff1.n217 net3_ff1.n216 0.021
R2936 net3_ff1.n149 net3_ff1.n148 0.021
R2937 net3_ff1.n23 net3_ff1.n16 0.021
R2938 net3_ff1.n19 net3_ff1.n18 0.021
R2939 net3_ff1.n71 net3_ff1.n60 0.021
R2940 net3_ff1.n242 net3_ff1.n197 0.019
R2941 net3_ff1.n213 net3_ff1.n212 0.019
R2942 net3_ff1.n212 net3_ff1.n211 0.019
R2943 net3_ff1.n210 net3_ff1.n205 0.019
R2944 net3_ff1.n150 net3_ff1.n149 0.019
R2945 net3_ff1.n107 net3_ff1.n106 0.019
R2946 net3_ff1.n113 net3_ff1.n112 0.019
R2947 net3_ff1.n134 net3_ff1.n129 0.019
R2948 net3_ff1.n4 net3_ff1.n3 0.019
R2949 net3_ff1.n5 net3_ff1.n4 0.019
R2950 net3_ff1.n70 net3_ff1.n69 0.019
R2951 net3_ff1.n78 net3_ff1.n77 0.019
R2952 net3_ff1.n83 net3_ff1.n82 0.019
R2953 net3_ff1.n93 net3_ff1.n90 0.019
R2954 net3_ff1.n99 net3_ff1.n96 0.019
R2955 net3_ff1.n242 net3_ff1.n237 0.017
R2956 net3_ff1.n233 net3_ff1.n232 0.017
R2957 net3_ff1.n211 net3_ff1.n210 0.017
R2958 net3_ff1.n204 net3_ff1.n203 0.017
R2959 net3_ff1.n112 net3_ff1.n107 0.017
R2960 net3_ff1.n123 net3_ff1.n122 0.017
R2961 net3_ff1.n134 net3_ff1.n127 0.017
R2962 net3_ff1.n14 net3_ff1.n5 0.017
R2963 net3_ff1.n34 net3_ff1.n29 0.017
R2964 net3_ff1.n83 net3_ff1.n78 0.017
R2965 net3_ff1.n186 net3_ff1.n185 0.016
R2966 net3_ff1.n145 net3_ff1.n144 0.016
R2967 net3_ff1.n222 net3_ff1.n217 0.015
R2968 net3_ff1.n162 net3_ff1.n161 0.015
R2969 net3_ff1.n155 net3_ff1.n150 0.015
R2970 net3_ff1.n23 net3_ff1.n19 0.015
R2971 net3_ff1.n58 net3_ff1.n57 0.015
R2972 net3_ff1.n71 net3_ff1.n70 0.015
R2973 net3_ff1.n245 net3_ff1.n244 0.014
R2974 net3_ff1.n194 net3_ff1.n193 0.014
R2975 net3_ff1.n189 net3_ff1.n188 0.014
R2976 net3_ff1.n142 net3_ff1.n141 0.014
R2977 net3_ff1.n138 net3_ff1.n137 0.014
R2978 net3_ff1.n103 net3_ff1.n102 0.014
R2979 net3_ff1.n35 net3_ff1.n27 0.014
R2980 net3_ff1.n72 net3_ff1.n59 0.014
R2981 net3_ff1.n182 net3_ff1.n181 0.013
R2982 net3_ff1.n177 net3_ff1.n171 0.013
R2983 net3_ff1.n163 net3_ff1.n156 0.013
R2984 net3_ff1.n135 net3_ff1.n103 0.013
R2985 net3_ff1.n36 net3_ff1.n35 0.013
R2986 net3_ff1.n42 net3_ff1.n37 0.013
R2987 net3_ff1.n51 net3_ff1.n50 0.013
R2988 net3_ff1.n59 net3_ff1.n52 0.013
R2989 net3_ff1.n208 net3_ff1.n207 0.012
R2990 net3_ff1.n152 net3_ff1.n151 0.012
R2991 net3_ff1.n232 net3_ff1.n227 0.012
R2992 net3_ff1.n205 net3_ff1.n204 0.012
R2993 net3_ff1.n161 net3_ff1.n160 0.012
R2994 net3_ff1.n122 net3_ff1.n117 0.012
R2995 net3_ff1.n244 net3_ff1.n243 0.012
R2996 net3_ff1.n178 net3_ff1.n177 0.012
R2997 net3_ff1.n29 net3_ff1.n28 0.012
R2998 net3_ff1.n171 net3_ff1.n166 0.011
R2999 net3_ff1.n246 net3_ff1.n245 0.01
R3000 net3_ff1.n193 net3_ff1.n192 0.01
R3001 net3_ff1.n183 net3_ff1.n182 0.01
R3002 net3_ff1.n164 net3_ff1.n163 0.01
R3003 net3_ff1.n139 net3_ff1.n138 0.01
R3004 net3_ff1.n102 net3_ff1.n101 0.01
R3005 net3_ff1.n27 net3_ff1.n26 0.01
R3006 net3_ff1.n73 net3_ff1.n72 0.01
R3007 net3_ff1.n191 net3_ff1.n190 0.009
R3008 net3_ff1.n181 net3_ff1.n180 0.009
R3009 net3_ff1.n156 net3_ff1.n147 0.009
R3010 net3_ff1.n141 net3_ff1.n140 0.009
R3011 net3_ff1.n202 net3_ff1.n201 0.008
R3012 net3_ff1.n168 net3_ff1.n167 0.008
R3013 net3_ff1.n195 net3_ff1.n194 0.008
R3014 net3_ff1.n185 net3_ff1.n184 0.008
R3015 net3_ff1.n146 net3_ff1.n145 0.008
R3016 net3_ff1.n143 net3_ff1.n142 0.008
R3017 net3_ff1.n39 net3_ff1.n38 0.008
R3018 net3_ff1.n54 net3_ff1.n53 0.008
R3019 net3_ff1.n24 net3_ff1.n15 0.008
R3020 net3_ff1.n188 net3_ff1.n187 0.007
R3021 net3_ff1.n187 net3_ff1.n186 0.007
R3022 net3_ff1.n144 net3_ff1.n143 0.007
R3023 net3_ff1.n137 net3_ff1.n136 0.007
R3024 net3_ff1.n43 net3_ff1.n42 0.007
R3025 net3_ff1.n50 net3_ff1.n43 0.007
R3026 net3_ff1.n85 net3_ff1.n84 0.007
R3027 net3_ff1.n234 net3_ff1.n233 0.006
R3028 net3_ff1.n224 net3_ff1.n223 0.006
R3029 net3_ff1.n114 net3_ff1.n113 0.006
R3030 net3_ff1.n124 net3_ff1.n123 0.006
R3031 net3_ff1.n74 net3_ff1.n73 0.006
R3032 net3_ff1.n184 net3_ff1.n183 0.005
R3033 net3_ff1.n147 net3_ff1.n146 0.005
R3034 net3_ff1.n26 net3_ff1.n25 0.005
R3035 net3_ff1.n90 net3_ff1.n89 0.004
R3036 net3_ff1.n96 net3_ff1.n95 0.004
R3037 net3_ff1.n247 net3_ff1.n246 0.004
R3038 net3_ff1.n243 net3_ff1.n195 0.004
R3039 net3_ff1.n192 net3_ff1.n191 0.004
R3040 net3_ff1.n140 net3_ff1.n139 0.004
R3041 net3_ff1.n136 net3_ff1.n135 0.004
R3042 net3_ff1.n101 net3_ff1.n100 0.004
R3043 net3_ff1.n180 net3_ff1.n179 0.002
R3044 net3_ff1.n179 net3_ff1.n178 0.002
R3045 net3_ff1.n166 net3_ff1.n165 0.002
R3046 net3_ff1.n165 net3_ff1.n164 0.002
R3047 net3_ff1.n37 net3_ff1.n36 0.002
R3048 net3_ff1.n52 net3_ff1.n51 0.002
R3049 net3_ff1.n190 net3_ff1.n189 0.001
R3050 net4_ff1.n13 net4_ff1.n10 9.3
R3051 net4_ff1.n5 net4_ff1.n3 9.3
R3052 net4_ff1.n24 net4_ff1.n21 9.3
R3053 net4_ff1.n16 net4_ff1.n14 9.3
R3054 net4_ff1.n35 net4_ff1.n32 9.3
R3055 net4_ff1.n30 net4_ff1.n28 9.3
R3056 net4_ff1.n41 net4_ff1.n39 9.3
R3057 net4_ff1.n41 net4_ff1.n40 9.3
R3058 net4_ff1.n59 net4_ff1.n57 9.3
R3059 net4_ff1.n59 net4_ff1.n58 9.3
R3060 net4_ff1.n70 net4_ff1.n68 9.3
R3061 net4_ff1.n70 net4_ff1.n69 9.3
R3062 net4_ff1.n95 net4_ff1.n76 9.3
R3063 net4_ff1.n95 net4_ff1.n94 9.3
R3064 net4_ff1.n27 net4_ff1.n25 9.3
R3065 net4_ff1.n35 net4_ff1.n34 9.3
R3066 net4_ff1.n38 net4_ff1.n36 9.3
R3067 net4_ff1.n44 net4_ff1.n42 9.3
R3068 net4_ff1.n56 net4_ff1.n53 9.3
R3069 net4_ff1.n62 net4_ff1.n60 9.3
R3070 net4_ff1.n67 net4_ff1.n64 9.3
R3071 net4_ff1.n73 net4_ff1.n71 9.3
R3072 net4_ff1.n98 net4_ff1.n75 9.3
R3073 net4_ff1.n93 net4_ff1.n77 9.3
R3074 net4_ff1.n91 net4_ff1.n79 9.3
R3075 net4_ff1.n86 net4_ff1.n81 9.3
R3076 net4_ff1.n88 net4_ff1.n80 9.3
R3077 net4_ff1.n38 net4_ff1.n37 9.3
R3078 net4_ff1.n44 net4_ff1.n43 9.3
R3079 net4_ff1.n56 net4_ff1.n55 9.3
R3080 net4_ff1.n62 net4_ff1.n61 9.3
R3081 net4_ff1.n67 net4_ff1.n66 9.3
R3082 net4_ff1.n73 net4_ff1.n72 9.3
R3083 net4_ff1.n98 net4_ff1.n97 9.3
R3084 net4_ff1.n93 net4_ff1.n92 9.3
R3085 net4_ff1.n91 net4_ff1.n90 9.3
R3086 net4_ff1.n86 net4_ff1.n85 9.3
R3087 net4_ff1.n88 net4_ff1.n87 9.3
R3088 net4_ff1.n30 net4_ff1.n29 9.3
R3089 net4_ff1.n27 net4_ff1.n26 9.3
R3090 net4_ff1.n24 net4_ff1.n23 9.3
R3091 net4_ff1.n19 net4_ff1.n17 9.3
R3092 net4_ff1.n19 net4_ff1.n18 9.3
R3093 net4_ff1.n16 net4_ff1.n15 9.3
R3094 net4_ff1.n13 net4_ff1.n12 9.3
R3095 net4_ff1.n8 net4_ff1.n6 9.3
R3096 net4_ff1.n8 net4_ff1.n7 9.3
R3097 net4_ff1.n5 net4_ff1.n4 9.3
R3098 net4_ff1.n48 net4_ff1.t0 7.141
R3099 net4_ff1.n45 net4_ff1.t1 7.141
R3100 net4_ff1.n47 net4_ff1.n46 5.418
R3101 net4_ff1.n50 net4_ff1.n49 5.418
R3102 net4_ff1.n2 net4_ff1.n0 4.728
R3103 net4_ff1.n84 net4_ff1.n82 4.728
R3104 net4_ff1.n84 net4_ff1.n83 4.728
R3105 net4_ff1.n2 net4_ff1.n1 4.727
R3106 net4_ff1.n51 net4_ff1.n47 4.65
R3107 net4_ff1.n51 net4_ff1.n50 4.65
R3108 net4_ff1.n46 net4_ff1.n45 1.844
R3109 net4_ff1.n49 net4_ff1.n48 1.844
R3110 net4_ff1.n12 net4_ff1.n11 0.144
R3111 net4_ff1.n10 net4_ff1.n9 0.144
R3112 net4_ff1.n79 net4_ff1.n78 0.144
R3113 net4_ff1.n90 net4_ff1.n89 0.144
R3114 net4_ff1.n23 net4_ff1.n22 0.133
R3115 net4_ff1.n97 net4_ff1.n96 0.133
R3116 net4_ff1.n21 net4_ff1.n20 0.133
R3117 net4_ff1.n75 net4_ff1.n74 0.132
R3118 net4_ff1.n34 net4_ff1.n33 0.121
R3119 net4_ff1.n32 net4_ff1.n31 0.121
R3120 net4_ff1.n64 net4_ff1.n63 0.121
R3121 net4_ff1.n66 net4_ff1.n65 0.121
R3122 net4_ff1.n55 net4_ff1.n54 0.11
R3123 net4_ff1.n53 net4_ff1.n52 0.109
R3124 net4_ff1.n51 net4_ff1.n44 0.036
R3125 net4_ff1.n56 net4_ff1.n51 0.036
R3126 net4_ff1.n5 net4_ff1.n2 0.029
R3127 net4_ff1.n86 net4_ff1.n84 0.029
R3128 net4_ff1.n16 net4_ff1.n13 0.027
R3129 net4_ff1.n27 net4_ff1.n24 0.027
R3130 net4_ff1.n38 net4_ff1.n35 0.027
R3131 net4_ff1.n67 net4_ff1.n62 0.027
R3132 net4_ff1.n93 net4_ff1.n91 0.027
R3133 net4_ff1 net4_ff1.n73 0.016
R3134 net4_ff1 net4_ff1.n98 0.01
R3135 net4_ff1.n41 net4_ff1.n38 0.007
R3136 net4_ff1.n62 net4_ff1.n59 0.007
R3137 net4_ff1.n30 net4_ff1.n27 0.006
R3138 net4_ff1.n73 net4_ff1.n70 0.006
R3139 net4_ff1.n19 net4_ff1.n16 0.005
R3140 net4_ff1.n95 net4_ff1.n93 0.005
R3141 net4_ff1.n8 net4_ff1.n5 0.004
R3142 net4_ff1.n13 net4_ff1.n8 0.004
R3143 net4_ff1.n91 net4_ff1.n88 0.004
R3144 net4_ff1.n88 net4_ff1.n86 0.004
R3145 net4_ff1.n24 net4_ff1.n19 0.003
R3146 net4_ff1.n98 net4_ff1.n95 0.003
R3147 net4_ff1.n35 net4_ff1.n30 0.002
R3148 net4_ff1.n70 net4_ff1.n67 0.002
R3149 net4_ff1.n44 net4_ff1.n41 0.001
R3150 net4_ff1.n59 net4_ff1.n56 0.001
R3151 P.n0 P.t0 1037.77
R3152 P P.t1 796.138
R3153 P.n17 P.n16 2.25
R3154 P.n16 P.n15 1.742
R3155 P.n6 P.n5 1.705
R3156 P.n12 P.n11 1.705
R3157 P P.n17 0.616
R3158 P.n15 P.n14 0.301
R3159 P.n1 P.n0 0.108
R3160 P.n2 P.n1 0.108
R3161 P.n17 P.n2 0.108
R3162 P.n5 P.n4 0.03
R3163 P.n8 P.n7 0.026
R3164 P.n6 P.n3 0.023
R3165 P.n16 P.n12 0.023
R3166 P.n11 P.n10 0.021
R3167 P.n10 P.n9 0.014
R3168 P.n7 P.n6 0.003
R3169 P.n12 P.n8 0.003
R3170 P.n14 P.n13 0.001
R3171 net1_nand3.n1 net1_nand3.n0 13.361
R3172 net1_nand3.n86 net1_nand3.n85 13.361
R3173 net1_nand3.n11 net1_nand3.n9 9.3
R3174 net1_nand3.n5 net1_nand3.n3 9.3
R3175 net1_nand3.n16 net1_nand3.n13 9.3
R3176 net1_nand3.n148 net1_nand3.n140 9.3
R3177 net1_nand3.n148 net1_nand3.n147 9.3
R3178 net1_nand3.n22 net1_nand3.n20 9.3
R3179 net1_nand3.n33 net1_nand3.n31 9.3
R3180 net1_nand3.n30 net1_nand3.n28 9.3
R3181 net1_nand3.n41 net1_nand3.n39 9.3
R3182 net1_nand3.n41 net1_nand3.n40 9.3
R3183 net1_nand3.n52 net1_nand3.n50 9.3
R3184 net1_nand3.n52 net1_nand3.n51 9.3
R3185 net1_nand3.n63 net1_nand3.n61 9.3
R3186 net1_nand3.n63 net1_nand3.n62 9.3
R3187 net1_nand3.n74 net1_nand3.n72 9.3
R3188 net1_nand3.n74 net1_nand3.n73 9.3
R3189 net1_nand3.n98 net1_nand3.n96 9.3
R3190 net1_nand3.n98 net1_nand3.n97 9.3
R3191 net1_nand3.n109 net1_nand3.n107 9.3
R3192 net1_nand3.n109 net1_nand3.n108 9.3
R3193 net1_nand3.n120 net1_nand3.n118 9.3
R3194 net1_nand3.n120 net1_nand3.n119 9.3
R3195 net1_nand3.n167 net1_nand3.n129 9.3
R3196 net1_nand3.n167 net1_nand3.n166 9.3
R3197 net1_nand3.n160 net1_nand3.n133 9.3
R3198 net1_nand3.n160 net1_nand3.n159 9.3
R3199 net1_nand3.n27 net1_nand3.n24 9.3
R3200 net1_nand3.n33 net1_nand3.n32 9.3
R3201 net1_nand3.n38 net1_nand3.n35 9.3
R3202 net1_nand3.n44 net1_nand3.n42 9.3
R3203 net1_nand3.n49 net1_nand3.n46 9.3
R3204 net1_nand3.n55 net1_nand3.n53 9.3
R3205 net1_nand3.n60 net1_nand3.n57 9.3
R3206 net1_nand3.n66 net1_nand3.n64 9.3
R3207 net1_nand3.n71 net1_nand3.n68 9.3
R3208 net1_nand3.n77 net1_nand3.n75 9.3
R3209 net1_nand3.n82 net1_nand3.n79 9.3
R3210 net1_nand3.n92 net1_nand3.n89 9.3
R3211 net1_nand3.n95 net1_nand3.n93 9.3
R3212 net1_nand3.n103 net1_nand3.n100 9.3
R3213 net1_nand3.n106 net1_nand3.n104 9.3
R3214 net1_nand3.n114 net1_nand3.n111 9.3
R3215 net1_nand3.n117 net1_nand3.n115 9.3
R3216 net1_nand3.n127 net1_nand3.n123 9.3
R3217 net1_nand3.n169 net1_nand3.n128 9.3
R3218 net1_nand3.n165 net1_nand3.n131 9.3
R3219 net1_nand3.n162 net1_nand3.n132 9.3
R3220 net1_nand3.n158 net1_nand3.n135 9.3
R3221 net1_nand3.n155 net1_nand3.n136 9.3
R3222 net1_nand3.n151 net1_nand3.n139 9.3
R3223 net1_nand3.n153 net1_nand3.n137 9.3
R3224 net1_nand3.n38 net1_nand3.n37 9.3
R3225 net1_nand3.n44 net1_nand3.n43 9.3
R3226 net1_nand3.n49 net1_nand3.n48 9.3
R3227 net1_nand3.n55 net1_nand3.n54 9.3
R3228 net1_nand3.n60 net1_nand3.n59 9.3
R3229 net1_nand3.n66 net1_nand3.n65 9.3
R3230 net1_nand3.n71 net1_nand3.n70 9.3
R3231 net1_nand3.n77 net1_nand3.n76 9.3
R3232 net1_nand3.n82 net1_nand3.n81 9.3
R3233 net1_nand3.n92 net1_nand3.n91 9.3
R3234 net1_nand3.n95 net1_nand3.n94 9.3
R3235 net1_nand3.n103 net1_nand3.n102 9.3
R3236 net1_nand3.n106 net1_nand3.n105 9.3
R3237 net1_nand3.n114 net1_nand3.n113 9.3
R3238 net1_nand3.n117 net1_nand3.n116 9.3
R3239 net1_nand3.n127 net1_nand3.n126 9.3
R3240 net1_nand3.n169 net1_nand3.n168 9.3
R3241 net1_nand3.n165 net1_nand3.n164 9.3
R3242 net1_nand3.n162 net1_nand3.n161 9.3
R3243 net1_nand3.n158 net1_nand3.n157 9.3
R3244 net1_nand3.n155 net1_nand3.n154 9.3
R3245 net1_nand3.n151 net1_nand3.n150 9.3
R3246 net1_nand3.n153 net1_nand3.n152 9.3
R3247 net1_nand3.n30 net1_nand3.n29 9.3
R3248 net1_nand3.n27 net1_nand3.n26 9.3
R3249 net1_nand3.n22 net1_nand3.n21 9.3
R3250 net1_nand3.n19 net1_nand3.n17 9.3
R3251 net1_nand3.n19 net1_nand3.n18 9.3
R3252 net1_nand3.n16 net1_nand3.n15 9.3
R3253 net1_nand3.n144 net1_nand3.n142 9.3
R3254 net1_nand3.n146 net1_nand3.n141 9.3
R3255 net1_nand3.n146 net1_nand3.n145 9.3
R3256 net1_nand3.n144 net1_nand3.n143 9.3
R3257 net1_nand3.n11 net1_nand3.n10 9.3
R3258 net1_nand3.n8 net1_nand3.n6 9.3
R3259 net1_nand3.n8 net1_nand3.n7 9.3
R3260 net1_nand3.n5 net1_nand3.n4 9.3
R3261 net1_nand3.n122 net1_nand3.n121 8.043
R3262 net1_nand3.n125 net1_nand3.n124 8.043
R3263 net1_nand3.n84 net1_nand3.n2 4.558
R3264 net1_nand3.n87 net1_nand3.n1 4.558
R3265 net1_nand3.n84 net1_nand3.n83 4.558
R3266 net1_nand3.n87 net1_nand3.n86 4.558
R3267 net1_nand3.n124 net1_nand3.t1 2.9
R3268 net1_nand3.n121 net1_nand3.t0 2.9
R3269 net1_nand3.n79 net1_nand3.n78 0.536
R3270 net1_nand3.n89 net1_nand3.n88 0.536
R3271 net1_nand3.n81 net1_nand3.n80 0.536
R3272 net1_nand3.n91 net1_nand3.n90 0.536
R3273 net1_nand3.n70 net1_nand3.n69 0.506
R3274 net1_nand3.n102 net1_nand3.n101 0.506
R3275 net1_nand3.n68 net1_nand3.n67 0.506
R3276 net1_nand3.n100 net1_nand3.n99 0.506
R3277 net1_nand3.n57 net1_nand3.n56 0.475
R3278 net1_nand3.n111 net1_nand3.n110 0.475
R3279 net1_nand3.n59 net1_nand3.n58 0.475
R3280 net1_nand3.n113 net1_nand3.n112 0.475
R3281 net1_nand3.n126 net1_nand3.n125 0.445
R3282 net1_nand3.n46 net1_nand3.n45 0.445
R3283 net1_nand3.n123 net1_nand3.n122 0.445
R3284 net1_nand3.n48 net1_nand3.n47 0.445
R3285 net1_nand3.n35 net1_nand3.n34 0.413
R3286 net1_nand3.n131 net1_nand3.n130 0.413
R3287 net1_nand3.n37 net1_nand3.n36 0.413
R3288 net1_nand3.n164 net1_nand3.n163 0.413
R3289 net1_nand3.n26 net1_nand3.n25 0.382
R3290 net1_nand3.n157 net1_nand3.n156 0.382
R3291 net1_nand3.n135 net1_nand3.n134 0.382
R3292 net1_nand3.n24 net1_nand3.n23 0.382
R3293 net1_nand3.n13 net1_nand3.n12 0.349
R3294 net1_nand3.n15 net1_nand3.n14 0.349
R3295 net1_nand3.n139 net1_nand3.n138 0.349
R3296 net1_nand3.n150 net1_nand3.n149 0.349
R3297 net1_nand3.n87 net1_nand3.n84 0.055
R3298 net1_nand3.n16 net1_nand3.n11 0.041
R3299 net1_nand3.n27 net1_nand3.n22 0.041
R3300 net1_nand3.n38 net1_nand3.n33 0.041
R3301 net1_nand3.n49 net1_nand3.n44 0.041
R3302 net1_nand3.n60 net1_nand3.n55 0.041
R3303 net1_nand3.n71 net1_nand3.n66 0.041
R3304 net1_nand3.n82 net1_nand3.n77 0.041
R3305 net1_nand3.n95 net1_nand3.n92 0.041
R3306 net1_nand3.n106 net1_nand3.n103 0.041
R3307 net1_nand3.n117 net1_nand3.n114 0.041
R3308 net1_nand3.n165 net1_nand3.n162 0.041
R3309 net1_nand3.n158 net1_nand3.n155 0.041
R3310 net1_nand3.n151 net1_nand3.n148 0.041
R3311 net1_nand3 net1_nand3.n169 0.039
R3312 net1_nand3.n84 net1_nand3.n82 0.012
R3313 net1_nand3.n92 net1_nand3.n87 0.012
R3314 net1_nand3.n11 net1_nand3.n8 0.011
R3315 net1_nand3.n74 net1_nand3.n71 0.011
R3316 net1_nand3.n103 net1_nand3.n98 0.011
R3317 net1_nand3.n148 net1_nand3.n146 0.011
R3318 net1_nand3.n22 net1_nand3.n19 0.01
R3319 net1_nand3.n155 net1_nand3.n153 0.01
R3320 net1_nand3.n63 net1_nand3.n60 0.009
R3321 net1_nand3.n114 net1_nand3.n109 0.009
R3322 net1_nand3.n33 net1_nand3.n30 0.008
R3323 net1_nand3.n162 net1_nand3.n160 0.008
R3324 net1_nand3.n44 net1_nand3.n41 0.007
R3325 net1_nand3.n52 net1_nand3.n49 0.007
R3326 net1_nand3.n127 net1_nand3.n120 0.007
R3327 net1_nand3.n169 net1_nand3.n167 0.007
R3328 net1_nand3.n41 net1_nand3.n38 0.006
R3329 net1_nand3.n167 net1_nand3.n165 0.006
R3330 net1_nand3.n55 net1_nand3.n52 0.005
R3331 net1_nand3.n120 net1_nand3.n117 0.005
R3332 net1_nand3.n30 net1_nand3.n27 0.004
R3333 net1_nand3.n160 net1_nand3.n158 0.004
R3334 net1_nand3.n19 net1_nand3.n16 0.003
R3335 net1_nand3.n66 net1_nand3.n63 0.003
R3336 net1_nand3.n109 net1_nand3.n106 0.003
R3337 net1_nand3.n153 net1_nand3.n151 0.003
R3338 net1_nand3.n77 net1_nand3.n74 0.002
R3339 net1_nand3.n98 net1_nand3.n95 0.002
R3340 net1_nand3 net1_nand3.n127 0.002
R3341 net1_nand3.n8 net1_nand3.n5 0.001
R3342 net1_nand3.n146 net1_nand3.n144 0.001
R3343 net3_ff2.n257 net3_ff2.t3 735.052
R3344 net3_ff2.n87 net3_ff2.t2 399.297
R3345 net3_ff2.n32 net3_ff2.n31 92.5
R3346 net3_ff2.n47 net3_ff2.n46 92.5
R3347 net3_ff2.n46 net3_ff2.t0 70.344
R3348 net3_ff2.n10 net3_ff2.n9 31.034
R3349 net3_ff2.n66 net3_ff2.n65 31.034
R3350 net3_ff2.n216 net3_ff2.n215 9.3
R3351 net3_ff2.n106 net3_ff2.n105 9.3
R3352 net3_ff2.n18 net3_ff2.n17 9.3
R3353 net3_ff2.n67 net3_ff2.n66 9.3
R3354 net3_ff2.n11 net3_ff2.n10 9.3
R3355 net3_ff2.n77 net3_ff2.n76 9.3
R3356 net3_ff2.n174 net3_ff2.n173 9.154
R3357 net3_ff2.n33 net3_ff2.n32 8.282
R3358 net3_ff2.n48 net3_ff2.n47 8.282
R3359 net3_ff2.n173 net3_ff2.t1 7.141
R3360 net3_ff2.n99 net3_ff2.n98 7.033
R3361 net3_ff2.n93 net3_ff2.n92 7.033
R3362 net3_ff2.n11 net3_ff2.n7 5.647
R3363 net3_ff2.n67 net3_ff2.n63 5.647
R3364 net3_ff2.n175 net3_ff2.n174 4.65
R3365 net3_ff2.n45 net3_ff2.n44 4.65
R3366 net3_ff2.n134 net3_ff2.n133 4.5
R3367 net3_ff2.n112 net3_ff2.n111 4.5
R3368 net3_ff2.n155 net3_ff2.n154 4.5
R3369 net3_ff2.n162 net3_ff2.n159 4.5
R3370 net3_ff2.n170 net3_ff2.n169 4.5
R3371 net3_ff2.n176 net3_ff2.n172 4.5
R3372 net3_ff2.n203 net3_ff2.n200 4.5
R3373 net3_ff2.n210 net3_ff2.n209 4.5
R3374 net3_ff2.n222 net3_ff2.n221 4.5
R3375 net3_ff2.n232 net3_ff2.n231 4.5
R3376 net3_ff2.n242 net3_ff2.n241 4.5
R3377 net3_ff2.n122 net3_ff2.n121 4.5
R3378 net3_ff2.n83 net3_ff2.n81 4.5
R3379 net3_ff2.n71 net3_ff2.n68 4.5
R3380 net3_ff2.n58 net3_ff2.n56 4.5
R3381 net3_ff2.n34 net3_ff2.n33 4.5
R3382 net3_ff2.n41 net3_ff2.n40 4.5
R3383 net3_ff2.n49 net3_ff2.n48 4.5
R3384 net3_ff2.n14 net3_ff2.n13 4.5
R3385 net3_ff2.n23 net3_ff2.n22 4.5
R3386 net3_ff2.n231 net3_ff2.n228 4.141
R3387 net3_ff2.n121 net3_ff2.n120 4.141
R3388 net3_ff2.n9 net3_ff2.n8 4.137
R3389 net3_ff2.n65 net3_ff2.n64 4.137
R3390 net3_ff2.n221 net3_ff2.n218 3.764
R3391 net3_ff2.n154 net3_ff2.n152 3.764
R3392 net3_ff2.n22 net3_ff2.n20 3.764
R3393 net3_ff2.n68 net3_ff2.n61 3.764
R3394 net3_ff2.n241 net3_ff2.n238 3.388
R3395 net3_ff2.n209 net3_ff2.n208 3.388
R3396 net3_ff2.n111 net3_ff2.n110 3.388
R3397 net3_ff2.n133 net3_ff2.n132 3.388
R3398 net3_ff2.n13 net3_ff2.n12 3.388
R3399 net3_ff2.n81 net3_ff2.n80 3.388
R3400 net3_ff2.n241 net3_ff2.n240 3.011
R3401 net3_ff2.n209 net3_ff2.n206 3.011
R3402 net3_ff2.n200 net3_ff2.n198 3.011
R3403 net3_ff2.n105 net3_ff2.n104 3.011
R3404 net3_ff2.n111 net3_ff2.n109 3.011
R3405 net3_ff2.n133 net3_ff2.n131 3.011
R3406 net3_ff2.n13 net3_ff2.n11 3.011
R3407 net3_ff2.n33 net3_ff2.n30 3.011
R3408 net3_ff2.n81 net3_ff2.n79 3.011
R3409 net3_ff2.n221 net3_ff2.n220 2.635
R3410 net3_ff2.n215 net3_ff2.n214 2.635
R3411 net3_ff2.n159 net3_ff2.n158 2.635
R3412 net3_ff2.n154 net3_ff2.n153 2.635
R3413 net3_ff2.n22 net3_ff2.n21 2.635
R3414 net3_ff2.n56 net3_ff2.n55 2.635
R3415 net3_ff2.n68 net3_ff2.n67 2.635
R3416 net3_ff2.n231 net3_ff2.n230 2.258
R3417 net3_ff2.n121 net3_ff2.n119 2.258
R3418 net3_ff2.n86 net3_ff2.n85 1.705
R3419 net3_ff2.n256 net3_ff2.n247 1.705
R3420 net3_ff2 net3_ff2.n87 1.689
R3421 net3_ff2.n159 net3_ff2.n157 1.505
R3422 net3_ff2.n156 net3_ff2.n155 1.5
R3423 net3_ff2.n163 net3_ff2.n162 1.5
R3424 net3_ff2.n171 net3_ff2.n170 1.5
R3425 net3_ff2.n177 net3_ff2.n176 1.5
R3426 net3_ff2.n84 net3_ff2.n83 1.5
R3427 net3_ff2.n72 net3_ff2.n71 1.5
R3428 net3_ff2.n35 net3_ff2.n34 1.5
R3429 net3_ff2.n59 net3_ff2.n58 1.5
R3430 net3_ff2.n42 net3_ff2.n41 1.5
R3431 net3_ff2.n50 net3_ff2.n49 1.5
R3432 net3_ff2.n27 net3_ff2.n14 1.5
R3433 net3_ff2.n24 net3_ff2.n23 1.5
R3434 net3_ff2.n200 net3_ff2.n199 1.129
R3435 net3_ff2.n100 net3_ff2.n99 1.127
R3436 net3_ff2.n247 net3_ff2.n93 1.127
R3437 net3_ff2.n243 net3_ff2.n242 1.125
R3438 net3_ff2.n135 net3_ff2.n134 1.125
R3439 net3_ff2.n7 net3_ff2.n6 0.752
R3440 net3_ff2.n63 net3_ff2.n62 0.752
R3441 net3_ff2.n92 net3_ff2.n91 0.155
R3442 net3_ff2.n98 net3_ff2.n97 0.155
R3443 net3_ff2.n240 net3_ff2.n239 0.144
R3444 net3_ff2.n131 net3_ff2.n130 0.144
R3445 net3_ff2.n230 net3_ff2.n229 0.133
R3446 net3_ff2.n119 net3_ff2.n118 0.132
R3447 net3_ff2.n87 net3_ff2.n86 0.117
R3448 net3_ff2.n257 net3_ff2.n256 0.112
R3449 net3_ff2 net3_ff2.n257 0.085
R3450 net3_ff2.n236 net3_ff2.n235 0.053
R3451 net3_ff2.n226 net3_ff2.n225 0.053
R3452 net3_ff2.n216 net3_ff2.n213 0.053
R3453 net3_ff2.n116 net3_ff2.n115 0.053
R3454 net3_ff2.n126 net3_ff2.n125 0.053
R3455 net3_ff2.n77 net3_ff2.n75 0.053
R3456 net3_ff2.n1 net3_ff2.n0 0.05
R3457 net3_ff2.n2 net3_ff2.n1 0.05
R3458 net3_ff2.n86 net3_ff2.n2 0.05
R3459 net3_ff2.n256 net3_ff2.n255 0.05
R3460 net3_ff2.n255 net3_ff2.n254 0.05
R3461 net3_ff2.n254 net3_ff2.n253 0.05
R3462 net3_ff2.n253 net3_ff2.n252 0.05
R3463 net3_ff2.n252 net3_ff2.n251 0.05
R3464 net3_ff2.n251 net3_ff2.n250 0.05
R3465 net3_ff2.n250 net3_ff2.n249 0.05
R3466 net3_ff2.n249 net3_ff2.n248 0.05
R3467 net3_ff2.n41 net3_ff2.n39 0.045
R3468 net3_ff2.n58 net3_ff2.n54 0.045
R3469 net3_ff2.n203 net3_ff2.n202 0.043
R3470 net3_ff2.n170 net3_ff2.n168 0.043
R3471 net3_ff2.n89 net3_ff2.n88 0.034
R3472 net3_ff2.n125 net3_ff2.n124 0.032
R3473 net3_ff2.n95 net3_ff2.n94 0.032
R3474 net3_ff2.n237 net3_ff2.n236 0.03
R3475 net3_ff2.n235 net3_ff2.n234 0.03
R3476 net3_ff2.n115 net3_ff2.n114 0.03
R3477 net3_ff2.n225 net3_ff2.n224 0.028
R3478 net3_ff2.n127 net3_ff2.n126 0.028
R3479 net3_ff2.n129 net3_ff2.n128 0.028
R3480 net3_ff2.n25 net3_ff2.n24 0.027
R3481 net3_ff2.n84 net3_ff2.n74 0.027
R3482 net3_ff2.n197 net3_ff2.n196 0.025
R3483 net3_ff2.n227 net3_ff2.n226 0.025
R3484 net3_ff2.n49 net3_ff2.n45 0.025
R3485 net3_ff2.n220 net3_ff2.n219 0.024
R3486 net3_ff2.n109 net3_ff2.n108 0.024
R3487 net3_ff2.n176 net3_ff2.n175 0.023
R3488 net3_ff2.n117 net3_ff2.n116 0.023
R3489 net3_ff2.n223 net3_ff2.n222 0.021
R3490 net3_ff2.n217 net3_ff2.n216 0.021
R3491 net3_ff2.n149 net3_ff2.n148 0.021
R3492 net3_ff2.n23 net3_ff2.n16 0.021
R3493 net3_ff2.n19 net3_ff2.n18 0.021
R3494 net3_ff2.n71 net3_ff2.n60 0.021
R3495 net3_ff2.n242 net3_ff2.n197 0.019
R3496 net3_ff2.n213 net3_ff2.n212 0.019
R3497 net3_ff2.n212 net3_ff2.n211 0.019
R3498 net3_ff2.n210 net3_ff2.n205 0.019
R3499 net3_ff2.n150 net3_ff2.n149 0.019
R3500 net3_ff2.n107 net3_ff2.n106 0.019
R3501 net3_ff2.n113 net3_ff2.n112 0.019
R3502 net3_ff2.n134 net3_ff2.n129 0.019
R3503 net3_ff2.n4 net3_ff2.n3 0.019
R3504 net3_ff2.n5 net3_ff2.n4 0.019
R3505 net3_ff2.n70 net3_ff2.n69 0.019
R3506 net3_ff2.n78 net3_ff2.n77 0.019
R3507 net3_ff2.n83 net3_ff2.n82 0.019
R3508 net3_ff2.n93 net3_ff2.n90 0.019
R3509 net3_ff2.n99 net3_ff2.n96 0.019
R3510 net3_ff2.n242 net3_ff2.n237 0.017
R3511 net3_ff2.n233 net3_ff2.n232 0.017
R3512 net3_ff2.n211 net3_ff2.n210 0.017
R3513 net3_ff2.n204 net3_ff2.n203 0.017
R3514 net3_ff2.n112 net3_ff2.n107 0.017
R3515 net3_ff2.n123 net3_ff2.n122 0.017
R3516 net3_ff2.n134 net3_ff2.n127 0.017
R3517 net3_ff2.n14 net3_ff2.n5 0.017
R3518 net3_ff2.n34 net3_ff2.n29 0.017
R3519 net3_ff2.n83 net3_ff2.n78 0.017
R3520 net3_ff2.n186 net3_ff2.n185 0.016
R3521 net3_ff2.n145 net3_ff2.n144 0.016
R3522 net3_ff2.n222 net3_ff2.n217 0.015
R3523 net3_ff2.n162 net3_ff2.n161 0.015
R3524 net3_ff2.n155 net3_ff2.n150 0.015
R3525 net3_ff2.n23 net3_ff2.n19 0.015
R3526 net3_ff2.n58 net3_ff2.n57 0.015
R3527 net3_ff2.n71 net3_ff2.n70 0.015
R3528 net3_ff2.n245 net3_ff2.n244 0.014
R3529 net3_ff2.n194 net3_ff2.n193 0.014
R3530 net3_ff2.n189 net3_ff2.n188 0.014
R3531 net3_ff2.n142 net3_ff2.n141 0.014
R3532 net3_ff2.n138 net3_ff2.n137 0.014
R3533 net3_ff2.n103 net3_ff2.n102 0.014
R3534 net3_ff2.n35 net3_ff2.n27 0.014
R3535 net3_ff2.n72 net3_ff2.n59 0.014
R3536 net3_ff2.n182 net3_ff2.n181 0.013
R3537 net3_ff2.n177 net3_ff2.n171 0.013
R3538 net3_ff2.n163 net3_ff2.n156 0.013
R3539 net3_ff2.n135 net3_ff2.n103 0.013
R3540 net3_ff2.n36 net3_ff2.n35 0.013
R3541 net3_ff2.n42 net3_ff2.n37 0.013
R3542 net3_ff2.n51 net3_ff2.n50 0.013
R3543 net3_ff2.n59 net3_ff2.n52 0.013
R3544 net3_ff2.n208 net3_ff2.n207 0.012
R3545 net3_ff2.n152 net3_ff2.n151 0.012
R3546 net3_ff2.n232 net3_ff2.n227 0.012
R3547 net3_ff2.n205 net3_ff2.n204 0.012
R3548 net3_ff2.n161 net3_ff2.n160 0.012
R3549 net3_ff2.n122 net3_ff2.n117 0.012
R3550 net3_ff2.n244 net3_ff2.n243 0.012
R3551 net3_ff2.n178 net3_ff2.n177 0.012
R3552 net3_ff2.n29 net3_ff2.n28 0.012
R3553 net3_ff2.n171 net3_ff2.n166 0.011
R3554 net3_ff2.n246 net3_ff2.n245 0.01
R3555 net3_ff2.n193 net3_ff2.n192 0.01
R3556 net3_ff2.n183 net3_ff2.n182 0.01
R3557 net3_ff2.n164 net3_ff2.n163 0.01
R3558 net3_ff2.n139 net3_ff2.n138 0.01
R3559 net3_ff2.n102 net3_ff2.n101 0.01
R3560 net3_ff2.n27 net3_ff2.n26 0.01
R3561 net3_ff2.n73 net3_ff2.n72 0.01
R3562 net3_ff2.n191 net3_ff2.n190 0.009
R3563 net3_ff2.n181 net3_ff2.n180 0.009
R3564 net3_ff2.n156 net3_ff2.n147 0.009
R3565 net3_ff2.n141 net3_ff2.n140 0.009
R3566 net3_ff2.n202 net3_ff2.n201 0.008
R3567 net3_ff2.n168 net3_ff2.n167 0.008
R3568 net3_ff2.n195 net3_ff2.n194 0.008
R3569 net3_ff2.n185 net3_ff2.n184 0.008
R3570 net3_ff2.n146 net3_ff2.n145 0.008
R3571 net3_ff2.n143 net3_ff2.n142 0.008
R3572 net3_ff2.n39 net3_ff2.n38 0.008
R3573 net3_ff2.n54 net3_ff2.n53 0.008
R3574 net3_ff2.n24 net3_ff2.n15 0.008
R3575 net3_ff2.n188 net3_ff2.n187 0.007
R3576 net3_ff2.n187 net3_ff2.n186 0.007
R3577 net3_ff2.n144 net3_ff2.n143 0.007
R3578 net3_ff2.n137 net3_ff2.n136 0.007
R3579 net3_ff2.n43 net3_ff2.n42 0.007
R3580 net3_ff2.n50 net3_ff2.n43 0.007
R3581 net3_ff2.n85 net3_ff2.n84 0.007
R3582 net3_ff2.n234 net3_ff2.n233 0.006
R3583 net3_ff2.n224 net3_ff2.n223 0.006
R3584 net3_ff2.n114 net3_ff2.n113 0.006
R3585 net3_ff2.n124 net3_ff2.n123 0.006
R3586 net3_ff2.n74 net3_ff2.n73 0.006
R3587 net3_ff2.n184 net3_ff2.n183 0.005
R3588 net3_ff2.n147 net3_ff2.n146 0.005
R3589 net3_ff2.n26 net3_ff2.n25 0.005
R3590 net3_ff2.n90 net3_ff2.n89 0.004
R3591 net3_ff2.n96 net3_ff2.n95 0.004
R3592 net3_ff2.n247 net3_ff2.n246 0.004
R3593 net3_ff2.n243 net3_ff2.n195 0.004
R3594 net3_ff2.n192 net3_ff2.n191 0.004
R3595 net3_ff2.n140 net3_ff2.n139 0.004
R3596 net3_ff2.n136 net3_ff2.n135 0.004
R3597 net3_ff2.n101 net3_ff2.n100 0.004
R3598 net3_ff2.n180 net3_ff2.n179 0.002
R3599 net3_ff2.n179 net3_ff2.n178 0.002
R3600 net3_ff2.n166 net3_ff2.n165 0.002
R3601 net3_ff2.n165 net3_ff2.n164 0.002
R3602 net3_ff2.n37 net3_ff2.n36 0.002
R3603 net3_ff2.n52 net3_ff2.n51 0.002
R3604 net3_ff2.n190 net3_ff2.n189 0.001
R3605 net5_ff2.n35 net5_ff2.n34 92.5
R3606 net5_ff2.n33 net5_ff2.n32 92.5
R3607 net5_ff2.n28 net5_ff2.n27 92.5
R3608 net5_ff2.n30 net5_ff2.n29 92.5
R3609 net5_ff2.n32 net5_ff2.t1 70.344
R3610 net5_ff2.n27 net5_ff2.t0 70.344
R3611 net5_ff2.n17 net5_ff2.n16 31.034
R3612 net5_ff2.n58 net5_ff2.n57 31.034
R3613 net5_ff2.n23 net5_ff2.n22 31.034
R3614 net5_ff2.n43 net5_ff2.n42 31.034
R3615 net5_ff2.n36 net5_ff2.n33 12.8
R3616 net5_ff2.n36 net5_ff2.n35 12.8
R3617 net5_ff2.n31 net5_ff2.n28 12.8
R3618 net5_ff2.n31 net5_ff2.n30 12.8
R3619 net5_ff2.n12 net5_ff2.n10 9.3
R3620 net5_ff2.n6 net5_ff2.n4 9.3
R3621 net5_ff2.n25 net5_ff2.n18 9.3
R3622 net5_ff2.n18 net5_ff2.n17 9.3
R3623 net5_ff2.n53 net5_ff2.n45 9.3
R3624 net5_ff2.n53 net5_ff2.n52 9.3
R3625 net5_ff2.n60 net5_ff2.n44 9.3
R3626 net5_ff2.n44 net5_ff2.n43 9.3
R3627 net5_ff2.n60 net5_ff2.n59 9.3
R3628 net5_ff2.n59 net5_ff2.n58 9.3
R3629 net5_ff2.n25 net5_ff2.n24 9.3
R3630 net5_ff2.n24 net5_ff2.n23 9.3
R3631 net5_ff2.n49 net5_ff2.n47 9.3
R3632 net5_ff2.n51 net5_ff2.n46 9.3
R3633 net5_ff2.n51 net5_ff2.n50 9.3
R3634 net5_ff2.n49 net5_ff2.n48 9.3
R3635 net5_ff2.n12 net5_ff2.n11 9.3
R3636 net5_ff2.n9 net5_ff2.n7 9.3
R3637 net5_ff2.n9 net5_ff2.n8 9.3
R3638 net5_ff2.n6 net5_ff2.n5 9.3
R3639 net5_ff2.n18 net5_ff2.n14 5.647
R3640 net5_ff2.n59 net5_ff2.n55 5.647
R3641 net5_ff2.n24 net5_ff2.n20 5.647
R3642 net5_ff2.n44 net5_ff2.n40 5.647
R3643 net5_ff2.n37 net5_ff2.n31 4.65
R3644 net5_ff2.n37 net5_ff2.n36 4.65
R3645 net5_ff2.n26 net5_ff2.n3 4.47
R3646 net5_ff2.n38 net5_ff2.n1 4.47
R3647 net5_ff2.n38 net5_ff2.n0 4.47
R3648 net5_ff2.n26 net5_ff2.n2 4.47
R3649 net5_ff2.n16 net5_ff2.n15 4.137
R3650 net5_ff2.n57 net5_ff2.n56 4.137
R3651 net5_ff2.n22 net5_ff2.n21 4.137
R3652 net5_ff2.n42 net5_ff2.n41 4.137
R3653 net5_ff2.n14 net5_ff2.n13 0.752
R3654 net5_ff2.n55 net5_ff2.n54 0.752
R3655 net5_ff2.n20 net5_ff2.n19 0.752
R3656 net5_ff2.n40 net5_ff2.n39 0.752
R3657 net5_ff2.n37 net5_ff2.n26 0.032
R3658 net5_ff2.n38 net5_ff2.n37 0.032
R3659 net5_ff2.n25 net5_ff2.n12 0.024
R3660 net5_ff2.n60 net5_ff2.n53 0.024
R3661 net5_ff2.n26 net5_ff2.n25 0.007
R3662 net5_ff2.n9 net5_ff2.n6 0.006
R3663 net5_ff2.n51 net5_ff2.n49 0.006
R3664 net5_ff2 net5_ff2.n38 0.005
R3665 net5_ff2.n12 net5_ff2.n9 0.001
R3666 net5_ff2 net5_ff2.n60 0.001
R3667 net5_ff2.n53 net5_ff2.n51 0.001
R3668 3.n354 3.t2 732.452
R3669 3.n354 3.t3 397.573
R3670 3.n252 3.n251 92.5
R3671 3.n315 3.n314 92.5
R3672 3.n251 3.t1 70.344
R3673 3.n265 3.n264 31.034
R3674 3.n332 3.n331 31.034
R3675 3.n275 3.n274 9.3
R3676 3.n341 3.n340 9.3
R3677 3.n333 3.n332 9.3
R3678 3.n266 3.n265 9.3
R3679 3.n62 3.n61 9.3
R3680 3.n164 3.n163 9.3
R3681 3.n128 3.n127 9.154
R3682 3.n253 3.n252 8.282
R3683 3.n316 3.n315 8.282
R3684 3.n127 3.t0 7.141
R3685 3.n222 3.n221 7.03
R3686 3.n5 3.n4 7.03
R3687 3.n266 3.n262 5.647
R3688 3.n333 3.n329 5.647
R3689 3.n313 3.n312 4.65
R3690 3.n129 3.n128 4.65
R3691 3.n353 3.n352 4.569
R3692 3.n317 3.n316 4.5
R3693 3.n324 3.n323 4.5
R3694 3.n258 3.n253 4.5
R3695 3.n335 3.n334 4.5
R3696 3.n311 3.n310 4.5
R3697 3.n269 3.n268 4.5
R3698 3.n347 3.n345 4.5
R3699 3.n280 3.n279 4.5
R3700 3.n28 3.n22 4.5
R3701 3.n167 3.n159 4.5
R3702 3.n189 3.n183 4.5
R3703 3.n146 3.n145 4.5
R3704 3.n116 3.n113 4.5
R3705 3.n131 3.n125 4.5
R3706 3.n105 3.n93 4.5
R3707 3.n121 3.n120 4.5
R3708 3.n102 3.n97 4.5
R3709 3.n73 3.n72 4.5
R3710 3.n47 3.n43 4.5
R3711 3.n210 3.n209 4.5
R3712 3.n353 3.n236 4.483
R3713 3.n183 3.n180 4.141
R3714 3.n43 3.n42 4.141
R3715 3.n264 3.n263 4.137
R3716 3.n331 3.n330 4.137
R3717 3.n279 3.n277 3.764
R3718 3.n334 3.n327 3.764
R3719 3.n159 3.n156 3.764
R3720 3.n97 3.n95 3.764
R3721 3.n268 3.n267 3.388
R3722 3.n345 3.n344 3.388
R3723 3.n209 3.n206 3.388
R3724 3.n145 3.n144 3.388
R3725 3.n72 3.n71 3.388
R3726 3.n22 3.n21 3.388
R3727 3.n268 3.n266 3.011
R3728 3.n253 3.n250 3.011
R3729 3.n345 3.n343 3.011
R3730 3.n209 3.n208 3.011
R3731 3.n145 3.n142 3.011
R3732 3.n113 3.n111 3.011
R3733 3.n61 3.n60 3.011
R3734 3.n72 3.n70 3.011
R3735 3.n22 3.n20 3.011
R3736 3.n279 3.n278 2.635
R3737 3.n323 3.n322 2.635
R3738 3.n334 3.n333 2.635
R3739 3.n159 3.n158 2.635
R3740 3.n163 3.n162 2.635
R3741 3.n93 3.n92 2.635
R3742 3.n97 3.n96 2.635
R3743 3.n183 3.n182 2.258
R3744 3.n43 3.n41 2.258
R3745 3.n93 3.n91 1.505
R3746 3.n348 3.n347 1.5
R3747 3.n281 3.n280 1.5
R3748 3.n8 3.n6 1.5
R3749 3.n29 3.n28 1.5
R3750 3.n190 3.n189 1.5
R3751 3.n228 3.n227 1.5
R3752 3.n168 3.n167 1.5
R3753 3.n147 3.n146 1.5
R3754 3.n117 3.n116 1.5
R3755 3.n132 3.n131 1.5
R3756 3.n106 3.n105 1.5
R3757 3.n122 3.n121 1.5
R3758 3.n74 3.n73 1.5
R3759 3.n48 3.n47 1.5
R3760 3.n211 3.n210 1.5
R3761 3 3.n353 1.297
R3762 3.n10 3.n9 1.137
R3763 3.n31 3.n30 1.137
R3764 3.n50 3.n49 1.137
R3765 3.n58 3.n57 1.137
R3766 3.n76 3.n75 1.137
R3767 3.n83 3.n82 1.137
R3768 3.n176 3.n175 1.137
R3769 3.n234 3.n233 1.137
R3770 3.n195 3.n194 1.137
R3771 3.n151 3.n150 1.137
R3772 3.n172 3.n171 1.137
R3773 3.n134 3.n133 1.137
R3774 3.n110 3.n109 1.137
R3775 3.n218 3.n217 1.137
R3776 3.n113 3.n112 1.129
R3777 3 3.n354 1.057
R3778 3.n351 3.n350 0.853
R3779 3.n262 3.n261 0.752
R3780 3.n329 3.n328 0.752
R3781 3.n283 3.n282 0.704
R3782 3.n221 3.n220 0.155
R3783 3.n4 3.n3 0.155
R3784 3.n208 3.n207 0.144
R3785 3.n20 3.n19 0.144
R3786 3.n182 3.n181 0.133
R3787 3.n41 3.n40 0.132
R3788 3.n234 3.n218 0.049
R3789 3.n134 3.n110 0.049
R3790 3.n31 3.n10 0.049
R3791 3.n203 3.n202 0.047
R3792 3.n149 3.n148 0.045
R3793 3.n133 3.n132 0.045
R3794 3.n164 3.n161 0.043
R3795 3.n48 3.n36 0.043
R3796 3.n29 3.n15 0.041
R3797 3.n105 3.n90 0.039
R3798 3.n233 3.n232 0.039
R3799 3.n116 3.n115 0.037
R3800 3.n9 3.n0 0.037
R3801 3.n255 3.n254 0.035
R3802 3.n319 3.n318 0.035
R3803 3.n238 3.n237 0.035
R3804 3.n300 3.n299 0.035
R3805 3.n186 3.n185 0.035
R3806 3.n100 3.n99 0.035
R3807 3.n248 3.n247 0.034
R3808 3.n309 3.n308 0.034
R3809 3.n25 3.n24 0.034
R3810 3.n231 3.n230 0.034
R3811 3.n124 3.n123 0.034
R3812 3.n14 3.n13 0.034
R3813 3.n338 3.n337 0.032
R3814 3.n307 3.n306 0.032
R3815 3.n228 3.n219 0.032
R3816 3.n107 3.n106 0.032
R3817 3.n88 3.n87 0.032
R3818 3.n284 3.n283 0.031
R3819 3.n295 3.n294 0.031
R3820 3.n196 3.n195 0.031
R3821 3.n151 3.n136 0.031
R3822 3.n84 3.n83 0.031
R3823 3.n50 3.n33 0.031
R3824 3.n272 3.n271 0.03
R3825 3.n341 3.n339 0.03
R3826 3.n246 3.n245 0.03
R3827 3.n305 3.n304 0.03
R3828 3.n225 3.n224 0.03
R3829 3.n214 3.n213 0.03
R3830 3.n147 3.n137 0.03
R3831 3.n118 3.n117 0.03
R3832 3.n275 3.n273 0.028
R3833 3.n257 3.n256 0.028
R3834 3.n321 3.n320 0.028
R3835 3.n243 3.n242 0.028
R3836 3.n240 3.n239 0.028
R3837 3.n302 3.n301 0.028
R3838 3.n348 3.n309 0.028
R3839 3.n35 3.n34 0.028
R3840 3.n282 3.n281 0.027
R3841 3.n288 3.n287 0.027
R3842 3.n291 3.n290 0.027
R3843 3.n176 3.n172 0.027
R3844 3.n76 3.n58 0.027
R3845 3.n281 3.n248 0.026
R3846 3.n204 3.n203 0.026
R3847 3.n67 3.n66 0.026
R3848 3.n216 3.n215 0.026
R3849 3.n17 3.n16 0.024
R3850 3.n27 3.n26 0.024
R3851 3.n194 3.n193 0.024
R3852 3.n174 3.n173 0.024
R3853 3.n171 3.n170 0.024
R3854 3.n82 3.n81 0.024
R3855 3.n57 3.n56 0.024
R3856 3.n12 3.n11 0.024
R3857 3.n158 3.n157 0.024
R3858 3.n70 3.n69 0.024
R3859 3.n317 3.n313 0.022
R3860 3.n298 3.n297 0.022
R3861 3.n350 3.n348 0.022
R3862 3.n200 3.n199 0.022
R3863 3.n187 3.n186 0.022
R3864 3.n46 3.n45 0.022
R3865 3.n74 3.n59 0.022
R3866 3.n313 3.n311 0.02
R3867 3.n297 3.n296 0.02
R3868 3.n189 3.n179 0.02
R3869 3.n38 3.n37 0.02
R3870 3.n47 3.n46 0.02
R3871 3.n351 3.n295 0.019
R3872 3.n352 3.n351 0.019
R3873 3.n280 3.n249 0.018
R3874 3.n276 3.n275 0.018
R3875 3.n273 3.n272 0.018
R3876 3.n335 3.n326 0.018
R3877 3.n247 3.n246 0.018
R3878 3.n167 3.n155 0.018
R3879 3.n165 3.n164 0.018
R3880 3.n103 3.n102 0.018
R3881 3.n8 3.n7 0.017
R3882 3.n269 3.n260 0.017
R3883 3.n339 3.n338 0.017
R3884 3.n342 3.n341 0.017
R3885 3.n347 3.n346 0.017
R3886 3.n245 3.n244 0.017
R3887 3.n306 3.n305 0.017
R3888 3.n308 3.n307 0.017
R3889 3.n210 3.n200 0.017
R3890 3.n146 3.n141 0.017
R3891 3.n130 3.n129 0.017
R3892 3.n129 3.n126 0.017
R3893 3.n63 3.n62 0.017
R3894 3.n73 3.n68 0.017
R3895 3.n28 3.n27 0.017
R3896 3.n215 3.n214 0.017
R3897 3.n236 3.n235 0.016
R3898 3.n197 3.n196 0.016
R3899 3.n136 3.n135 0.016
R3900 3.n85 3.n84 0.016
R3901 3.n33 3.n32 0.016
R3902 3.n270 3.n269 0.015
R3903 3.n259 3.n258 0.015
R3904 3.n347 3.n342 0.015
R3905 3.n242 3.n241 0.015
R3906 3.n170 3.n169 0.015
R3907 3.n81 3.n80 0.015
R3908 3.n280 3.n276 0.013
R3909 3.n325 3.n324 0.013
R3910 3.n336 3.n335 0.013
R3911 3.n304 3.n303 0.013
R3912 3.n105 3.n104 0.013
R3913 3.n73 3.n64 0.013
R3914 3.n75 3.n74 0.013
R3915 3.n56 3.n55 0.013
R3916 3.n144 3.n143 0.012
R3917 3.n95 3.n94 0.012
R3918 3.n289 3.n288 0.012
R3919 3.n290 3.n289 0.012
R3920 3.n350 3.n349 0.012
R3921 3.n260 3.n259 0.011
R3922 3.n326 3.n325 0.011
R3923 3.n286 3.n285 0.011
R3924 3.n293 3.n292 0.011
R3925 3.n185 3.n184 0.011
R3926 3.n167 3.n166 0.011
R3927 3.n139 3.n138 0.011
R3928 3.n141 3.n140 0.011
R3929 3.n104 3.n103 0.011
R3930 3.n101 3.n100 0.011
R3931 3.n24 3.n23 0.011
R3932 3.n192 3.n191 0.011
R3933 3.n175 3.n174 0.011
R3934 3.n171 3.n168 0.011
R3935 3.n106 3.n88 0.011
R3936 3.n318 3.n317 0.009
R3937 3.n299 3.n298 0.009
R3938 3.n227 3.n226 0.009
R3939 3.n226 3.n225 0.009
R3940 3.n224 3.n223 0.009
R3941 3.n205 3.n204 0.009
R3942 3.n66 3.n65 0.009
R3943 3.n18 3.n17 0.009
R3944 3.n2 3.n1 0.009
R3945 3.n6 3.n2 0.009
R3946 3.n233 3.n228 0.009
R3947 3.n232 3.n231 0.009
R3948 3.n217 3.n216 0.009
R3949 3.n57 3.n53 0.009
R3950 3.n30 3.n12 0.009
R3951 3.n9 3.n8 0.009
R3952 3.n195 3.n178 0.009
R3953 3.n177 3.n176 0.009
R3954 3.n172 3.n153 0.009
R3955 3.n152 3.n151 0.009
R3956 3.n83 3.n78 0.009
R3957 3.n77 3.n76 0.009
R3958 3.n58 3.n52 0.009
R3959 3.n51 3.n50 0.009
R3960 3.n256 3.n255 0.007
R3961 3.n320 3.n319 0.007
R3962 3.n239 3.n238 0.007
R3963 3.n301 3.n300 0.007
R3964 3.n119 3.n118 0.007
R3965 3.n108 3.n107 0.007
R3966 3.n285 3.n284 0.006
R3967 3.n287 3.n286 0.006
R3968 3.n292 3.n291 0.006
R3969 3.n294 3.n293 0.006
R3970 3.n210 3.n205 0.005
R3971 3.n189 3.n188 0.005
R3972 3.n188 3.n187 0.005
R3973 3.n155 3.n154 0.005
R3974 3.n68 3.n67 0.005
R3975 3.n39 3.n38 0.005
R3976 3.n47 3.n39 0.005
R3977 3.n45 3.n44 0.005
R3978 3.n28 3.n18 0.005
R3979 3.n217 3.n211 0.005
R3980 3.n194 3.n190 0.005
R3981 3.n123 3.n122 0.005
R3982 3.n49 3.n48 0.005
R3983 3.n36 3.n35 0.005
R3984 3.n30 3.n29 0.005
R3985 3.n178 3.n177 0.005
R3986 3.n153 3.n152 0.005
R3987 3.n78 3.n77 0.005
R3988 3.n52 3.n51 0.005
R3989 3.n227 3.n222 0.004
R3990 3.n6 3.n5 0.004
R3991 3.n271 3.n270 0.003
R3992 3.n324 3.n321 0.003
R3993 3.n337 3.n336 0.003
R3994 3.n303 3.n302 0.003
R3995 3.n199 3.n198 0.003
R3996 3.n202 3.n201 0.003
R3997 3.n161 3.n160 0.003
R3998 3.n146 3.n139 0.003
R3999 3.n131 3.n130 0.003
R4000 3.n230 3.n229 0.003
R4001 3.n213 3.n212 0.003
R4002 3.n193 3.n192 0.003
R4003 3.n150 3.n149 0.003
R4004 3.n148 3.n147 0.003
R4005 3.n132 3.n124 0.003
R4006 3.n235 3.n234 0.003
R4007 3.n218 3.n197 0.003
R4008 3.n135 3.n134 0.003
R4009 3.n110 3.n85 0.003
R4010 3.n32 3.n31 0.003
R4011 3.n258 3.n257 0.001
R4012 3.n244 3.n243 0.001
R4013 3.n241 3.n240 0.001
R4014 3.n166 3.n165 0.001
R4015 3.n115 3.n114 0.001
R4016 3.n90 3.n89 0.001
R4017 3.n102 3.n101 0.001
R4018 3.n99 3.n98 0.001
R4019 3.n64 3.n63 0.001
R4020 3.n26 3.n25 0.001
R4021 3.n133 3.n119 0.001
R4022 3.n109 3.n108 0.001
R4023 3.n87 3.n86 0.001
R4024 3.n82 3.n79 0.001
R4025 3.n55 3.n54 0.001
R4026 3.n15 3.n14 0.001
R4027 finb.n67 finb.t5 733.434
R4028 finb.n137 finb.t2 733.434
R4029 finb.n29 finb.t3 396.757
R4030 finb.n105 finb.t4 396.757
R4031 finb.n392 finb.n391 92.5
R4032 finb.n455 finb.n454 92.5
R4033 finb.n391 finb.t0 70.344
R4034 finb.n405 finb.n404 31.034
R4035 finb.n472 finb.n471 31.034
R4036 finb.n415 finb.n414 9.3
R4037 finb.n481 finb.n480 9.3
R4038 finb.n473 finb.n472 9.3
R4039 finb.n406 finb.n405 9.3
R4040 finb.n202 finb.n201 9.3
R4041 finb.n304 finb.n303 9.3
R4042 finb.n268 finb.n267 9.154
R4043 finb.n393 finb.n392 8.282
R4044 finb.n456 finb.n455 8.282
R4045 finb.n267 finb.t1 7.141
R4046 finb.n362 finb.n361 7.03
R4047 finb.n145 finb.n144 7.03
R4048 finb.n493 finb.n376 6.38
R4049 finb.n406 finb.n402 5.647
R4050 finb.n473 finb.n469 5.647
R4051 finb.n453 finb.n452 4.65
R4052 finb.n269 finb.n268 4.65
R4053 finb.n457 finb.n456 4.5
R4054 finb.n464 finb.n463 4.5
R4055 finb.n398 finb.n393 4.5
R4056 finb.n475 finb.n474 4.5
R4057 finb.n451 finb.n450 4.5
R4058 finb.n409 finb.n408 4.5
R4059 finb.n487 finb.n485 4.5
R4060 finb.n420 finb.n419 4.5
R4061 finb.n168 finb.n162 4.5
R4062 finb.n307 finb.n299 4.5
R4063 finb.n329 finb.n323 4.5
R4064 finb.n286 finb.n285 4.5
R4065 finb.n256 finb.n253 4.5
R4066 finb.n271 finb.n265 4.5
R4067 finb.n245 finb.n233 4.5
R4068 finb.n261 finb.n260 4.5
R4069 finb.n242 finb.n237 4.5
R4070 finb.n213 finb.n212 4.5
R4071 finb.n187 finb.n183 4.5
R4072 finb.n350 finb.n349 4.5
R4073 finb.n323 finb.n320 4.141
R4074 finb.n183 finb.n182 4.141
R4075 finb.n404 finb.n403 4.137
R4076 finb.n471 finb.n470 4.137
R4077 finb.n419 finb.n417 3.764
R4078 finb.n474 finb.n467 3.764
R4079 finb.n299 finb.n296 3.764
R4080 finb.n237 finb.n235 3.764
R4081 finb.n408 finb.n407 3.388
R4082 finb.n485 finb.n484 3.388
R4083 finb.n349 finb.n346 3.388
R4084 finb.n285 finb.n284 3.388
R4085 finb.n212 finb.n211 3.388
R4086 finb.n162 finb.n161 3.388
R4087 finb.n408 finb.n406 3.011
R4088 finb.n393 finb.n390 3.011
R4089 finb.n485 finb.n483 3.011
R4090 finb.n349 finb.n348 3.011
R4091 finb.n285 finb.n282 3.011
R4092 finb.n253 finb.n251 3.011
R4093 finb.n201 finb.n200 3.011
R4094 finb.n212 finb.n210 3.011
R4095 finb.n162 finb.n160 3.011
R4096 finb.n419 finb.n418 2.635
R4097 finb.n463 finb.n462 2.635
R4098 finb.n474 finb.n473 2.635
R4099 finb.n299 finb.n298 2.635
R4100 finb.n303 finb.n302 2.635
R4101 finb.n233 finb.n232 2.635
R4102 finb.n237 finb.n236 2.635
R4103 finb.n493 finb.n492 2.632
R4104 finb.n323 finb.n322 2.258
R4105 finb.n183 finb.n181 2.258
R4106 finb.n233 finb.n231 1.505
R4107 finb.n488 finb.n487 1.5
R4108 finb.n421 finb.n420 1.5
R4109 finb.n148 finb.n146 1.5
R4110 finb.n169 finb.n168 1.5
R4111 finb.n330 finb.n329 1.5
R4112 finb.n368 finb.n367 1.5
R4113 finb.n308 finb.n307 1.5
R4114 finb.n287 finb.n286 1.5
R4115 finb.n257 finb.n256 1.5
R4116 finb.n272 finb.n271 1.5
R4117 finb.n246 finb.n245 1.5
R4118 finb.n262 finb.n261 1.5
R4119 finb.n214 finb.n213 1.5
R4120 finb.n188 finb.n187 1.5
R4121 finb.n351 finb.n350 1.5
R4122 finb.n22 finb.n21 1.435
R4123 finb.n55 finb.n54 1.435
R4124 finb.n121 finb.n120 1.435
R4125 finb.n500 finb.n499 1.435
R4126 finb.n31 finb.n29 1.354
R4127 finb.n68 finb.n67 1.354
R4128 finb.n107 finb.n105 1.354
R4129 finb.n138 finb.n137 1.354
R4130 finb.n108 finb.n107 1.142
R4131 finb.n23 finb.n22 1.142
R4132 finb.n56 finb.n55 1.142
R4133 finb.n139 finb.n138 1.142
R4134 finb.n69 finb.n68 1.14
R4135 finb.n24 finb.n23 1.138
R4136 finb.n509 finb.n139 1.138
R4137 finb.n57 finb.n56 1.138
R4138 finb.n109 finb.n108 1.138
R4139 finb.n8 finb.n7 1.137
R4140 finb.n37 finb.n36 1.137
R4141 finb.n4 finb.n3 1.137
R4142 finb.n14 finb.n13 1.137
R4143 finb.n32 finb.n31 1.137
R4144 finb.n80 finb.n79 1.137
R4145 finb.n47 finb.n46 1.137
R4146 finb.n61 finb.n60 1.137
R4147 finb.n74 finb.n73 1.137
R4148 finb.n122 finb.n121 1.137
R4149 finb.n92 finb.n91 1.137
R4150 finb.n114 finb.n113 1.137
R4151 finb.n89 finb.n88 1.137
R4152 finb.n98 finb.n97 1.137
R4153 finb.n150 finb.n149 1.137
R4154 finb.n171 finb.n170 1.137
R4155 finb.n190 finb.n189 1.137
R4156 finb.n198 finb.n197 1.137
R4157 finb.n216 finb.n215 1.137
R4158 finb.n223 finb.n222 1.137
R4159 finb.n316 finb.n315 1.137
R4160 finb.n374 finb.n373 1.137
R4161 finb.n335 finb.n334 1.137
R4162 finb.n291 finb.n290 1.137
R4163 finb.n312 finb.n311 1.137
R4164 finb.n274 finb.n273 1.137
R4165 finb.n250 finb.n249 1.137
R4166 finb.n358 finb.n357 1.137
R4167 finb.n518 finb.n517 1.137
R4168 finb.n505 finb.n504 1.137
R4169 finb.n513 finb.n512 1.137
R4170 finb.n129 finb.n128 1.137
R4171 finb.n501 finb.n500 1.137
R4172 finb.n94 finb.n93 1.136
R4173 finb.n508 finb.n507 1.136
R4174 finb.n520 finb.n519 1.136
R4175 finb.n124 finb.n123 1.136
R4176 finb.n82 finb.n81 1.136
R4177 finb.n40 finb.n39 1.136
R4178 finb.n10 finb.n9 1.136
R4179 finb.n253 finb.n252 1.129
R4180 finb.n491 finb.n490 0.853
R4181 finb.n402 finb.n401 0.752
R4182 finb.n469 finb.n468 0.752
R4183 finb.n423 finb.n422 0.704
R4184 finb.n361 finb.n360 0.155
R4185 finb.n144 finb.n143 0.155
R4186 finb.n348 finb.n347 0.144
R4187 finb.n160 finb.n159 0.144
R4188 finb.n322 finb.n321 0.133
R4189 finb.n181 finb.n180 0.132
R4190 finb.n84 finb.n83 0.106
R4191 finb.n42 finb.n41 0.099
R4192 finb.n29 finb.n28 0.083
R4193 finb.n67 finb.n66 0.083
R4194 finb.n105 finb.n104 0.083
R4195 finb.n137 finb.n136 0.083
R4196 finb.n494 finb.n493 0.061
R4197 finb finb.n125 0.058
R4198 finb.n374 finb.n358 0.049
R4199 finb.n274 finb.n250 0.049
R4200 finb.n171 finb.n150 0.049
R4201 finb.n343 finb.n342 0.047
R4202 finb.n289 finb.n288 0.045
R4203 finb.n273 finb.n272 0.045
R4204 finb.n304 finb.n301 0.043
R4205 finb.n188 finb.n176 0.043
R4206 finb.n169 finb.n155 0.041
R4207 finb finb.n521 0.041
R4208 finb.n245 finb.n230 0.039
R4209 finb.n373 finb.n372 0.039
R4210 finb.n256 finb.n255 0.037
R4211 finb.n149 finb.n140 0.037
R4212 finb.n395 finb.n394 0.035
R4213 finb.n459 finb.n458 0.035
R4214 finb.n378 finb.n377 0.035
R4215 finb.n440 finb.n439 0.035
R4216 finb.n326 finb.n325 0.035
R4217 finb.n240 finb.n239 0.035
R4218 finb.n388 finb.n387 0.034
R4219 finb.n449 finb.n448 0.034
R4220 finb.n165 finb.n164 0.034
R4221 finb.n371 finb.n370 0.034
R4222 finb.n264 finb.n263 0.034
R4223 finb.n154 finb.n153 0.034
R4224 finb.n478 finb.n477 0.032
R4225 finb.n447 finb.n446 0.032
R4226 finb.n3 finb.n2 0.032
R4227 finb.n79 finb.n76 0.032
R4228 finb.n88 finb.n87 0.032
R4229 finb.n368 finb.n359 0.032
R4230 finb.n247 finb.n246 0.032
R4231 finb.n228 finb.n227 0.032
R4232 finb.n517 finb.n515 0.032
R4233 finb.n424 finb.n423 0.031
R4234 finb.n435 finb.n434 0.031
R4235 finb.n336 finb.n335 0.031
R4236 finb.n291 finb.n276 0.031
R4237 finb.n224 finb.n223 0.031
R4238 finb.n190 finb.n173 0.031
R4239 finb.n412 finb.n411 0.03
R4240 finb.n481 finb.n479 0.03
R4241 finb.n386 finb.n385 0.03
R4242 finb.n445 finb.n444 0.03
R4243 finb.n365 finb.n364 0.03
R4244 finb.n354 finb.n353 0.03
R4245 finb.n287 finb.n277 0.03
R4246 finb.n258 finb.n257 0.03
R4247 finb.n415 finb.n413 0.028
R4248 finb.n397 finb.n396 0.028
R4249 finb.n461 finb.n460 0.028
R4250 finb.n383 finb.n382 0.028
R4251 finb.n380 finb.n379 0.028
R4252 finb.n442 finb.n441 0.028
R4253 finb.n488 finb.n449 0.028
R4254 finb.n28 finb.n27 0.028
R4255 finb.n26 finb.n25 0.028
R4256 finb.n19 finb.n18 0.028
R4257 finb.n21 finb.n20 0.028
R4258 finb.n36 finb.n35 0.028
R4259 finb.n3 finb.n1 0.028
R4260 finb.n7 finb.n6 0.028
R4261 finb.n13 finb.n11 0.028
R4262 finb.n54 finb.n53 0.028
R4263 finb.n52 finb.n51 0.028
R4264 finb.n64 finb.n63 0.028
R4265 finb.n66 finb.n65 0.028
R4266 finb.n46 finb.n45 0.028
R4267 finb.n60 finb.n59 0.028
R4268 finb.n79 finb.n78 0.028
R4269 finb.n104 finb.n103 0.028
R4270 finb.n102 finb.n101 0.028
R4271 finb.n118 finb.n117 0.028
R4272 finb.n120 finb.n119 0.028
R4273 finb.n97 finb.n96 0.028
R4274 finb.n88 finb.n86 0.028
R4275 finb.n91 finb.n90 0.028
R4276 finb.n113 finb.n111 0.028
R4277 finb.n175 finb.n174 0.028
R4278 finb.n499 finb.n498 0.028
R4279 finb.n497 finb.n496 0.028
R4280 finb.n134 finb.n133 0.028
R4281 finb.n136 finb.n135 0.028
R4282 finb.n504 finb.n503 0.028
R4283 finb.n512 finb.n511 0.028
R4284 finb.n517 finb.n516 0.028
R4285 finb.n128 finb.n126 0.028
R4286 finb.n422 finb.n421 0.027
R4287 finb.n428 finb.n427 0.027
R4288 finb.n431 finb.n430 0.027
R4289 finb.n316 finb.n312 0.027
R4290 finb.n216 finb.n198 0.027
R4291 finb.n421 finb.n388 0.026
R4292 finb.n344 finb.n343 0.026
R4293 finb.n207 finb.n206 0.026
R4294 finb.n356 finb.n355 0.026
R4295 finb.n157 finb.n156 0.024
R4296 finb.n167 finb.n166 0.024
R4297 finb.n334 finb.n333 0.024
R4298 finb.n314 finb.n313 0.024
R4299 finb.n311 finb.n310 0.024
R4300 finb.n222 finb.n221 0.024
R4301 finb.n197 finb.n196 0.024
R4302 finb.n152 finb.n151 0.024
R4303 finb.n298 finb.n297 0.024
R4304 finb.n210 finb.n209 0.024
R4305 finb.n457 finb.n453 0.022
R4306 finb.n438 finb.n437 0.022
R4307 finb.n490 finb.n488 0.022
R4308 finb.n340 finb.n339 0.022
R4309 finb.n327 finb.n326 0.022
R4310 finb.n186 finb.n185 0.022
R4311 finb.n214 finb.n199 0.022
R4312 finb.n453 finb.n451 0.02
R4313 finb.n437 finb.n436 0.02
R4314 finb.n329 finb.n319 0.02
R4315 finb.n178 finb.n177 0.02
R4316 finb.n187 finb.n186 0.02
R4317 finb.n491 finb.n435 0.019
R4318 finb.n492 finb.n491 0.019
R4319 finb.n420 finb.n389 0.018
R4320 finb.n416 finb.n415 0.018
R4321 finb.n413 finb.n412 0.018
R4322 finb.n475 finb.n466 0.018
R4323 finb.n387 finb.n386 0.018
R4324 finb.n307 finb.n295 0.018
R4325 finb.n305 finb.n304 0.018
R4326 finb.n243 finb.n242 0.018
R4327 finb.n148 finb.n147 0.017
R4328 finb.n409 finb.n400 0.017
R4329 finb.n479 finb.n478 0.017
R4330 finb.n482 finb.n481 0.017
R4331 finb.n487 finb.n486 0.017
R4332 finb.n385 finb.n384 0.017
R4333 finb.n446 finb.n445 0.017
R4334 finb.n448 finb.n447 0.017
R4335 finb.n31 finb.n30 0.017
R4336 finb.n36 finb.n34 0.017
R4337 finb.n13 finb.n12 0.017
R4338 finb.n22 finb.n17 0.017
R4339 finb.n55 finb.n50 0.017
R4340 finb.n46 finb.n44 0.017
R4341 finb.n73 finb.n72 0.017
R4342 finb.n68 finb.n62 0.017
R4343 finb.n107 finb.n106 0.017
R4344 finb.n97 finb.n95 0.017
R4345 finb.n113 finb.n112 0.017
R4346 finb.n121 finb.n116 0.017
R4347 finb.n350 finb.n340 0.017
R4348 finb.n286 finb.n281 0.017
R4349 finb.n270 finb.n269 0.017
R4350 finb.n269 finb.n266 0.017
R4351 finb.n203 finb.n202 0.017
R4352 finb.n213 finb.n208 0.017
R4353 finb.n168 finb.n167 0.017
R4354 finb.n355 finb.n354 0.017
R4355 finb.n500 finb.n495 0.017
R4356 finb.n504 finb.n502 0.017
R4357 finb.n128 finb.n127 0.017
R4358 finb.n138 finb.n132 0.017
R4359 finb.n8 finb.n5 0.016
R4360 finb.n61 finb.n58 0.016
R4361 finb.n80 finb.n75 0.016
R4362 finb.n89 finb.n85 0.016
R4363 finb.n513 finb.n510 0.016
R4364 finb.n518 finb.n514 0.016
R4365 finb.n376 finb.n375 0.016
R4366 finb.n337 finb.n336 0.016
R4367 finb.n276 finb.n275 0.016
R4368 finb.n225 finb.n224 0.016
R4369 finb.n173 finb.n172 0.016
R4370 finb.n410 finb.n409 0.015
R4371 finb.n399 finb.n398 0.015
R4372 finb.n487 finb.n482 0.015
R4373 finb.n382 finb.n381 0.015
R4374 finb.n27 finb.n26 0.015
R4375 finb.n20 finb.n19 0.015
R4376 finb.n53 finb.n52 0.015
R4377 finb.n65 finb.n64 0.015
R4378 finb.n78 finb.n77 0.015
R4379 finb.n103 finb.n102 0.015
R4380 finb.n119 finb.n118 0.015
R4381 finb.n310 finb.n309 0.015
R4382 finb.n221 finb.n220 0.015
R4383 finb.n498 finb.n497 0.015
R4384 finb.n135 finb.n134 0.015
R4385 finb.n420 finb.n416 0.013
R4386 finb.n465 finb.n464 0.013
R4387 finb.n476 finb.n475 0.013
R4388 finb.n444 finb.n443 0.013
R4389 finb.n245 finb.n244 0.013
R4390 finb.n213 finb.n204 0.013
R4391 finb.n215 finb.n214 0.013
R4392 finb.n196 finb.n195 0.013
R4393 finb.n284 finb.n283 0.012
R4394 finb.n235 finb.n234 0.012
R4395 finb.n429 finb.n428 0.012
R4396 finb.n430 finb.n429 0.012
R4397 finb.n9 finb.n4 0.012
R4398 finb.n9 finb.n8 0.012
R4399 finb.n81 finb.n61 0.012
R4400 finb.n81 finb.n80 0.012
R4401 finb.n93 finb.n89 0.012
R4402 finb.n93 finb.n92 0.012
R4403 finb.n519 finb.n513 0.012
R4404 finb.n519 finb.n518 0.012
R4405 finb.n490 finb.n489 0.012
R4406 finb.n400 finb.n399 0.011
R4407 finb.n466 finb.n465 0.011
R4408 finb.n426 finb.n425 0.011
R4409 finb.n433 finb.n432 0.011
R4410 finb.n39 finb.n38 0.011
R4411 finb.n16 finb.n15 0.011
R4412 finb.n49 finb.n48 0.011
R4413 finb.n71 finb.n70 0.011
R4414 finb.n100 finb.n99 0.011
R4415 finb.n123 finb.n115 0.011
R4416 finb.n325 finb.n324 0.011
R4417 finb.n307 finb.n306 0.011
R4418 finb.n279 finb.n278 0.011
R4419 finb.n281 finb.n280 0.011
R4420 finb.n244 finb.n243 0.011
R4421 finb.n241 finb.n240 0.011
R4422 finb.n164 finb.n163 0.011
R4423 finb.n332 finb.n331 0.011
R4424 finb.n315 finb.n314 0.011
R4425 finb.n311 finb.n308 0.011
R4426 finb.n246 finb.n228 0.011
R4427 finb.n507 finb.n506 0.011
R4428 finb.n131 finb.n130 0.011
R4429 finb.n37 finb.n33 0.01
R4430 finb.n75 finb.n74 0.01
R4431 finb.n114 finb.n110 0.01
R4432 finb.n458 finb.n457 0.009
R4433 finb.n439 finb.n438 0.009
R4434 finb.n367 finb.n366 0.009
R4435 finb.n366 finb.n365 0.009
R4436 finb.n364 finb.n363 0.009
R4437 finb.n345 finb.n344 0.009
R4438 finb.n206 finb.n205 0.009
R4439 finb.n158 finb.n157 0.009
R4440 finb.n142 finb.n141 0.009
R4441 finb.n146 finb.n142 0.009
R4442 finb.n373 finb.n368 0.009
R4443 finb.n372 finb.n371 0.009
R4444 finb.n357 finb.n356 0.009
R4445 finb.n197 finb.n193 0.009
R4446 finb.n170 finb.n152 0.009
R4447 finb.n149 finb.n148 0.009
R4448 finb.n335 finb.n318 0.009
R4449 finb.n317 finb.n316 0.009
R4450 finb.n312 finb.n293 0.009
R4451 finb.n292 finb.n291 0.009
R4452 finb.n223 finb.n218 0.009
R4453 finb.n217 finb.n216 0.009
R4454 finb.n198 finb.n192 0.009
R4455 finb.n191 finb.n190 0.009
R4456 finb.n396 finb.n395 0.007
R4457 finb.n460 finb.n459 0.007
R4458 finb.n379 finb.n378 0.007
R4459 finb.n441 finb.n440 0.007
R4460 finb.n259 finb.n258 0.007
R4461 finb.n248 finb.n247 0.007
R4462 finb.n425 finb.n424 0.006
R4463 finb.n427 finb.n426 0.006
R4464 finb.n432 finb.n431 0.006
R4465 finb.n434 finb.n433 0.006
R4466 finb.n39 finb.n32 0.006
R4467 finb.n38 finb.n37 0.006
R4468 finb.n15 finb.n14 0.006
R4469 finb.n48 finb.n47 0.006
R4470 finb.n74 finb.n71 0.006
R4471 finb.n99 finb.n98 0.006
R4472 finb.n115 finb.n114 0.006
R4473 finb.n123 finb.n122 0.006
R4474 finb.n507 finb.n501 0.006
R4475 finb.n506 finb.n505 0.006
R4476 finb.n130 finb.n129 0.006
R4477 finb.n350 finb.n345 0.005
R4478 finb.n329 finb.n328 0.005
R4479 finb.n328 finb.n327 0.005
R4480 finb.n295 finb.n294 0.005
R4481 finb.n208 finb.n207 0.005
R4482 finb.n179 finb.n178 0.005
R4483 finb.n187 finb.n179 0.005
R4484 finb.n185 finb.n184 0.005
R4485 finb.n168 finb.n158 0.005
R4486 finb.n357 finb.n351 0.005
R4487 finb.n334 finb.n330 0.005
R4488 finb.n263 finb.n262 0.005
R4489 finb.n189 finb.n188 0.005
R4490 finb.n176 finb.n175 0.005
R4491 finb.n170 finb.n169 0.005
R4492 finb.n318 finb.n317 0.005
R4493 finb.n293 finb.n292 0.005
R4494 finb.n218 finb.n217 0.005
R4495 finb.n192 finb.n191 0.005
R4496 finb.n367 finb.n362 0.004
R4497 finb.n146 finb.n145 0.004
R4498 finb.n94 finb.n84 0.004
R4499 finb.n70 finb.n69 0.003
R4500 finb.n10 finb.n0 0.003
R4501 finb.n41 finb.n40 0.003
R4502 finb.n83 finb.n82 0.003
R4503 finb.n125 finb.n124 0.003
R4504 finb.n521 finb.n520 0.003
R4505 finb.n508 finb.n494 0.003
R4506 finb.n411 finb.n410 0.003
R4507 finb.n464 finb.n461 0.003
R4508 finb.n477 finb.n476 0.003
R4509 finb.n443 finb.n442 0.003
R4510 finb.n339 finb.n338 0.003
R4511 finb.n342 finb.n341 0.003
R4512 finb.n301 finb.n300 0.003
R4513 finb.n286 finb.n279 0.003
R4514 finb.n271 finb.n270 0.003
R4515 finb.n370 finb.n369 0.003
R4516 finb.n353 finb.n352 0.003
R4517 finb.n333 finb.n332 0.003
R4518 finb.n290 finb.n289 0.003
R4519 finb.n288 finb.n287 0.003
R4520 finb.n272 finb.n264 0.003
R4521 finb.n375 finb.n374 0.003
R4522 finb.n358 finb.n337 0.003
R4523 finb.n275 finb.n274 0.003
R4524 finb.n250 finb.n225 0.003
R4525 finb.n172 finb.n171 0.003
R4526 finb.n56 finb.n49 0.003
R4527 finb.n108 finb.n100 0.003
R4528 finb.n139 finb.n131 0.003
R4529 finb.n23 finb.n16 0.003
R4530 finb.n43 finb.n42 0.002
R4531 finb.n57 finb.n43 0.002
R4532 finb.n109 finb.n94 0.002
R4533 finb.n509 finb.n508 0.002
R4534 finb.n124 finb.n109 0.002
R4535 finb.n520 finb.n509 0.002
R4536 finb.n82 finb.n57 0.002
R4537 finb.n40 finb.n24 0.002
R4538 finb.n24 finb.n10 0.002
R4539 finb.n398 finb.n397 0.001
R4540 finb.n384 finb.n383 0.001
R4541 finb.n381 finb.n380 0.001
R4542 finb.n306 finb.n305 0.001
R4543 finb.n255 finb.n254 0.001
R4544 finb.n230 finb.n229 0.001
R4545 finb.n242 finb.n241 0.001
R4546 finb.n239 finb.n238 0.001
R4547 finb.n204 finb.n203 0.001
R4548 finb.n166 finb.n165 0.001
R4549 finb.n273 finb.n259 0.001
R4550 finb.n249 finb.n248 0.001
R4551 finb.n227 finb.n226 0.001
R4552 finb.n222 finb.n219 0.001
R4553 finb.n195 finb.n194 0.001
R4554 finb.n155 finb.n154 0.001
R4555 net1.n3 net1.n2 13.361
R4556 net1.n88 net1.n87 13.361
R4557 net1.n13 net1.n11 9.3
R4558 net1.n7 net1.n5 9.3
R4559 net1.n18 net1.n15 9.3
R4560 net1.n134 net1.n126 9.3
R4561 net1.n134 net1.n133 9.3
R4562 net1.n24 net1.n22 9.3
R4563 net1.n35 net1.n33 9.3
R4564 net1.n32 net1.n30 9.3
R4565 net1.n43 net1.n41 9.3
R4566 net1.n43 net1.n42 9.3
R4567 net1.n54 net1.n52 9.3
R4568 net1.n54 net1.n53 9.3
R4569 net1.n65 net1.n63 9.3
R4570 net1.n65 net1.n64 9.3
R4571 net1.n76 net1.n74 9.3
R4572 net1.n76 net1.n75 9.3
R4573 net1.n100 net1.n98 9.3
R4574 net1.n100 net1.n99 9.3
R4575 net1.n168 net1.n106 9.3
R4576 net1.n168 net1.n167 9.3
R4577 net1.n160 net1.n111 9.3
R4578 net1.n160 net1.n159 9.3
R4579 net1.n153 net1.n115 9.3
R4580 net1.n153 net1.n152 9.3
R4581 net1.n146 net1.n119 9.3
R4582 net1.n146 net1.n145 9.3
R4583 net1.n29 net1.n26 9.3
R4584 net1.n35 net1.n34 9.3
R4585 net1.n40 net1.n37 9.3
R4586 net1.n46 net1.n44 9.3
R4587 net1.n51 net1.n48 9.3
R4588 net1.n57 net1.n55 9.3
R4589 net1.n62 net1.n59 9.3
R4590 net1.n68 net1.n66 9.3
R4591 net1.n73 net1.n70 9.3
R4592 net1.n79 net1.n77 9.3
R4593 net1.n84 net1.n81 9.3
R4594 net1.n94 net1.n91 9.3
R4595 net1.n97 net1.n95 9.3
R4596 net1.n105 net1.n102 9.3
R4597 net1 net1.n1 9.3
R4598 net1.n166 net1.n109 9.3
R4599 net1.n162 net1.n110 9.3
R4600 net1.n158 net1.n113 9.3
R4601 net1.n155 net1.n114 9.3
R4602 net1.n151 net1.n117 9.3
R4603 net1.n148 net1.n118 9.3
R4604 net1.n144 net1.n121 9.3
R4605 net1.n141 net1.n122 9.3
R4606 net1.n137 net1.n125 9.3
R4607 net1.n139 net1.n123 9.3
R4608 net1.n40 net1.n39 9.3
R4609 net1.n46 net1.n45 9.3
R4610 net1.n51 net1.n50 9.3
R4611 net1.n57 net1.n56 9.3
R4612 net1.n62 net1.n61 9.3
R4613 net1.n68 net1.n67 9.3
R4614 net1.n73 net1.n72 9.3
R4615 net1.n79 net1.n78 9.3
R4616 net1.n84 net1.n83 9.3
R4617 net1.n94 net1.n93 9.3
R4618 net1.n97 net1.n96 9.3
R4619 net1.n105 net1.n104 9.3
R4620 net1 net1.n0 9.3
R4621 net1.n166 net1.n165 9.3
R4622 net1.n162 net1.n161 9.3
R4623 net1.n158 net1.n157 9.3
R4624 net1.n155 net1.n154 9.3
R4625 net1.n151 net1.n150 9.3
R4626 net1.n148 net1.n147 9.3
R4627 net1.n144 net1.n143 9.3
R4628 net1.n141 net1.n140 9.3
R4629 net1.n137 net1.n136 9.3
R4630 net1.n139 net1.n138 9.3
R4631 net1.n32 net1.n31 9.3
R4632 net1.n29 net1.n28 9.3
R4633 net1.n24 net1.n23 9.3
R4634 net1.n21 net1.n19 9.3
R4635 net1.n21 net1.n20 9.3
R4636 net1.n18 net1.n17 9.3
R4637 net1.n130 net1.n128 9.3
R4638 net1.n132 net1.n127 9.3
R4639 net1.n132 net1.n131 9.3
R4640 net1.n130 net1.n129 9.3
R4641 net1.n13 net1.n12 9.3
R4642 net1.n10 net1.n8 9.3
R4643 net1.n10 net1.n9 9.3
R4644 net1.n7 net1.n6 9.3
R4645 net1.n164 net1.n163 8.016
R4646 net1.n108 net1.n107 8.016
R4647 net1.n86 net1.n4 4.558
R4648 net1.n89 net1.n3 4.558
R4649 net1.n86 net1.n85 4.558
R4650 net1.n89 net1.n88 4.558
R4651 net1.n163 net1.t0 2.9
R4652 net1.n107 net1.t1 2.9
R4653 net1.n81 net1.n80 0.536
R4654 net1.n91 net1.n90 0.536
R4655 net1.n83 net1.n82 0.536
R4656 net1.n93 net1.n92 0.536
R4657 net1.n72 net1.n71 0.506
R4658 net1.n104 net1.n103 0.506
R4659 net1.n70 net1.n69 0.506
R4660 net1.n102 net1.n101 0.506
R4661 net1.n59 net1.n58 0.475
R4662 net1.n109 net1.n108 0.475
R4663 net1.n61 net1.n60 0.475
R4664 net1.n165 net1.n164 0.475
R4665 net1.n157 net1.n156 0.445
R4666 net1.n48 net1.n47 0.445
R4667 net1.n113 net1.n112 0.445
R4668 net1.n50 net1.n49 0.445
R4669 net1.n37 net1.n36 0.413
R4670 net1.n117 net1.n116 0.413
R4671 net1.n39 net1.n38 0.413
R4672 net1.n150 net1.n149 0.413
R4673 net1.n28 net1.n27 0.382
R4674 net1.n143 net1.n142 0.382
R4675 net1.n121 net1.n120 0.382
R4676 net1.n26 net1.n25 0.382
R4677 net1.n15 net1.n14 0.349
R4678 net1.n17 net1.n16 0.349
R4679 net1.n125 net1.n124 0.349
R4680 net1.n136 net1.n135 0.349
R4681 net1.n89 net1.n86 0.039
R4682 net1.n18 net1.n13 0.03
R4683 net1.n29 net1.n24 0.03
R4684 net1.n40 net1.n35 0.03
R4685 net1.n51 net1.n46 0.03
R4686 net1.n62 net1.n57 0.03
R4687 net1.n73 net1.n68 0.03
R4688 net1.n84 net1.n79 0.03
R4689 net1.n97 net1.n94 0.03
R4690 net1 net1.n105 0.03
R4691 net1.n166 net1.n162 0.03
R4692 net1.n158 net1.n155 0.03
R4693 net1.n151 net1.n148 0.03
R4694 net1.n144 net1.n141 0.03
R4695 net1.n137 net1.n134 0.03
R4696 net1.n86 net1.n84 0.009
R4697 net1.n94 net1.n89 0.009
R4698 net1.n13 net1.n10 0.008
R4699 net1.n134 net1.n132 0.008
R4700 net1.n24 net1.n21 0.007
R4701 net1.n76 net1.n73 0.007
R4702 net1.n105 net1.n100 0.007
R4703 net1.n141 net1.n139 0.007
R4704 net1.n35 net1.n32 0.006
R4705 net1.n65 net1.n62 0.006
R4706 net1.n168 net1.n166 0.006
R4707 net1.n148 net1.n146 0.006
R4708 net1.n46 net1.n43 0.005
R4709 net1.n54 net1.n51 0.005
R4710 net1.n160 net1.n158 0.005
R4711 net1.n155 net1.n153 0.005
R4712 net1.n43 net1.n40 0.004
R4713 net1.n153 net1.n151 0.004
R4714 net1.n32 net1.n29 0.003
R4715 net1.n57 net1.n54 0.003
R4716 net1.n162 net1.n160 0.003
R4717 net1.n146 net1.n144 0.003
R4718 net1.n21 net1.n18 0.002
R4719 net1.n68 net1.n65 0.002
R4720 net1 net1.n168 0.002
R4721 net1.n139 net1.n137 0.002
R4722 net1.n10 net1.n7 0.001
R4723 net1.n79 net1.n76 0.001
R4724 net1.n100 net1.n97 0.001
R4725 net1.n132 net1.n130 0.001
R4726 fin fin.t6 1038.56
R4727 fin.n121 fin.t2 795.567
R4728 fin.n80 fin.t5 731.671
R4729 fin.n51 fin.t3 731.671
R4730 fin.n14 fin.t7 730.672
R4731 fin.n100 fin.t1 400.617
R4732 fin.n57 fin.t4 400.616
R4733 fin.n14 fin.t0 395.84
R4734 fin.n89 fin.n87 1.435
R4735 fin.n22 fin.n21 1.435
R4736 fin.n130 fin.n120 1.354
R4737 fin.n81 fin.n80 1.354
R4738 fin.n52 fin.n51 1.354
R4739 fin.n82 fin.n81 1.142
R4740 fin.n23 fin.n22 1.14
R4741 fin.n83 fin.n82 1.138
R4742 fin.n90 fin.n89 1.137
R4743 fin.n66 fin.n65 1.137
R4744 fin.n72 fin.n71 1.137
R4745 fin.n61 fin.n60 1.137
R4746 fin.n95 fin.n94 1.137
R4747 fin.n28 fin.n27 1.137
R4748 fin.n33 fin.n32 1.137
R4749 fin.n53 fin.n52 1.137
R4750 fin.n43 fin.n42 1.137
R4751 fin.n37 fin.n36 1.137
R4752 fin.n120 fin.n119 1.137
R4753 fin.n68 fin.n67 1.136
R4754 fin.n118 fin.n106 1.136
R4755 fin.n55 fin.n54 1.136
R4756 fin.n98 fin.n97 1.136
R4757 fin fin.n130 0.392
R4758 fin.n102 fin.n101 0.154
R4759 fin.n57 fin.n56 0.123
R4760 fin.n100 fin.n99 0.123
R4761 fin.n58 fin.n57 0.091
R4762 fin.n80 fin.n79 0.083
R4763 fin.n51 fin.n50 0.083
R4764 fin.n130 fin.n129 0.076
R4765 fin.n122 fin.n121 0.076
R4766 fin.n101 fin.n100 0.072
R4767 fin.n47 fin.n46 0.064
R4768 fin.n126 fin.n125 0.059
R4769 fin.n65 fin.n63 0.032
R4770 fin.n36 fin.n35 0.032
R4771 fin.n8 fin.n7 0.032
R4772 fin.n7 fin.n6 0.032
R4773 fin.n13 fin.n12 0.03
R4774 fin.n2 fin.n1 0.03
R4775 fin.n87 fin.n86 0.028
R4776 fin.n85 fin.n84 0.028
R4777 fin.n77 fin.n76 0.028
R4778 fin.n79 fin.n78 0.028
R4779 fin.n94 fin.n93 0.028
R4780 fin.n60 fin.n59 0.028
R4781 fin.n65 fin.n64 0.028
R4782 fin.n71 fin.n69 0.028
R4783 fin.n21 fin.n20 0.028
R4784 fin.n48 fin.n47 0.028
R4785 fin.n50 fin.n49 0.028
R4786 fin.n32 fin.n31 0.028
R4787 fin.n42 fin.n40 0.028
R4788 fin.n11 fin.n10 0.028
R4789 fin.n9 fin.n8 0.028
R4790 fin.n6 fin.n5 0.028
R4791 fin.n4 fin.n3 0.028
R4792 fin.n129 fin.n128 0.026
R4793 fin.n127 fin.n126 0.026
R4794 fin.n125 fin.n124 0.026
R4795 fin.n123 fin.n122 0.026
R4796 fin.n89 fin.n88 0.017
R4797 fin.n94 fin.n92 0.017
R4798 fin.n71 fin.n70 0.017
R4799 fin.n81 fin.n75 0.017
R4800 fin.n22 fin.n18 0.017
R4801 fin.n27 fin.n26 0.017
R4802 fin.n42 fin.n41 0.017
R4803 fin.n52 fin.n45 0.017
R4804 fin.n120 fin.n13 0.017
R4805 fin.n12 fin.n11 0.017
R4806 fin.n3 fin.n2 0.017
R4807 fin.n1 fin.n0 0.017
R4808 fin.n66 fin.n62 0.016
R4809 fin.n115 fin.n114 0.016
R4810 fin.n112 fin.n111 0.016
R4811 fin.n33 fin.n29 0.016
R4812 fin.n38 fin.n37 0.016
R4813 fin.n86 fin.n85 0.015
R4814 fin.n78 fin.n77 0.015
R4815 fin.n20 fin.n19 0.015
R4816 fin.n49 fin.n48 0.015
R4817 fin.n31 fin.n30 0.015
R4818 fin.n40 fin.n39 0.015
R4819 fin.n10 fin.n9 0.015
R4820 fin.n5 fin.n4 0.015
R4821 fin.n128 fin.n127 0.013
R4822 fin.n124 fin.n123 0.013
R4823 fin.n67 fin.n61 0.012
R4824 fin.n67 fin.n66 0.012
R4825 fin.n114 fin.n113 0.012
R4826 fin.n113 fin.n112 0.012
R4827 fin.n34 fin.n33 0.012
R4828 fin.n37 fin.n34 0.012
R4829 fin.n97 fin.n96 0.011
R4830 fin.n74 fin.n73 0.011
R4831 fin.n118 fin.n117 0.011
R4832 fin.n109 fin.n108 0.011
R4833 fin.n25 fin.n24 0.011
R4834 fin.n54 fin.n44 0.011
R4835 fin.n95 fin.n91 0.01
R4836 fin.n116 fin.n115 0.01
R4837 fin.n111 fin.n110 0.01
R4838 fin.n29 fin.n28 0.01
R4839 fin.n43 fin.n38 0.01
R4840 fin.n97 fin.n90 0.006
R4841 fin.n96 fin.n95 0.006
R4842 fin.n73 fin.n72 0.006
R4843 fin.n119 fin.n118 0.006
R4844 fin.n117 fin.n116 0.006
R4845 fin.n110 fin.n109 0.006
R4846 fin.n28 fin.n25 0.006
R4847 fin.n44 fin.n43 0.006
R4848 fin.n54 fin.n53 0.006
R4849 fin.n103 fin.n102 0.004
R4850 fin.n68 fin.n58 0.004
R4851 fin.n24 fin.n23 0.003
R4852 fin.n56 fin.n55 0.003
R4853 fin.n99 fin.n98 0.003
R4854 fin.n106 fin.n105 0.003
R4855 fin.n82 fin.n74 0.003
R4856 fin.n16 fin.n15 0.003
R4857 fin.n108 fin.n107 0.002
R4858 fin.n17 fin.n16 0.002
R4859 fin.n104 fin.n103 0.002
R4860 fin.n83 fin.n68 0.002
R4861 fin.n106 fin.n104 0.002
R4862 fin.n98 fin.n83 0.002
R4863 fin.n55 fin.n17 0.002
R4864 fin.n101 fin.n14 0.002
R4865 1.n257 1.t3 1039.53
R4866 1.n257 1.t2 795.332
R4867 1.n30 1.n29 92.5
R4868 1.n46 1.n45 92.5
R4869 1.n45 1.t1 70.344
R4870 1.n8 1.n7 31.034
R4871 1.n65 1.n64 31.034
R4872 1.n113 1.n112 9.3
R4873 1.n190 1.n189 9.3
R4874 1.n15 1.n14 9.3
R4875 1.n66 1.n65 9.3
R4876 1.n9 1.n8 9.3
R4877 1.n77 1.n76 9.3
R4878 1.n229 1.n228 9.154
R4879 1.n31 1.n30 8.282
R4880 1.n47 1.n46 8.282
R4881 1.n228 1.t0 7.141
R4882 1.n149 1.n148 7.033
R4883 1.n92 1.n91 7.033
R4884 1.n9 1.n5 5.647
R4885 1.n66 1.n62 5.647
R4886 1.n230 1.n229 4.65
R4887 1.n44 1.n43 4.65
R4888 1.n176 1.n175 4.5
R4889 1.n196 1.n195 4.5
R4890 1.n210 1.n209 4.5
R4891 1.n217 1.n214 4.5
R4892 1.n225 1.n224 4.5
R4893 1.n231 1.n227 4.5
R4894 1.n100 1.n97 4.5
R4895 1.n107 1.n106 4.5
R4896 1.n119 1.n118 4.5
R4897 1.n129 1.n128 4.5
R4898 1.n139 1.n138 4.5
R4899 1.n163 1.n162 4.5
R4900 1.n83 1.n81 4.5
R4901 1.n70 1.n67 4.5
R4902 1.n57 1.n55 4.5
R4903 1.n32 1.n31 4.5
R4904 1.n39 1.n38 4.5
R4905 1.n48 1.n47 4.5
R4906 1.n12 1.n11 4.5
R4907 1.n20 1.n19 4.5
R4908 1 1.n257 4.265
R4909 1.n128 1.n125 4.141
R4910 1.n162 1.n161 4.141
R4911 1.n7 1.n6 4.137
R4912 1.n64 1.n63 4.137
R4913 1.n118 1.n115 3.764
R4914 1.n209 1.n207 3.764
R4915 1.n19 1.n17 3.764
R4916 1.n67 1.n60 3.764
R4917 1.n138 1.n135 3.388
R4918 1.n106 1.n105 3.388
R4919 1.n195 1.n194 3.388
R4920 1.n175 1.n174 3.388
R4921 1.n11 1.n10 3.388
R4922 1.n81 1.n80 3.388
R4923 1.n138 1.n137 3.011
R4924 1.n106 1.n103 3.011
R4925 1.n97 1.n95 3.011
R4926 1.n189 1.n188 3.011
R4927 1.n195 1.n193 3.011
R4928 1.n175 1.n173 3.011
R4929 1.n11 1.n9 3.011
R4930 1.n31 1.n28 3.011
R4931 1.n81 1.n79 3.011
R4932 1 1.n256 2.652
R4933 1.n118 1.n117 2.635
R4934 1.n112 1.n111 2.635
R4935 1.n214 1.n213 2.635
R4936 1.n209 1.n208 2.635
R4937 1.n19 1.n18 2.635
R4938 1.n55 1.n54 2.635
R4939 1.n67 1.n66 2.635
R4940 1.n128 1.n127 2.258
R4941 1.n162 1.n160 2.258
R4942 1.n25 1.n0 1.755
R4943 1.n179 1.n150 1.755
R4944 1.n25 1.n24 1.705
R4945 1.n42 1.n41 1.705
R4946 1.n72 1.n71 1.705
R4947 1.n86 1.n85 1.705
R4948 1.n255 1.n144 1.705
R4949 1.n199 1.n198 1.705
R4950 1.n248 1.n247 1.705
R4951 1.n254 1.n253 1.705
R4952 1.n242 1.n241 1.705
R4953 1.n236 1.n235 1.705
R4954 1.n185 1.n184 1.705
R4955 1.n179 1.n178 1.705
R4956 1.n256 1.n86 1.527
R4957 1.n214 1.n212 1.505
R4958 1.n197 1.n196 1.5
R4959 1.n211 1.n210 1.5
R4960 1.n218 1.n217 1.5
R4961 1.n226 1.n225 1.5
R4962 1.n232 1.n231 1.5
R4963 1.n84 1.n83 1.5
R4964 1.n71 1.n70 1.5
R4965 1.n33 1.n32 1.5
R4966 1.n58 1.n57 1.5
R4967 1.n40 1.n39 1.5
R4968 1.n49 1.n48 1.5
R4969 1.n24 1.n12 1.5
R4970 1.n21 1.n20 1.5
R4971 1.n97 1.n96 1.129
R4972 1.n150 1.n149 1.127
R4973 1.n144 1.n92 1.127
R4974 1.n140 1.n139 1.125
R4975 1.n177 1.n176 1.125
R4976 1.n5 1.n4 0.752
R4977 1.n62 1.n61 0.752
R4978 1.n256 1.n255 0.476
R4979 1.n91 1.n90 0.155
R4980 1.n148 1.n147 0.155
R4981 1.n137 1.n136 0.144
R4982 1.n173 1.n172 0.144
R4983 1.n127 1.n126 0.133
R4984 1.n160 1.n159 0.132
R4985 1.n133 1.n132 0.053
R4986 1.n123 1.n122 0.053
R4987 1.n113 1.n110 0.053
R4988 1.n157 1.n156 0.053
R4989 1.n167 1.n166 0.053
R4990 1.n170 1.n169 0.053
R4991 1.n77 1.n75 0.053
R4992 1.n42 1.n25 0.05
R4993 1.n72 1.n42 0.05
R4994 1.n86 1.n72 0.05
R4995 1.n255 1.n254 0.05
R4996 1.n254 1.n248 0.05
R4997 1.n248 1.n242 0.05
R4998 1.n242 1.n236 0.05
R4999 1.n236 1.n200 0.05
R5000 1.n200 1.n199 0.05
R5001 1.n199 1.n185 0.05
R5002 1.n185 1.n179 0.05
R5003 1.n39 1.n37 0.045
R5004 1.n57 1.n53 0.045
R5005 1.n100 1.n99 0.043
R5006 1.n225 1.n223 0.043
R5007 1.n88 1.n87 0.034
R5008 1.n166 1.n165 0.032
R5009 1.n134 1.n133 0.03
R5010 1.n132 1.n131 0.03
R5011 1.n156 1.n155 0.03
R5012 1.n22 1.n21 0.03
R5013 1.n84 1.n74 0.03
R5014 1.n122 1.n121 0.028
R5015 1.n168 1.n167 0.028
R5016 1.n171 1.n170 0.028
R5017 1.n94 1.n93 0.025
R5018 1.n124 1.n123 0.025
R5019 1.n48 1.n44 0.025
R5020 1.n117 1.n116 0.024
R5021 1.n193 1.n192 0.024
R5022 1.n231 1.n230 0.023
R5023 1.n158 1.n157 0.023
R5024 1.n120 1.n119 0.021
R5025 1.n114 1.n113 0.021
R5026 1.n204 1.n203 0.021
R5027 1.n20 1.n13 0.021
R5028 1.n16 1.n15 0.021
R5029 1.n70 1.n59 0.021
R5030 1.n139 1.n94 0.019
R5031 1.n110 1.n109 0.019
R5032 1.n109 1.n108 0.019
R5033 1.n107 1.n102 0.019
R5034 1.n205 1.n204 0.019
R5035 1.n191 1.n190 0.019
R5036 1.n176 1.n171 0.019
R5037 1.n2 1.n1 0.019
R5038 1.n3 1.n2 0.019
R5039 1.n69 1.n68 0.019
R5040 1.n78 1.n77 0.019
R5041 1.n83 1.n82 0.019
R5042 1.n92 1.n89 0.019
R5043 1.n149 1.n146 0.019
R5044 1.n198 1.n197 0.018
R5045 1.n139 1.n134 0.017
R5046 1.n130 1.n129 0.017
R5047 1.n108 1.n107 0.017
R5048 1.n101 1.n100 0.017
R5049 1.n196 1.n191 0.017
R5050 1.n164 1.n163 0.017
R5051 1.n176 1.n168 0.017
R5052 1.n12 1.n3 0.017
R5053 1.n32 1.n27 0.017
R5054 1.n83 1.n78 0.017
R5055 1.n142 1.n141 0.016
R5056 1.n252 1.n251 0.016
R5057 1.n246 1.n245 0.016
R5058 1.n181 1.n180 0.016
R5059 1.n153 1.n152 0.016
R5060 1.n71 1.n58 0.016
R5061 1.n119 1.n114 0.015
R5062 1.n217 1.n216 0.015
R5063 1.n210 1.n205 0.015
R5064 1.n238 1.n237 0.015
R5065 1.n232 1.n226 0.015
R5066 1.n218 1.n211 0.015
R5067 1.n20 1.n16 0.015
R5068 1.n57 1.n56 0.015
R5069 1.n70 1.n69 0.015
R5070 1.n40 1.n35 0.015
R5071 1.n58 1.n51 0.015
R5072 1.n177 1.n153 0.014
R5073 1.n34 1.n33 0.014
R5074 1.n50 1.n49 0.014
R5075 1.n141 1.n140 0.013
R5076 1.n233 1.n232 0.013
R5077 1.n226 1.n221 0.013
R5078 1.n105 1.n104 0.012
R5079 1.n207 1.n206 0.012
R5080 1.n129 1.n124 0.012
R5081 1.n102 1.n101 0.012
R5082 1.n216 1.n215 0.012
R5083 1.n163 1.n158 0.012
R5084 1.n27 1.n26 0.012
R5085 1.n143 1.n142 0.011
R5086 1.n251 1.n250 0.011
R5087 1.n239 1.n238 0.011
R5088 1.n219 1.n218 0.011
R5089 1.n182 1.n181 0.011
R5090 1.n152 1.n151 0.011
R5091 1.n24 1.n23 0.011
R5092 1.n211 1.n202 0.01
R5093 1.n184 1.n183 0.01
R5094 1.n253 1.n252 0.009
R5095 1.n241 1.n240 0.009
R5096 1.n187 1.n186 0.009
R5097 1.n99 1.n98 0.008
R5098 1.n223 1.n222 0.008
R5099 1.n245 1.n244 0.008
R5100 1.n244 1.n243 0.008
R5101 1.n37 1.n36 0.008
R5102 1.n53 1.n52 0.008
R5103 1.n85 1.n84 0.008
R5104 1.n197 1.n187 0.007
R5105 1.n41 1.n40 0.007
R5106 1.n74 1.n73 0.007
R5107 1.n131 1.n130 0.006
R5108 1.n121 1.n120 0.006
R5109 1.n155 1.n154 0.006
R5110 1.n165 1.n164 0.006
R5111 1.n202 1.n201 0.006
R5112 1.n23 1.n22 0.006
R5113 1.n144 1.n143 0.005
R5114 1.n250 1.n249 0.005
R5115 1.n240 1.n239 0.005
R5116 1.n183 1.n182 0.005
R5117 1.n178 1.n177 0.005
R5118 1.n89 1.n88 0.004
R5119 1.n146 1.n145 0.004
R5120 1.n235 1.n234 0.002
R5121 1.n234 1.n233 0.002
R5122 1.n221 1.n220 0.002
R5123 1.n220 1.n219 0.002
R5124 1.n35 1.n34 0.002
R5125 1.n51 1.n50 0.002
R5126 1.n247 1.n246 0.001
R5127 net2_ff1.n35 net2_ff1.n34 92.5
R5128 net2_ff1.n33 net2_ff1.n32 92.5
R5129 net2_ff1.n28 net2_ff1.n27 92.5
R5130 net2_ff1.n30 net2_ff1.n29 92.5
R5131 net2_ff1.n34 net2_ff1.t0 70.344
R5132 net2_ff1.n27 net2_ff1.t1 70.344
R5133 net2_ff1.n17 net2_ff1.n16 31.034
R5134 net2_ff1.n49 net2_ff1.n48 31.034
R5135 net2_ff1.n23 net2_ff1.n22 31.034
R5136 net2_ff1.n43 net2_ff1.n42 31.034
R5137 net2_ff1.n36 net2_ff1.n33 12.8
R5138 net2_ff1.n36 net2_ff1.n35 12.8
R5139 net2_ff1.n31 net2_ff1.n28 12.8
R5140 net2_ff1.n31 net2_ff1.n30 12.8
R5141 net2_ff1.n12 net2_ff1.n10 9.3
R5142 net2_ff1.n6 net2_ff1.n4 9.3
R5143 net2_ff1.n25 net2_ff1.n18 9.3
R5144 net2_ff1.n18 net2_ff1.n17 9.3
R5145 net2_ff1.n60 net2_ff1.n52 9.3
R5146 net2_ff1.n60 net2_ff1.n59 9.3
R5147 net2_ff1.n51 net2_ff1.n44 9.3
R5148 net2_ff1.n44 net2_ff1.n43 9.3
R5149 net2_ff1.n51 net2_ff1.n50 9.3
R5150 net2_ff1.n50 net2_ff1.n49 9.3
R5151 net2_ff1.n25 net2_ff1.n24 9.3
R5152 net2_ff1.n24 net2_ff1.n23 9.3
R5153 net2_ff1.n56 net2_ff1.n54 9.3
R5154 net2_ff1.n58 net2_ff1.n53 9.3
R5155 net2_ff1.n58 net2_ff1.n57 9.3
R5156 net2_ff1.n56 net2_ff1.n55 9.3
R5157 net2_ff1.n12 net2_ff1.n11 9.3
R5158 net2_ff1.n9 net2_ff1.n7 9.3
R5159 net2_ff1.n9 net2_ff1.n8 9.3
R5160 net2_ff1.n6 net2_ff1.n5 9.3
R5161 net2_ff1.n18 net2_ff1.n14 5.647
R5162 net2_ff1.n50 net2_ff1.n46 5.647
R5163 net2_ff1.n24 net2_ff1.n20 5.647
R5164 net2_ff1.n44 net2_ff1.n40 5.647
R5165 net2_ff1.n37 net2_ff1.n31 4.65
R5166 net2_ff1.n37 net2_ff1.n36 4.65
R5167 net2_ff1.n26 net2_ff1.n3 4.47
R5168 net2_ff1.n38 net2_ff1.n1 4.47
R5169 net2_ff1.n38 net2_ff1.n0 4.47
R5170 net2_ff1.n26 net2_ff1.n2 4.47
R5171 net2_ff1.n16 net2_ff1.n15 4.137
R5172 net2_ff1.n48 net2_ff1.n47 4.137
R5173 net2_ff1.n22 net2_ff1.n21 4.137
R5174 net2_ff1.n42 net2_ff1.n41 4.137
R5175 net2_ff1.n14 net2_ff1.n13 0.752
R5176 net2_ff1.n46 net2_ff1.n45 0.752
R5177 net2_ff1.n20 net2_ff1.n19 0.752
R5178 net2_ff1.n40 net2_ff1.n39 0.752
R5179 net2_ff1.n37 net2_ff1.n26 0.032
R5180 net2_ff1.n38 net2_ff1.n37 0.032
R5181 net2_ff1.n25 net2_ff1.n12 0.024
R5182 net2_ff1 net2_ff1.n51 0.019
R5183 net2_ff1.n26 net2_ff1.n25 0.007
R5184 net2_ff1.n51 net2_ff1.n38 0.007
R5185 net2_ff1.n9 net2_ff1.n6 0.006
R5186 net2_ff1.n58 net2_ff1.n56 0.006
R5187 net2_ff1 net2_ff1.n60 0.005
R5188 net2_ff1.n12 net2_ff1.n9 0.001
R5189 net2_ff1.n60 net2_ff1.n58 0.001
R5190 net4_ff2.n65 net4_ff2.n63 9.3
R5191 net4_ff2.n65 net4_ff2.n64 9.3
R5192 net4_ff2.n68 net4_ff2.n62 9.3
R5193 net4_ff2.n2 net4_ff2.n0 9.3
R5194 net4_ff2.n98 net4_ff2.n4 9.3
R5195 net4_ff2.n93 net4_ff2.n6 9.3
R5196 net4_ff2.n95 net4_ff2.n5 9.3
R5197 net4_ff2.n68 net4_ff2.n67 9.3
R5198 net4_ff2.n2 net4_ff2.n1 9.3
R5199 net4_ff2.n98 net4_ff2.n97 9.3
R5200 net4_ff2.n93 net4_ff2.n92 9.3
R5201 net4_ff2.n95 net4_ff2.n94 9.3
R5202 net4_ff2.n89 net4_ff2.n84 8.907
R5203 net4_ff2.n33 net4_ff2.n28 8.907
R5204 net4_ff2.n33 net4_ff2.n19 8.897
R5205 net4_ff2.n33 net4_ff2.n32 8.896
R5206 net4_ff2.n89 net4_ff2.n47 8.896
R5207 net4_ff2.n89 net4_ff2.n88 8.896
R5208 net4_ff2.n89 net4_ff2.n43 8.886
R5209 net4_ff2.n33 net4_ff2.n15 8.886
R5210 net4_ff2.n33 net4_ff2.n11 8.875
R5211 net4_ff2.n89 net4_ff2.n39 8.875
R5212 net4_ff2.n34 net4_ff2.n33 8.864
R5213 net4_ff2.n33 net4_ff2.n7 8.864
R5214 net4_ff2.n90 net4_ff2.n89 8.864
R5215 net4_ff2.n89 net4_ff2.n35 8.864
R5216 net4_ff2.n33 net4_ff2.t1 7.141
R5217 net4_ff2.n89 net4_ff2.t3 7.141
R5218 net4_ff2.n22 net4_ff2.n21 5.647
R5219 net4_ff2.n26 net4_ff2.n25 5.647
R5220 net4_ff2.n78 net4_ff2.n77 5.647
R5221 net4_ff2.n82 net4_ff2.n81 5.647
R5222 net4_ff2.n24 net4_ff2.n20 5.418
R5223 net4_ff2.n80 net4_ff2.n76 5.418
R5224 net4_ff2.n24 net4_ff2.n23 5.38
R5225 net4_ff2.n80 net4_ff2.n79 5.38
R5226 net4_ff2.n17 net4_ff2.n16 4.894
R5227 net4_ff2.n30 net4_ff2.n29 4.894
R5228 net4_ff2.n45 net4_ff2.n44 4.894
R5229 net4_ff2.n86 net4_ff2.n85 4.894
R5230 net4_ff2.n91 net4_ff2.n34 4.728
R5231 net4_ff2.n91 net4_ff2.n90 4.728
R5232 net4_ff2.n76 net4_ff2.n75 4.65
R5233 net4_ff2.n13 net4_ff2.n12 4.141
R5234 net4_ff2.n41 net4_ff2.n40 4.141
R5235 net4_ff2.n9 net4_ff2.n8 3.388
R5236 net4_ff2.n37 net4_ff2.n36 3.388
R5237 net4_ff2.n10 net4_ff2.n9 3.011
R5238 net4_ff2.n38 net4_ff2.n37 3.011
R5239 net4_ff2.n14 net4_ff2.n13 2.258
R5240 net4_ff2.n42 net4_ff2.n41 2.258
R5241 net4_ff2.n89 net4_ff2.n80 1.844
R5242 net4_ff2.n33 net4_ff2.n24 1.844
R5243 net4_ff2.n18 net4_ff2.n17 1.505
R5244 net4_ff2.n31 net4_ff2.n30 1.505
R5245 net4_ff2.n46 net4_ff2.n45 1.505
R5246 net4_ff2.n87 net4_ff2.n86 1.505
R5247 net4_ff2.n23 net4_ff2.n22 0.752
R5248 net4_ff2.n27 net4_ff2.n26 0.752
R5249 net4_ff2.n79 net4_ff2.n78 0.752
R5250 net4_ff2.n83 net4_ff2.n82 0.752
R5251 net4_ff2.n11 net4_ff2.n10 0.144
R5252 net4_ff2.n39 net4_ff2.n38 0.144
R5253 net4_ff2.n4 net4_ff2.n3 0.144
R5254 net4_ff2.n97 net4_ff2.n96 0.144
R5255 net4_ff2.n15 net4_ff2.n14 0.133
R5256 net4_ff2.n43 net4_ff2.n42 0.133
R5257 net4_ff2.n62 net4_ff2.n61 0.133
R5258 net4_ff2.n67 net4_ff2.n66 0.132
R5259 net4_ff2.n19 net4_ff2.n18 0.121
R5260 net4_ff2.n47 net4_ff2.n46 0.121
R5261 net4_ff2.n88 net4_ff2.n87 0.121
R5262 net4_ff2.n32 net4_ff2.n31 0.121
R5263 net4_ff2.n84 net4_ff2.n83 0.11
R5264 net4_ff2.n28 net4_ff2.n27 0.109
R5265 net4_ff2.n75 net4_ff2.n60 0.035
R5266 net4_ff2.n75 net4_ff2.n74 0.035
R5267 net4_ff2.n49 net4_ff2.n48 0.029
R5268 net4_ff2.n93 net4_ff2.n91 0.029
R5269 net4_ff2.n52 net4_ff2.n51 0.027
R5270 net4_ff2.n55 net4_ff2.n54 0.027
R5271 net4_ff2.n58 net4_ff2.n57 0.027
R5272 net4_ff2.n72 net4_ff2.n71 0.027
R5273 net1_ff2 net4_ff2.n98 0.019
R5274 net4_ff2.n69 net4_ff2 0.018
R5275 net4_ff2 net4_ff2.n68 0.008
R5276 net4_ff2.n59 net4_ff2.n58 0.007
R5277 net4_ff2.n73 net4_ff2.n72 0.007
R5278 net1_ff2 net4_ff2.n2 0.007
R5279 net4_ff2.n56 net4_ff2.n55 0.006
R5280 net4_ff2.n70 net4_ff2.n69 0.006
R5281 net4_ff2.n53 net4_ff2.n52 0.005
R5282 net4_ff2.n65 net4_ff2.n2 0.005
R5283 net4_ff2.n50 net4_ff2.n49 0.004
R5284 net4_ff2.n51 net4_ff2.n50 0.004
R5285 net4_ff2.n98 net4_ff2.n95 0.004
R5286 net4_ff2.n95 net4_ff2.n93 0.004
R5287 net4_ff2.n54 net4_ff2.n53 0.003
R5288 net4_ff2.n68 net4_ff2.n65 0.003
R5289 net4_ff2.n57 net4_ff2.n56 0.002
R5290 net4_ff2.n71 net4_ff2.n70 0.002
R5291 net4_ff2.n60 net4_ff2.n59 0.001
R5292 net4_ff2.n74 net4_ff2.n73 0.001
R5293 net2_ff2.n40 net2_ff2.n39 92.5
R5294 net2_ff2.n38 net2_ff2.n37 92.5
R5295 net2_ff2.n32 net2_ff2.n31 92.5
R5296 net2_ff2.n34 net2_ff2.n33 92.5
R5297 net2_ff2.n39 net2_ff2.t1 70.344
R5298 net2_ff2.n33 net2_ff2.t0 70.344
R5299 net2_ff2.n26 net2_ff2.n25 31.034
R5300 net2_ff2.n56 net2_ff2.n55 31.034
R5301 net2_ff2.n19 net2_ff2.n18 31.034
R5302 net2_ff2.n49 net2_ff2.n48 31.034
R5303 net2_ff2.n41 net2_ff2.n38 12.8
R5304 net2_ff2.n41 net2_ff2.n40 12.8
R5305 net2_ff2.n35 net2_ff2.n32 12.8
R5306 net2_ff2.n35 net2_ff2.n34 12.8
R5307 net2_ff2.n6 net2_ff2.n4 9.303
R5308 net2_ff2.n61 net2_ff2.n59 9.303
R5309 net2_ff2.n10 net2_ff2.n9 9.3
R5310 net2_ff2.n6 net2_ff2.n5 9.3
R5311 net2_ff2.n28 net2_ff2.n27 9.3
R5312 net2_ff2.n27 net2_ff2.n26 9.3
R5313 net2_ff2.n65 net2_ff2.n64 9.3
R5314 net2_ff2.n69 net2_ff2.n68 9.3
R5315 net2_ff2.n51 net2_ff2.n50 9.3
R5316 net2_ff2.n50 net2_ff2.n49 9.3
R5317 net2_ff2.n58 net2_ff2.n57 9.3
R5318 net2_ff2.n57 net2_ff2.n56 9.3
R5319 net2_ff2.n21 net2_ff2.n20 9.3
R5320 net2_ff2.n20 net2_ff2.n19 9.3
R5321 net2_ff2.n61 net2_ff2.n60 9.3
R5322 net2_ff2.n67 net2_ff2.n66 9.3
R5323 net2_ff2.n63 net2_ff2.n62 9.3
R5324 net2_ff2.n14 net2_ff2.n13 9.3
R5325 net2_ff2.n12 net2_ff2.n11 9.3
R5326 net2_ff2.n8 net2_ff2.n7 9.3
R5327 net2_ff2.n27 net2_ff2.n23 5.647
R5328 net2_ff2.n57 net2_ff2.n53 5.647
R5329 net2_ff2.n20 net2_ff2.n16 5.647
R5330 net2_ff2.n50 net2_ff2.n46 5.647
R5331 net2_ff2.n36 net2_ff2.n35 4.65
R5332 net2_ff2.n42 net2_ff2.n41 4.65
R5333 net2_ff2.n29 net2_ff2.n3 4.47
R5334 net2_ff2.n43 net2_ff2.n1 4.47
R5335 net2_ff2.n44 net2_ff2.n0 4.47
R5336 net2_ff2.n30 net2_ff2.n2 4.47
R5337 net2_ff2.n25 net2_ff2.n24 4.137
R5338 net2_ff2.n55 net2_ff2.n54 4.137
R5339 net2_ff2.n18 net2_ff2.n17 4.137
R5340 net2_ff2.n48 net2_ff2.n47 4.137
R5341 net2_ff2.n23 net2_ff2.n22 0.752
R5342 net2_ff2.n53 net2_ff2.n52 0.752
R5343 net2_ff2.n16 net2_ff2.n15 0.752
R5344 net2_ff2.n46 net2_ff2.n45 0.752
R5345 net2_ff2.n36 net2_ff2.n30 0.029
R5346 net2_ff2.n43 net2_ff2.n42 0.029
R5347 net2_ff2.n21 net2_ff2.n14 0.021
R5348 net2_ff2 net2_ff2.n69 0.013
R5349 net2_ff2 net2_ff2.n58 0.008
R5350 net2_ff2.n28 net2_ff2.n21 0.003
R5351 net2_ff2.n29 net2_ff2.n28 0.003
R5352 net2_ff2.n42 net2_ff2.n36 0.003
R5353 net2_ff2.n51 net2_ff2.n44 0.003
R5354 net2_ff2.n58 net2_ff2.n51 0.003
R5355 net2_ff2.n8 net2_ff2.n6 0.002
R5356 net2_ff2.n30 net2_ff2.n29 0.002
R5357 net2_ff2.n44 net2_ff2.n43 0.002
R5358 net2_ff2.n63 net2_ff2.n61 0.002
R5359 net2_ff2.n10 net2_ff2.n8 0.001
R5360 net2_ff2.n12 net2_ff2.n10 0.001
R5361 net2_ff2.n14 net2_ff2.n12 0.001
R5362 net2_ff2.n69 net2_ff2.n67 0.001
R5363 net2_ff2.n67 net2_ff2.n65 0.001
R5364 net2_ff2.n65 net2_ff2.n63 0.001
R5365 net5_ff1.n35 net5_ff1.n34 92.5
R5366 net5_ff1.n33 net5_ff1.n32 92.5
R5367 net5_ff1.n28 net5_ff1.n27 92.5
R5368 net5_ff1.n30 net5_ff1.n29 92.5
R5369 net5_ff1.n34 net5_ff1.t0 70.344
R5370 net5_ff1.n27 net5_ff1.t1 70.344
R5371 net5_ff1.n17 net5_ff1.n16 31.034
R5372 net5_ff1.n49 net5_ff1.n48 31.034
R5373 net5_ff1.n23 net5_ff1.n22 31.034
R5374 net5_ff1.n43 net5_ff1.n42 31.034
R5375 net5_ff1.n36 net5_ff1.n33 12.8
R5376 net5_ff1.n36 net5_ff1.n35 12.8
R5377 net5_ff1.n31 net5_ff1.n28 12.8
R5378 net5_ff1.n31 net5_ff1.n30 12.8
R5379 net5_ff1.n12 net5_ff1.n10 9.3
R5380 net5_ff1.n6 net5_ff1.n4 9.3
R5381 net5_ff1.n25 net5_ff1.n18 9.3
R5382 net5_ff1.n18 net5_ff1.n17 9.3
R5383 net5_ff1.n60 net5_ff1.n52 9.3
R5384 net5_ff1.n60 net5_ff1.n59 9.3
R5385 net5_ff1.n51 net5_ff1.n44 9.3
R5386 net5_ff1.n44 net5_ff1.n43 9.3
R5387 net5_ff1.n51 net5_ff1.n50 9.3
R5388 net5_ff1.n50 net5_ff1.n49 9.3
R5389 net5_ff1.n25 net5_ff1.n24 9.3
R5390 net5_ff1.n24 net5_ff1.n23 9.3
R5391 net5_ff1.n56 net5_ff1.n54 9.3
R5392 net5_ff1.n58 net5_ff1.n53 9.3
R5393 net5_ff1.n58 net5_ff1.n57 9.3
R5394 net5_ff1.n56 net5_ff1.n55 9.3
R5395 net5_ff1.n12 net5_ff1.n11 9.3
R5396 net5_ff1.n9 net5_ff1.n7 9.3
R5397 net5_ff1.n9 net5_ff1.n8 9.3
R5398 net5_ff1.n6 net5_ff1.n5 9.3
R5399 net5_ff1.n18 net5_ff1.n14 5.647
R5400 net5_ff1.n50 net5_ff1.n46 5.647
R5401 net5_ff1.n24 net5_ff1.n20 5.647
R5402 net5_ff1.n44 net5_ff1.n40 5.647
R5403 net5_ff1.n37 net5_ff1.n31 4.65
R5404 net5_ff1.n37 net5_ff1.n36 4.65
R5405 net5_ff1.n26 net5_ff1.n3 4.47
R5406 net5_ff1.n38 net5_ff1.n1 4.47
R5407 net5_ff1.n38 net5_ff1.n0 4.47
R5408 net5_ff1.n26 net5_ff1.n2 4.47
R5409 net5_ff1.n16 net5_ff1.n15 4.137
R5410 net5_ff1.n48 net5_ff1.n47 4.137
R5411 net5_ff1.n22 net5_ff1.n21 4.137
R5412 net5_ff1.n42 net5_ff1.n41 4.137
R5413 net5_ff1.n14 net5_ff1.n13 0.752
R5414 net5_ff1.n46 net5_ff1.n45 0.752
R5415 net5_ff1.n20 net5_ff1.n19 0.752
R5416 net5_ff1.n40 net5_ff1.n39 0.752
R5417 net5_ff1.n37 net5_ff1.n26 0.032
R5418 net5_ff1.n38 net5_ff1.n37 0.032
R5419 net5_ff1.n25 net5_ff1.n12 0.024
R5420 net5_ff1 net5_ff1.n51 0.016
R5421 net5_ff1 net5_ff1.n60 0.008
R5422 net5_ff1.n26 net5_ff1.n25 0.006
R5423 net5_ff1.n51 net5_ff1.n38 0.006
R5424 net5_ff1.n9 net5_ff1.n6 0.005
R5425 net5_ff1.n58 net5_ff1.n56 0.005
R5426 net5_ff1.n12 net5_ff1.n9 0.001
R5427 net5_ff1.n60 net5_ff1.n58 0.001
R5428 net1_ff2.n75 net1_ff2.n74 50.948
R5429 net1_ff2.n93 net1_ff2.n92 50.948
R5430 net1_ff2.n69 net1_ff2.n68 50.948
R5431 net1_ff2.n87 net1_ff2.n86 50.948
R5432 net1_ff2.n50 net1_ff2.n49 44.155
R5433 net1_ff2.n112 net1_ff2.n111 44.155
R5434 net1_ff2.n56 net1_ff2.n55 44.155
R5435 net1_ff2.n106 net1_ff2.n105 44.155
R5436 net1_ff2.n37 net1_ff2.n36 37.362
R5437 net1_ff2.n159 net1_ff2.n158 37.362
R5438 net1_ff2.n31 net1_ff2.n30 37.362
R5439 net1_ff2.n125 net1_ff2.n124 37.362
R5440 net1_ff2.n18 net1_ff2.n17 30.568
R5441 net1_ff2.n148 net1_ff2.n147 30.568
R5442 net1_ff2.n12 net1_ff2.n11 30.568
R5443 net1_ff2.n133 net1_ff2.n132 30.568
R5444 net1_ff2.n19 net1_ff2.n18 27.172
R5445 net1_ff2.n149 net1_ff2.n148 27.172
R5446 net1_ff2.n13 net1_ff2.n12 27.172
R5447 net1_ff2.n134 net1_ff2.n133 27.172
R5448 net1_ff2.n38 net1_ff2.n37 20.379
R5449 net1_ff2.n160 net1_ff2.n159 20.379
R5450 net1_ff2.n32 net1_ff2.n31 20.379
R5451 net1_ff2.n126 net1_ff2.n125 20.379
R5452 net1_ff2.n51 net1_ff2.n50 13.586
R5453 net1_ff2.n113 net1_ff2.n112 13.586
R5454 net1_ff2.n57 net1_ff2.n56 13.586
R5455 net1_ff2.n107 net1_ff2.n106 13.586
R5456 net1_ff2.n21 net1_ff2.n14 9.3
R5457 net1_ff2.n14 net1_ff2.n13 9.3
R5458 net1_ff2.n5 net1_ff2.n3 9.3
R5459 net1_ff2.n40 net1_ff2.n33 9.3
R5460 net1_ff2.n33 net1_ff2.n32 9.3
R5461 net1_ff2.n24 net1_ff2.n22 9.3
R5462 net1_ff2.n59 net1_ff2.n52 9.3
R5463 net1_ff2.n52 net1_ff2.n51 9.3
R5464 net1_ff2.n46 net1_ff2.n44 9.3
R5465 net1_ff2.n65 net1_ff2.n63 9.3
R5466 net1_ff2.n65 net1_ff2.n64 9.3
R5467 net1_ff2.n99 net1_ff2.n97 9.3
R5468 net1_ff2.n99 net1_ff2.n98 9.3
R5469 net1_ff2.n118 net1_ff2.n116 9.3
R5470 net1_ff2.n118 net1_ff2.n117 9.3
R5471 net1_ff2.n155 net1_ff2.n128 9.3
R5472 net1_ff2.n155 net1_ff2.n154 9.3
R5473 net1_ff2.n43 net1_ff2.n41 9.3
R5474 net1_ff2.n59 net1_ff2.n58 9.3
R5475 net1_ff2.n58 net1_ff2.n57 9.3
R5476 net1_ff2.n62 net1_ff2.n60 9.3
R5477 net1_ff2.n78 net1_ff2.n71 9.3
R5478 net1_ff2.n71 net1_ff2.n70 9.3
R5479 net1_ff2.n96 net1_ff2.n89 9.3
R5480 net1_ff2.n89 net1_ff2.n88 9.3
R5481 net1_ff2.n102 net1_ff2.n100 9.3
R5482 net1_ff2.n115 net1_ff2.n108 9.3
R5483 net1_ff2.n108 net1_ff2.n107 9.3
R5484 net1_ff2.n121 net1_ff2.n119 9.3
R5485 net1_ff2.n162 net1_ff2.n127 9.3
R5486 net1_ff2.n127 net1_ff2.n126 9.3
R5487 net1_ff2.n153 net1_ff2.n129 9.3
R5488 net1_ff2.n151 net1_ff2.n135 9.3
R5489 net1_ff2.n135 net1_ff2.n134 9.3
R5490 net1_ff2.n142 net1_ff2.n137 9.3
R5491 net1_ff2.n144 net1_ff2.n136 9.3
R5492 net1_ff2.n62 net1_ff2.n61 9.3
R5493 net1_ff2.n78 net1_ff2.n77 9.3
R5494 net1_ff2.n77 net1_ff2.n76 9.3
R5495 net1_ff2.n96 net1_ff2.n95 9.3
R5496 net1_ff2.n95 net1_ff2.n94 9.3
R5497 net1_ff2.n102 net1_ff2.n101 9.3
R5498 net1_ff2.n115 net1_ff2.n114 9.3
R5499 net1_ff2.n114 net1_ff2.n113 9.3
R5500 net1_ff2.n121 net1_ff2.n120 9.3
R5501 net1_ff2.n162 net1_ff2.n161 9.3
R5502 net1_ff2.n161 net1_ff2.n160 9.3
R5503 net1_ff2.n153 net1_ff2.n152 9.3
R5504 net1_ff2.n151 net1_ff2.n150 9.3
R5505 net1_ff2.n150 net1_ff2.n149 9.3
R5506 net1_ff2.n142 net1_ff2.n141 9.3
R5507 net1_ff2.n144 net1_ff2.n143 9.3
R5508 net1_ff2.n46 net1_ff2.n45 9.3
R5509 net1_ff2.n43 net1_ff2.n42 9.3
R5510 net1_ff2.n40 net1_ff2.n39 9.3
R5511 net1_ff2.n39 net1_ff2.n38 9.3
R5512 net1_ff2.n27 net1_ff2.n25 9.3
R5513 net1_ff2.n27 net1_ff2.n26 9.3
R5514 net1_ff2.n24 net1_ff2.n23 9.3
R5515 net1_ff2.n21 net1_ff2.n20 9.3
R5516 net1_ff2.n20 net1_ff2.n19 9.3
R5517 net1_ff2.n8 net1_ff2.n6 9.3
R5518 net1_ff2.n8 net1_ff2.n7 9.3
R5519 net1_ff2.n5 net1_ff2.n4 9.3
R5520 net1_ff2.n80 net1_ff2.n79 9.154
R5521 net1_ff2.n82 net1_ff2.n81 9.154
R5522 net1_ff2.n76 net1_ff2.n75 6.793
R5523 net1_ff2.n94 net1_ff2.n93 6.793
R5524 net1_ff2.n70 net1_ff2.n69 6.793
R5525 net1_ff2.n88 net1_ff2.n87 6.793
R5526 net1_ff2.n73 net1_ff2.n72 5.647
R5527 net1_ff2.n91 net1_ff2.n90 5.647
R5528 net1_ff2.n67 net1_ff2.n66 5.647
R5529 net1_ff2.n85 net1_ff2.n84 5.647
R5530 net1_ff2.n2 net1_ff2.n0 5.428
R5531 net1_ff2.n140 net1_ff2.n138 5.428
R5532 net1_ff2.n140 net1_ff2.n139 5.427
R5533 net1_ff2.n2 net1_ff2.n1 5.427
R5534 net1_ff2.n48 net1_ff2.n47 4.894
R5535 net1_ff2.n110 net1_ff2.n109 4.894
R5536 net1_ff2.n54 net1_ff2.n53 4.894
R5537 net1_ff2.n104 net1_ff2.n103 4.894
R5538 net1_ff2.n83 net1_ff2.n80 4.65
R5539 net1_ff2.n83 net1_ff2.n82 4.65
R5540 net1_ff2.n35 net1_ff2.n34 4.141
R5541 net1_ff2.n157 net1_ff2.n156 4.141
R5542 net1_ff2.n29 net1_ff2.n28 4.141
R5543 net1_ff2.n123 net1_ff2.n122 4.141
R5544 net1_ff2.n16 net1_ff2.n15 3.388
R5545 net1_ff2.n146 net1_ff2.n145 3.388
R5546 net1_ff2.n10 net1_ff2.n9 3.388
R5547 net1_ff2.n131 net1_ff2.n130 3.388
R5548 net1_ff2.n20 net1_ff2.n16 3.011
R5549 net1_ff2.n150 net1_ff2.n146 3.011
R5550 net1_ff2.n14 net1_ff2.n10 3.011
R5551 net1_ff2.n135 net1_ff2.n131 3.011
R5552 net1_ff2.n39 net1_ff2.n35 2.258
R5553 net1_ff2.n161 net1_ff2.n157 2.258
R5554 net1_ff2.n33 net1_ff2.n29 2.258
R5555 net1_ff2.n127 net1_ff2.n123 2.258
R5556 net1_ff2.n52 net1_ff2.n48 1.505
R5557 net1_ff2.n114 net1_ff2.n110 1.505
R5558 net1_ff2.n58 net1_ff2.n54 1.505
R5559 net1_ff2.n108 net1_ff2.n104 1.505
R5560 net1_ff2.n77 net1_ff2.n73 0.752
R5561 net1_ff2.n95 net1_ff2.n91 0.752
R5562 net1_ff2.n71 net1_ff2.n67 0.752
R5563 net1_ff2.n89 net1_ff2.n85 0.752
R5564 net1_ff2.n83 net1_ff2.n78 0.035
R5565 net1_ff2.n96 net1_ff2.n83 0.035
R5566 net1_ff2.n5 net1_ff2.n2 0.029
R5567 net1_ff2.n142 net1_ff2.n140 0.029
R5568 net1_ff2.n24 net1_ff2.n21 0.027
R5569 net1_ff2.n43 net1_ff2.n40 0.027
R5570 net1_ff2.n62 net1_ff2.n59 0.027
R5571 net1_ff2.n115 net1_ff2.n102 0.027
R5572 net1_ff2.n153 net1_ff2.n151 0.027
R5573 net1_ff2 net1_ff2.n121 0.024
R5574 net1_ff2.n65 net1_ff2.n62 0.007
R5575 net1_ff2.n102 net1_ff2.n99 0.007
R5576 net1_ff2.n46 net1_ff2.n43 0.006
R5577 net1_ff2.n121 net1_ff2.n118 0.006
R5578 net1_ff2.n27 net1_ff2.n24 0.005
R5579 net1_ff2.n155 net1_ff2.n153 0.005
R5580 net1_ff2.n8 net1_ff2.n5 0.004
R5581 net1_ff2.n21 net1_ff2.n8 0.004
R5582 net1_ff2.n151 net1_ff2.n144 0.004
R5583 net1_ff2.n144 net1_ff2.n142 0.004
R5584 net1_ff2.n40 net1_ff2.n27 0.003
R5585 net1_ff2 net1_ff2.n162 0.003
R5586 net1_ff2.n162 net1_ff2.n155 0.003
R5587 net1_ff2.n59 net1_ff2.n46 0.002
R5588 net1_ff2.n118 net1_ff2.n115 0.002
R5589 net1_ff2.n78 net1_ff2.n65 0.001
R5590 net1_ff2.n99 net1_ff2.n96 0.001
C0 1 net3_ff1 0.84fF
C1 fin net4_ff1 0.04fF
C2 fout modi 0.96fF
C3 modo net1_ff2 0.06fF
C4 net1 net2_nand3 0.02fF
C5 3 modo 0.53fF
C6 finb 1 0.62fF
C7 net5_ff2 31 0.03fF
C8 finb net5_ff2 0.02fF
C9 net3_ff2 net4_ff1 0.07fF
C10 VDD fin 1.49fF
C11 net5_ff1 net3_ff2 0.04fF
C12 3 net2_ff2 0.01fF
C13 2 VDD 4.56fF
C14 modo P 0.56fF
C15 fout net3_ff1 0.25fF
C16 fin net1_ff2 0.04fF
C17 fout 31 1.16fF
C18 net3_ff2 VDD 1.27fF
C19 3 fin 0.37fF
C20 net1 1 0.03fF
C21 finb fout 2.72fF
C22 net2_ff2 modo 0.05fF
C23 modi 31 0.46fF
C24 1 net4_ff2 0.06fF
C25 finb modi 0.14fF
C26 net3_ff2 net1_ff2 0.66fF
C27 P fin 0.89fF
C28 3 net3_ff2 0.21fF
C29 2 P 0.39fF
C30 modo fin 1.17fF
C31 modo 2 0.80fF
C32 1 net1_ff1 0.09fF
C33 fout net2 0.05fF
C34 net2_ff2 fin 0.05fF
C35 net2_ff1 1 0.04fF
C36 finb net3_ff1 0.87fF
C37 net3_ff2 modo 0.79fF
C38 net1 fout 1.07fF
C39 modi net2 0.06fF
C40 finb 31 0.18fF
C41 net2_ff2 net3_ff2 0.33fF
C42 2 fin 0.60fF
C43 net1_nand3 P 0.02fF
C44 a_n100_n729# VDD 0.03fF
C45 modo net1_nand3 0.07fF
C46 fout net1_ff1 0.03fF
C47 1 net4_ff1 0.67fF
C48 net3_ff2 fin 0.75fF
C49 net1 net3_ff1 0.04fF
C50 net5_ff1 1 0.34fF
C51 net2_ff1 fout 0.04fF
C52 31 net2 1.06fF
C53 finb net2 0.01fF
C54 finb net1 0.08fF
C55 31 net4_ff2 0.04fF
C56 net1_nand3 fin 0.03fF
C57 1 VDD 1.21fF
C58 modo net2_nand3 0.09fF
C59 2 net1_nand3 1.00fF
C60 1 net1_ff2 0.12fF
C61 net3_ff1 net1_ff1 0.66fF
C62 net2_ff1 net3_ff1 0.35fF
C63 3 1 0.09fF
C64 finb net1_ff1 0.12fF
C65 3 net5_ff2 0.03fF
C66 finb net2_ff1 0.07fF
C67 fout VDD 3.20fF
C68 1 P 0.01fF
C69 net2_nand3 fin 0.04fF
C70 modo 1 0.25fF
C71 2 net2_nand3 0.12fF
C72 VDD modi 0.24fF
C73 modo net5_ff2 0.35fF
C74 net3_ff1 net4_ff1 0.15fF
C75 net3_ff2 a_n100_n729# 0.01fF
C76 net2_ff2 1 0.06fF
C77 net5_ff1 net3_ff1 0.08fF
C78 3 fout 1.06fF
C79 net2_ff2 net5_ff2 0.01fF
C80 finb net4_ff1 0.06fF
C81 3 modi 0.74fF
C82 finb net5_ff1 0.05fF
C83 net3_ff1 VDD 1.29fF
C84 fout P 0.09fF
C85 1 fin 1.54fF
C86 net1_nand3 net2_nand3 0.97fF
C87 modo fout 0.51fF
C88 2 1 0.44fF
C89 VDD 31 2.52fF
C90 modo modi 0.06fF
C91 finb VDD 2.32fF
C92 net3_ff1 net1_ff2 0.06fF
C93 3 net3_ff1 0.05fF
C94 net3_ff2 1 0.50fF
C95 31 net1_ff2 0.01fF
C96 net3_ff2 net5_ff2 0.08fF
C97 3 31 1.51fF
C98 finb net1_ff2 0.01fF
C99 finb 3 0.79fF
C100 fout fin 2.86fF
C101 2 fout 0.84fF
C102 modo net3_ff1 0.10fF
C103 fin modi 0.12fF
C104 modo 31 1.43fF
C105 finb P 0.04fF
C106 finb modo 0.74fF
C107 net3_ff2 fout 0.16fF
C108 net2_ff2 net3_ff1 0.03fF
C109 VDD net4_ff2 0.99fF
C110 net1_ff1 net4_ff1 0.02fF
C111 net3_ff2 modi 0.05fF
C112 net2_ff2 31 0.01fF
C113 3 net2 0.11fF
C114 net2_ff1 net5_ff1 0.01fF
C115 finb net2_ff2 0.01fF
C116 net1_ff2 net4_ff2 0.02fF
C117 net3_ff1 fin 0.88fF
C118 2 net3_ff1 0.02fF
C119 1 a_n100_n729# 0.01fF
C120 net1_nand3 fout 0.12fF
C121 a_n3136_n729# VDD 0.03fF
C122 3 net4_ff2 0.06fF
C123 fin 31 0.17fF
C124 VDD net1_ff1 0.91fF
C125 modo net2 0.04fF
C126 finb fin 2.10fF
C127 net1 modo 0.08fF
C128 finb 2 0.20fF
C129 net3_ff2 net3_ff1 0.09fF
C130 modo net4_ff2 0.64fF
C131 net3_ff2 31 0.19fF
C132 finb net3_ff2 0.44fF
C133 net2_nand3 fout 0.13fF
C134 VDD net4_ff1 1.01fF
C135 1 net5_ff2 0.03fF
C136 net1 fin 0.05fF
C137 net2_ff1 modo 0.02fF
C138 net1 2 0.13fF
C139 finb net1_nand3 0.04fF
C140 fin net4_ff2 0.04fF
C141 net4_ff1 net1_ff2 0.02fF
C142 net3_ff2 net2 0.06fF
C143 net3_ff1 a_n100_n729# 0.01fF
C144 1 fout 0.41fF
C145 net3_ff2 net4_ff2 0.15fF
C146 2 a_n3136_n729# 0.01fF
C147 VDD net1_ff2 1.02fF
C148 fin net1_ff1 0.03fF
C149 3 VDD 1.67fF
C150 net2_ff1 fin 0.06fF
C151 finb net2_nand3 0.05fF
C152 net1 net1_nand3 0.02fF
C153 net5_ff1 modo 0.02fF
C154 3 net1_ff2 0.02fF
C155 VDD P 0.27fF
C156 net5_ff1 net2_ff2 0.01fF
C157 modo VDD 0.90fF
.ends

