** Test bench for BGR

.include ../spice_files/divider.ckt

{{ corner_setup }}

xdiv vdd fout gnd p2 p7 p1 p6 p5 p4 p3 p0 fin float divider

C1 fout GND 25f m=1
I0 opennet GND 0
V5 p5 GND 0
V6 p6 GND 0
V7 p7 GND 0
**** begin user architecture code

.control
    set wr_singlescale
    set wr_vecnames
    set appendwrite
    tran 0.01n 5u
   
    print all

.endc
.measure tran tdiff TRIG v(fout) VAL=0.9 RISE=30 TARG v(fout) VAL=0.9 RISE=31
.measure tran frequency param = {1/tdiff}

.GLOBAL GND
.GLOBAL VDD
.end
*.end