* Extracted by KLayout with SKY130 LVS runset on : 16/11/2022 16:34

.SUBCKT DIVIDER modi5 modi4 modi3 modi6 fout6 fout fout5 fout4 modi P7 P6 P5 P4
+ fout3 VDD fout0 modo fout1 modi0 fout2 modi1 modi2 P0 P1 P2 P3 fin GND
M$1 \$124 fout5 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$2 \$126 fout4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$3 modi5 fout5 \$153 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$4 \$153 \$6 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$5 \$6 \$124 \$156 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$6 \$156 \$45 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$7 \$8 fout5 \$195 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$8 \$195 \$11 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$9 \$11 \$124 \$161 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$10 \$161 fout6 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$11 \$150 fout3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$12 \$149 fout6 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$13 modi4 fout4 \$164 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$14 \$164 \$18 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$15 \$18 \$126 \$167 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$16 \$167 \$58 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$17 \$21 fout4 \$170 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$18 \$170 \$25 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$19 \$25 \$126 \$173 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$20 \$173 fout5 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$21 modi3 fout3 \$205 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$22 \$205 \$30 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$23 \$30 \$150 \$175 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$24 \$175 \$66 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$25 \$31 fout3 \$176 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$26 \$176 \$32 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$27 \$32 \$150 \$212 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$28 \$212 fout4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$29 modi6 fout6 \$180 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$30 \$180 \$36 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$31 \$36 \$149 \$183 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$32 \$183 \$80 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$33 \$2 fout6 \$186 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$34 \$186 \$41 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$35 \$41 \$149 \$189 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$36 \$189 fout VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$37 \$45 \$49 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$38 VDD fout6 \$49 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$39 VDD modi6 \$49 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$40 VDD \$8 fout6 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$41 VDD \$96 fout6 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$42 VDD modi5 \$96 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$43 VDD fout5 \$96 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$44 VDD P6 \$96 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$45 \$58 \$61 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$46 VDD fout5 \$61 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$47 VDD modi5 \$61 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$48 VDD \$21 fout5 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$49 VDD \$65 fout5 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$50 VDD modi4 \$65 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$51 VDD fout4 \$65 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$52 VDD P5 \$65 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$53 \$66 \$69 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$54 VDD modi3 \$79 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$55 VDD fout3 \$79 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$56 VDD P4 \$79 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$57 \$329 P0 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$58 \$80 \$84 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$59 \$329 fin VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$60 VDD fout \$84 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$61 \$329 modo VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$62 VDD modi \$84 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$63 fout0 \$329 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$64 fout0 \$255 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$65 VDD fin \$276 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$66 VDD fout0 \$249 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$67 \$249 \$276 \$251 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$68 VDD \$251 \$253 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$69 \$253 fin \$255 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$70 VDD \$331 \$330 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$71 \$330 \$276 \$258 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$72 VDD \$258 \$260 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$73 \$260 fin modo VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$74 VDD \$2 fout VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$75 VDD \$44 fout VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$76 \$264 modi0 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$77 VDD modi6 \$44 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$78 \$264 fout0 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$79 VDD fout6 \$44 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$80 VDD \$264 \$331 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$81 VDD P7 \$44 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$82 \$332 P1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$83 \$332 fout0 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$84 \$332 modi0 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$85 fout1 \$332 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$86 fout1 \$283 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$87 VDD fout1 \$333 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$88 \$333 \$277 \$280 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$89 VDD \$280 \$334 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$90 \$334 fout0 \$283 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$91 VDD \$335 \$285 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$92 \$285 \$277 \$287 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$93 VDD \$287 \$289 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$94 \$289 fout0 modi0 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$95 \$270 modi1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$96 \$270 fout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$97 VDD \$270 \$335 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$98 \$336 P2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$99 \$336 fout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$100 \$336 modi1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$101 fout2 \$336 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$102 fout2 \$337 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$103 \$311 modi2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$104 \$311 fout2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$105 VDD \$311 \$313 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$106 \$339 P3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$107 \$339 fout2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$108 VDD fout4 \$69 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$109 \$339 modi2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$110 VDD modi4 \$69 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$111 fout3 \$339 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$112 fout3 \$319 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$113 VDD \$31 fout4 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$114 VDD \$79 fout4 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P AD=1.16P
+ PS=8.58U PD=8.58U
M$115 \$343 modi3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$116 \$343 fout3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$117 VDD \$343 \$328 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$118 VDD fout0 \$277 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$119 VDD fout1 \$295 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$120 VDD fout2 \$297 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$121 \$297 \$295 \$299 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$122 VDD \$299 \$301 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$123 \$301 fout1 \$337 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$124 VDD \$313 \$338 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$125 \$338 \$295 \$305 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$126 VDD \$305 \$307 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$127 \$307 fout1 modi1 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$128 VDD fout2 \$314 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$129 VDD fout3 \$340 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$130 \$340 \$314 \$341 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$131 VDD \$341 \$342 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$132 \$342 fout2 \$319 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$133 VDD \$328 \$321 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$134 \$321 \$314 \$323 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$135 VDD \$323 \$325 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$136 \$325 fout2 modi2 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U AS=1.16P
+ AD=1.16P PS=8.58U PD=8.58U
M$137 \$51 \$45 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$138 \$20 \$58 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$139 \$86 \$80 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$140 \$103 \$66 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$141 modi5 \$124 \$50 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$142 \$50 \$6 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$143 \$6 fout5 \$51 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$144 \$8 \$124 \$52 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$145 \$52 \$11 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$146 \$11 fout5 \$53 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$147 \$53 fout6 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$148 modi4 \$126 \$16 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$149 \$16 \$18 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$150 \$18 fout4 \$20 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$151 \$21 \$126 \$23 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$152 \$23 \$25 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$153 \$25 fout4 \$27 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$154 \$27 fout5 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$155 modi3 \$150 \$102 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$156 \$102 \$30 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$157 \$30 fout3 \$103 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$158 \$31 \$150 \$104 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$159 \$104 \$32 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$160 \$32 fout3 \$105 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$161 \$105 fout4 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$162 modi6 \$149 \$85 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$163 \$85 \$36 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$164 \$36 fout6 \$86 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$165 \$2 \$149 \$39 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$166 \$39 \$41 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$167 \$41 fout6 \$87 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$168 \$87 fout GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$169 GND fout6 \$149 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$170 GND fout6 \$47 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$171 \$47 modi6 \$49 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$172 GND fout5 \$124 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$173 GND \$8 \$55 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$174 \$55 \$96 fout6 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$175 GND modi5 \$94 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$176 \$94 fout5 \$95 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$177 \$95 P6 \$96 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$178 GND fout5 \$97 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$179 \$97 modi5 \$61 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$180 GND fout4 \$126 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$181 GND \$21 \$63 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$182 \$63 \$65 fout5 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$183 GND modi4 \$99 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$184 \$99 fout4 \$100 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$185 \$100 P5 \$65 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$186 GND fout3 \$150 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$187 GND modi3 \$108 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$188 \$108 fout3 \$109 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$189 \$109 P4 \$79 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$190 \$329 P0 \$383 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$191 GND \$84 \$80 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$192 \$383 fin \$384 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$193 GND fout \$82 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$194 \$384 modo GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$195 \$82 modi \$84 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$196 fout0 \$329 \$378 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$197 \$378 \$255 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$198 \$276 fin GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$199 GND fout0 \$411 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$200 \$411 fin \$251 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$201 GND \$251 \$414 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$202 \$414 \$276 \$255 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$203 \$420 fin \$258 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$204 GND \$258 \$418 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$205 \$418 \$276 modo GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$206 GND \$2 \$89 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$207 \$89 \$44 fout GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$208 \$264 modi0 \$385 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$209 GND modi6 \$92 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$210 \$385 fout0 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$211 \$92 fout6 \$93 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$212 \$331 \$264 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$213 \$93 P7 \$44 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$214 GND \$49 \$45 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$215 \$332 P1 \$386 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$216 \$386 fout0 \$387 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$217 \$387 modi0 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$218 fout1 \$332 \$389 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$219 \$389 \$283 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$220 \$270 modi1 \$392 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$221 \$392 fout1 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$222 \$335 \$270 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$223 GND \$61 \$58 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$224 \$336 P2 \$405 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$225 \$405 fout1 \$406 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$226 \$406 modi1 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$227 fout2 \$336 \$407 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$228 \$407 \$337 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$229 \$311 modi2 \$397 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$230 \$397 fout2 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$231 \$313 \$311 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$232 \$339 P3 \$408 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$233 GND \$69 \$66 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P AD=0.58P
+ PS=4.58U PD=4.58U
M$234 \$408 fout2 \$409 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$235 GND fout4 \$101 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$236 \$409 modi2 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$237 \$101 modi4 \$69 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$238 fout3 \$339 \$400 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$239 \$400 \$319 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$240 GND \$31 \$106 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P AD=1.74P
+ PS=12.58U PD=12.58U
M$241 \$106 \$79 fout4 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$242 \$343 modi3 \$403 GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$243 \$403 fout3 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=6U AS=1.74P
+ AD=1.74P PS=12.58U PD=12.58U
M$244 \$328 \$343 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$245 GND \$331 \$420 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$246 \$277 fout0 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$247 GND fout1 \$422 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$248 \$422 fout0 \$280 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$249 GND \$280 \$425 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$250 \$425 \$277 \$283 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$251 GND \$335 \$427 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$252 \$427 fout0 \$287 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$253 GND \$287 \$430 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$254 \$430 \$277 modi0 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$255 \$295 fout1 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$256 GND fout2 \$433 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$257 \$433 fout1 \$299 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$258 GND \$299 \$436 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$259 \$436 \$295 \$337 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$260 GND \$313 \$438 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$261 \$438 fout1 \$305 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$262 GND \$305 \$441 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$263 \$441 \$295 modi1 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$264 \$314 fout2 GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$265 GND fout3 \$444 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$266 \$444 fout2 \$341 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$267 GND \$341 \$447 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$268 \$447 \$314 \$319 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$269 GND \$328 \$449 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$270 \$449 fout2 \$323 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$271 GND \$323 \$452 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
M$272 \$452 \$314 modi2 GND sky130_fd_pr__nfet_01v8 L=0.15U W=2U AS=0.58P
+ AD=0.58P PS=4.58U PD=4.58U
.ENDS DIVIDER
