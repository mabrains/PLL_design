** Test bench for BGR
.include {{ current_path }}/../../../circuit/bgr_pex.ext
.include {{ current_path }}/../../../circuit/bgr_sch.ckt
.include {{ current_path }}/../../../circuit/vco_load.ckt

{{ corner_setup }}


** xbgr_pex out GND VDD bgr_pex
xbgr_sch out GND VDD bgr_sch
xvco_load out vco_load

.control
    set wr_singlescale
    set wr_vecnames
    set appendwrite

    op
    **const load**
    *let Iref = i(VTuner)*1000000

    **variant load**
    let Iref  = @m.xvco_load.xm8.msky130_fd_pr__nfet_01v8[id]*1000000
    print Iref
    print all

   
    
.endc

.GLOBAL GND
.GLOBAL VDD
.end