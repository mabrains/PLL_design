** sch_path: /home/ahmed/Mabrains_internship/VCO_Try3/VCO_Full_2.sch
**.subckt VCO_Full_2
*VDD VDD GND 1.8 
VDD VDD GND V_supply



XM11 vp vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=50 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
XM1 vn vp net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=50 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
XM2 vp vn GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
L1 vp net4 4n m=1
R1 vp vn 1182 m=1
R2 net4 vn 3 m=1
XM7 vn vp GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
C1 vp vn 5f m=10
C3 vp GND 5f m=5
C2 vn GND 5f m=5
VTuner net5 GND 1.5
C13 vp vn 10f m=15

* Varactor 
*******************old******************
XM6 net5 vn net5 gnd sky130_fd_pr__nfet_01v8_lvt L=0.6 W=17 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20
XM3 net5 vp net5 gnd sky130_fd_pr__nfet_01v8_lvt L=0.6 W=17 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20


*********************new******************
*XM6 net5 vn net5 net5 sky130_fd_pr__nfet_01v8_lvt L=2.7 W=49.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
*+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
*+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
*
*XM3 net5 vp net5 net5 sky130_fd_pr__nfet_01v8_lvt L=2.7 W=49.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
*+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
*+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2

*********************************************
XM4 net3 net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=50 m=50
XM5 net1 net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10

Isource net1 GND 450u
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /open_design_environment/foundry/pdks/skywaters/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /open_design_environment/foundry/pdks/skywaters/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice

*corners setup
.temp 27
.options tnom=27
.param V_supply = 1.8
.include /open_design_environment/foundry/pdks/skywaters/sky130A/libs.tech/ngspice/corners/tt.spice
.include /open_design_environment/foundry/pdks/skywaters/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


.save all
.nodeset v(vout)=0
.control

compose  vctrl_vector   start=0         stop=1.8          step=0.1
let vctrl_counter = 0
let f_osc = vector(length(vctrl_vector))
let curr_value = vctrl_vector[0]
set appendwrite
while vctrl_counter < length(vctrl_vector)
    print curr_value
    alter VTuner  $&curr_value
    op
    save  @m.xm4.msky130_fd_pr__pfet_01v8[id]

    save  @m.xm1.msky130_fd_pr__pfet_01v8[id]
    save  @m.xm11.msky130_fd_pr__pfet_01v8[id]

    save  @m.xm7.msky130_fd_pr__nfet_01v8[id]
    save  @m.xm2.msky130_fd_pr__nfet_01v8[id]

    save  vp
    save  vn

    wrdata csv_files/I_tail_tttt.csv   @m.xm4.msky130_fd_pr__pfet_01v8[id]
    wrdata csv_files/Ip_left_tttt.csv  @m.xm1.msky130_fd_pr__pfet_01v8[id]
    wrdata csv_files/Ip_right_tttt.csv @m.xm11.msky130_fd_pr__pfet_01v8[id]
    wrdata csv_files/In_left_tttt.csv  @m.xm7.msky130_fd_pr__nfet_01v8[id]
    wrdata csv_files/In_right_tttt.csv @m.xm2.msky130_fd_pr__nfet_01v8[id]
    wrdata csv_files/vp_tttt.csv vp
    wrdata csv_files/vn_tttt.csv vn

    tran 0.01ns 100ns
    let vdiff = v(vp)-v(vn)
    let vdiff_max =  vecmax(vp-vn)
    meas tran tperiod TRIG vdiff VAL=0.4 RISE=30 TARG vdiff VAL=0.4 RISE=31
    let freq = 1/tperiod
    setplot op
    let f_osc[vctrl_counter] = tran.freq

    wrdata csv_files/fosc_vs_vctrl_tttt.csv f_osc[vctrl_counter]
    wrdata csv_files/max_swing_tttt.csv tran.vdiff_max
    wrdata csv_files/time_swing_tttt.csv tran.vdiff

    reset
    let vctrl_counter = vctrl_counter + 1
    let curr_value = vctrl_vector[vctrl_counter]
end

let kvco = vecd(f_osc)
print f_osc
*plot f_osc vs vctrl_vector
*plot kvco vs vctrl_vector xlimit 0.5 1.6
*print kvco
quit
.endc


**** end user architecture code
**.ends

* expanding   symbol:  BGR_Banba.sym # of pins=3
** sym_path: /home/ahmed/Mabrains_internship/VCO_Try3/BGR_Banba.sym
** sch_path: /home/ahmed/Mabrains_internship/VCO_Try3/BGR_Banba.sch

.GLOBAL GND
.GLOBAL VDD
.end
