****************

.subckt BGR  Iref GND VDD VBE net1 net2 net3 net4 net6 
Q1 GND GND VBE GND sky130_fd_pr__pnp_05v5_W0p68L0p68 NE=1 m=1
Q2 GND GND net2 GND sky130_fd_pr__pnp_05v5_W0p68L0p68 NE=8


R4 net2 net3 GND sky130_fd_pr__res_xhigh_po_1p41 L=20.24u mult=1 m=1
R1 GND net3 GND sky130_fd_pr__res_xhigh_po_1p41 L=70u mult=1 m=1
R3 GND VBE GND sky130_fd_pr__res_xhigh_po_1p41 L=70u mult=1 m=1

Rd1 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 L=10.12u W=5.64umult=1 m=1

M15 net5 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5u W=4u nf=4    
M13 net3 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5u W=20u nf=4    
M14 VBE net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5u W=20u nf=4  
M16 net1 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=44u nf=44
M17 net6 net3 net5 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5u W=90u nf=6      
M18 net4 VBE net5 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5u W=90u nf=6            
M19 net1 net6 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5u W=0.42u m=10      
M20 net6 net4 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5u W=0.42u m=4             
M21 net4 net4 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5u W=0.42u m=4             
M22 net7 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1u W=40u nf=2     
M23 net7 net1 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=20u W=0.42u         
M24 VBE net7 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1u W=40u nf=2     
M2 Iref net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5u W=200u nf=40    
  
.ends
