** sch_path: /home/ahmed/PLL_Internship/transient_noise.sch
**.subckt transient_noise

.csparam W = 60
.csparam L = 0.15
.csparam R = 1e3 

XM1 net2 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=60 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1

VDD VDD GND 1.8
R1 VDD vout 1k m=1
Vsource vin GND DC 0.8 SIN (0.8 1m 1e9)

VmosNoise net1 vin DC 0 trnoise ( 0 0 0 0)
VresNoise vout net2 DC 0 trnoise (0 0 0 0)
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
**** begin user architecture code


.tran 0.05n 5000n

.control
*==============================DC SIMULATION===================================================================
  op
  let gm = @m.xm1.msky130_fd_pr__nfet_01v8[gm]
  save  @m.xm1.msky130_fd_pr__nfet_01v8[vds]
  save  @m.xm1.msky130_fd_pr__nfet_01v8[id]
  save  @m.xm1.msky130_fd_pr__nfet_01v8[gm]
  save  @m.xm1.msky130_fd_pr__nfet_01v8[vth]
  save gm
  save vin
  save vout
  save net1
  save net2
  
  echo ******************************************************************************************************
  echo DC Peremeters
  print  @m.xm1.msky130_fd_pr__nfet_01v8[vds]
  print  @m.xm1.msky130_fd_pr__nfet_01v8[id]
  print  @m.xm1.msky130_fd_pr__nfet_01v8[gm]
  print  @m.xm1.msky130_fd_pr__nfet_01v8[vds]-@m.xm1.msky130_fd_pr__nfet_01v8[vgs]+@m.xm1.msky130_fd_pr__nfet_01v8[vth]
  print vin
  print vout
  print v(net1)
  print v(net2)
  print gm
  echo ******************************************************************************************************
  set color0=white
  set color1=black
*==============================TRANSIENT SIMULATION WITHOUT NOISE=============================================
  alter @VmosNoise[trnoise] = 0 0 0 0 
  alter @VresNoise[trnoise] = 0 0 0 0 
  run
  save @m.xm1.msky130_fd_pr__nfet_01v8[gm]
  let gm_no_noise = @m.xm1.msky130_fd_pr__nfet_01v8[gm]
  save gm_no_noise
  *plot gm_no_noise
  
  plot vout xlimit 30n 50n
  linearize
  fft vout
  *spec 0.5 1.5e9 210e3 vout
  
  
*==============================CALCULATE RMS VALUES===========================================================
*=======CONSTANTS==========================
  let eps_o      = 8.854187817*1e-12
  let eps_r      = 12
  let t_ox       = 0.07*1e-6
  let k_flkr_mos = 10^-25
  let k          = 1.38*1e-23
  let temp       = 300
*========EQUATIONS=========================
  let cox        = eps_o*eps_r/t_ox
  let fc_flkr    = (3*tran1.gm_no_noise*k_flkr_mos)/(8*cox*k*temp*W*L)
  
  let v_flkr_mos = sqrt((k_flkr_mos)/(fc_flkr*cox*W*L))
  let v_whit_mos = sqrt((8*k*temp)/(3*tran1.gm_no_noise))
  let v_whit_res = sqrt(4*k*temp*R)
  
  print eps_o eps_r t_ox k_flkr_mos k temp cox length(fc_flkr) length(v_flkr_mos) v_whit_res 
  wrdata gm_no_noise.csv tran1.gm_no_noise
  
.endc

**** end user architecture code
.end
