* PLL subckt

.INCLUDE ../../BGR/circuit/bgr_cir.ckt
.INCLUDE ../../XCTL/behav/xctl_behave.ckt
.INCLUDE ../../CP/circuit/cp_cir.ckt
.INCLUDE ../../PFD/circuit/pfd_cir.ckt
.INCLUDE ../../LPF/circuit/lf_cir.ckt
.include ../../VCO/circuit/vco_cir.ckt
.include ../../VCO/circuit/inductor_model_cct.ckt
.include ../../Divider/circuit/div_cir.ckt


.param p0_val = {0}
.param p1_val=  {0}
.param p2_val=  {0}
.param p3_val=  {0}
.param p4_val=  {1}
.param p5_val=  {0}
.param p6_val=  {0}
.param p7_val=  {0}


.subckt pll_cir REF FB UP DWN iout vctrl vco_out VDD GND

Xctl_behave REF VDD GND xctl_behave

Xconventional_pfd  REF VDD GND FB UP DN conventional_pfd

Xcp  UP VOP DN VDD GND CP_with_buffer 

Vtest VOP ilf DC 0

Xloop_filter_3rd_order ilf vctrl GND loop_filter_3rd_order 

xvco vp vn vctrl ibias VDD GND vco_cir
* xinv_vco1 vdd vp vp2 gnd
* xinv_vco2 vdd vn vn2 gnd
xind1 vp vn ind_model
** xbgr ibias GND VDD BGR_Banba
Isource VDD ibias 90u          $ original
xdiv VDD FB GND p2 p7 p1 p6 p5 p4 p3 p0 vp opennet1 divider
xdivdumyy VDD fdummy GND p2 p7 p1 p6 p5 p4 p3 p0 vn opennet divider


.ic v(vctrl)=0

VP1 p2 GND {p2_val}
VP2 p4 GND {p4_val}
VP3 p1 GND {p1_val}
VP4 p3 GND {p3_val}
VP5 p5 GND {p5_val}
VP6 p6 GND {p6_val}
VP7 p0 GND {p0_val}
VP8 p7 GND {p7_val}

.ends