** sch_path: /home/ahmed/PLL_Internship/transient_noise.sch
**.subckt transient_noise

.csparam W = 60
.csparam L = 0.15
.csparam R = 1e3 

XM1 net2 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=60 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1

VDD VDD GND 1.8
R1 VDD vout 1k m=1
Vsource vin GND DC 0.8 SIN (0.8 1m 1e9)


**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
**** begin user architecture code


.tran 0.1n 500n

.control
*==============================DC SIMULATION===================================================================
  op
  let gm = @m.xm1.msky130_fd_pr__nfet_01v8[gm]
  save  @m.xm1.msky130_fd_pr__nfet_01v8[vds]
  save  @m.xm1.msky130_fd_pr__nfet_01v8[id]
  save  @m.xm1.msky130_fd_pr__nfet_01v8[gm]
  save  @m.xm1.msky130_fd_pr__nfet_01v8[vth]
  save vin
  save vout
  save net1
  save net2
  echo ******************************************************************************************************
  echo DC Peremeters
  print  @m.xm1.msky130_fd_pr__nfet_01v8[vds]
  print  @m.xm1.msky130_fd_pr__nfet_01v8[id]
  print  @m.xm1.msky130_fd_pr__nfet_01v8[gm]
  print  @m.xm1.msky130_fd_pr__nfet_01v8[vds]-@m.xm1.msky130_fd_pr__nfet_01v8[vgs]+@m.xm1.msky130_fd_pr__nfet_01v8[vth]
  print vin
  print vout
  print v(net1)
  print v(net2)
  echo ******************************************************************************************************
  set color0=white
  set color1=black
*==============================TRANSIENT SIMULATION WITH NOISE================================================
  run
  *plot vin xlimit 30n 50n
  linearize vin
  fft vin 

  setplot tran1
  *plot v(net1) xlimit 30n 50n
  linearize v(net1)
  fft v(net1)

  setplot tran1
  *plot vout xlimit 30n 50n
  linearize vout
  fft vout
  
  *plot mag(sp2.vout) mag(sp4.vin) mag(sp5.v(net1)) mag(sp6.vout) xlimit 0.9G 1.1G ylimit 0.1 1e-11 ylog
  *plot mag(sp2.vout)  mag(sp6.vout) xlimit 0.9G 1.1G ylimit 0.1 1e-11 ylog
  
  plot mag(sp2.vin) mag(sp4.vout) xlimit 0.9G 1.1G ylimit 3 1e-10 ylog
  wrdata vout_fft.csv mag(sp4.vout)
  
*==============================PHASE NOISE CALCULATION================================================
.endc

**** end user architecture code
.end
