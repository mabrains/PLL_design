** Test bench for VCO

.include ../circuit/inv.ckt
.include ../circuit/vco_sch.ckt
.include ../../BGR/circuit/bgr_sch.ckt 
.include ../circuit/inductor_model_cct.ckt



.lib /open_design_environment/foundry/pdks/skywaters/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.temp 27
.options tnom=27

VDD VDD GND 1.8
VTuner vctrl GND 0.5

xinv   vp  vp2 VDD GND inv
xinv2  vp2 vp3 VDD GND inv

xinv3 vn  vn2 VDD GND inv
xinv4 vn2 vn3 VDD GND inv

Vpulse vin GND PULSE(0 1.8 1ns 1ns 1ns 4ns 10ns)
xvco vp vn vctrl ibias VDD GND vco_sch
xind1 vp vn ind_model
XC_load vp vn sky130_fd_pr__cap_mim_m3_1 W=15 L=9 MF=1 m=1  $mim cap
xbgr ibias GND VDD bgr_sch
** Isource VDD ibias 90u

.control
    set appendwrite 
    op
    save all
    print all
    tran 0.01ns 200ns
    plot vp vp3
    plot vn vn3
    ** meas tran inv_delay  trig v(vin)  val=0.9  fall=10 targ v(vout) val=0.9   rise=10

    ** let inv_delay2 =  inv_delay*1G*1000
    ** print inv_delay2

    *quit

    let vdiff = v(vp)-v(vn)
    let vdiff_max =  vecmax(vp-vn)
    print vdiff_max
    meas tran tperiod TRIG vdiff VAL=0.4 RISE=30 TARG vdiff VAL=0.4 RISE=31
    let freq = 1/(tperiod*1000000000)
    print freq

    let vdiff2 = v(vp2)-v(vn2)
    let vdiff_max2 =  vecmax(vp2-vn2)
    print vdiff_max2
    meas tran tperiod2 TRIG vdiff2 VAL=0.4 RISE=30 TARG vdiff2 VAL=0.4 RISE=31
    let freq2 = 1/(tperiod2*1000000000)
    print freq2

    let vdiff3 = v(vp3)-v(vn3)
    let vdiff_max3 =  vecmax(vp3-vn3)
    print vdiff_max3
    meas tran tperiod3 TRIG vdiff3 VAL=0.4 RISE=30 TARG vdiff3 VAL=0.4 RISE=31
    let freq3 = 1/(tperiod3*1000000000)
    print freq3
    
    
    

.endc

.GLOBAL GND
.GLOBAL VDD
.end