*********************************************************
*******************charge pump cdl file****************** 
*********************************************************
.subckt CP VDD GND UP DN VOP ibias_cp 

***************non ideal current source*****************
M_cp_p1 ibias_cp ibias_cp VDD VDD sky130_fd_pr__pfet_01v8 L=0.15u W=40u nf=4 m=1
M_cp_p2 VBN      ibias_cp VDD VDD sky130_fd_pr__pfet_01v8 L=0.15u W=10u nf=1 m=1


M_cp_1 cp_net1 Nbais GND GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U nf=1 m=2
M_cp_2 cp_net2 Nbais GND GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U nf=1 m=1
M_cp_3 VBp VBN cp_net1 GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U nf=1 m=2
M_cp_4 Nbais VBN cp_net2 GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U nf=1 m=1

R_cp1 VBN Nbais VDD sky130_fd_pr__res_iso_pw r=23.0188679245k   m=1 L=60u  W=7.95u
R_cp2 p_bais VBp VDD sky130_fd_pr__res_iso_pw r=11.5094339623k  m=1 L=30u  W=7.95u  
Rdumy VDD VDD VDD sky130_fd_pr__res_iso_pw r=17.2641509434k     m=1 L=30u  W=5.3u  

M_cp_5 p_bais VBp cp_net3 VDD sky130_fd_pr__pfet_01v8 L=0.6U W=6.66U nf=1 m=2
M_cp_6 cp_net3 p_bais VDD VDD sky130_fd_pr__pfet_01v8 L=0.6U W=6.66U nf=1 m=2

M_cp_7 cp_net4 Nbais GND GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U nf=1 m=10
M_cp_8 cp_net5 VBN cp_net4 GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U nf=1 m=10
M_cp_9 VON DNB cp_net5 GND sky130_fd_pr__nfet_01v8 L=0.15U W=4U nf=1 m=1
M_cp_10 VOP DN cp_net5 GND sky130_fd_pr__nfet_01v8 L=0.15U W=4U nf=1 m=1
M_cp_11 VOP UBP cp_net6 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=10U nf=1 m=1
M_cp_12 VON UP cp_net6 VDD sky130_fd_pr__pfet_01v8 L=0.15U W=10U nf=1 m=1
M_cp_13 cp_net6 VBp cp_net7 VDD sky130_fd_pr__pfet_01v8 L=0.6U W=6.66U nf=1 m=10
M_cp_14 cp_net7 p_bais VDD VDD sky130_fd_pr__pfet_01v8 L=0.6U W=6.66U nf=1 m=10

M_cp_15 UBP UP GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_16 UBP UP VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=2U nf=1 m=1

M_cp_17 DNB DN GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_18 DNB DN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15U W=2U nf=1 m=1

M_cp_19 cp_net2_ota Nbais GND GND sky130_fd_pr__nfet_01v8 L=0.6U W=2U nf=1 m=2
M_cp_20 cp_net1_ota p_bais VDD VDD sky130_fd_pr__pfet_01v8 L=0.6U W=4U nf=1 m=2
M_cp_21 cp_net3_ota p_bais VDD VDD sky130_fd_pr__pfet_01v8 L=0.6U W=4U nf=1 m=2
M_cp_22 cp_net3_ota VON cp_net2_ota GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_23 cp_net1_ota VOP cp_net2_ota GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_24 cp_net5_ota cp_net4_ota GND GND sky130_fd_pr__nfet_01v8 L=1U W=1.3U nf=1 m=1
M_cp_25 GND cp_net4_ota GND GND sky130_fd_pr__nfet_01v8 L=1U W=1.3U nf=1 m=1
M_cp_26 cp_net4_ota VBN cp_net5_ota GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_27 VON VBN GND GND sky130_fd_pr__nfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_28 VON VBp cp_net3_ota VDD sky130_fd_pr__pfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_29 cp_net4_ota VBp cp_net1_ota VDD sky130_fd_pr__pfet_01v8 L=0.15U W=1U nf=1 m=1
M_cp_30 cp_net6_ota p_bais VDD VDD sky130_fd_pr__pfet_01v8 L=0.6U W=6.66U nf=1 m=1
M_cp_32 GND VON cp_net6_ota VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1
M_cp_33 cp_net5_ota VOP cp_net6_ota VDD sky130_fd_pr__pfet_01v8 L=0.15U W=4U nf=1 m=1


.ends