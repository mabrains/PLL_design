** sch_path: /home/ahmed/PLL_Internship/Ahmed Elshahat LC VCO/CMOS_LC_VCO/CMOS_VCO/varactor.sch
**.subckt varactor
.param len = 1
.param width = 90.2
.param mul = 2
.param fingNum = 1
XM1 v_tunN v_tunP v_tunN v_tunN sky130_fd_pr__nfet_01v8 L=len W=width nf=fingNum ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=mul


XM2 v_tunN v_tunP v_tunN v_tunN sky130_fd_pr__pfet_01v8 L=len W=width nf=fingNum ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=mul

XM3 v_tunN v_tunP v_tunN GND sky130_fd_pr__nfet_01v8 L=len W=width nf=fingNum ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=mul

XM4 v_tunN v_tunP v_tunN VDD sky130_fd_pr__pfet_01v8 L=len W=width nf=fingNum ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=mul

VDD VDD GND 1.8
V_tun v_tunN GND dc=0
V_tank v_tunP GND 1.3
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD

.control
let v_min  = 0
let v_step = 0.01
let v_max  = 2.5

save @m.xm1.msky130_fd_pr__nfet_01v8[cgg] 
save @m.xm1.msky130_fd_pr__nfet_01v8[cgs] 
save @m.xm1.msky130_fd_pr__nfet_01v8[cgd] 
save @m.xm1.msky130_fd_pr__nfet_01v8[cdd] 
save @m.xm1.msky130_fd_pr__nfet_01v8[cdb] 
save @m.xm1.msky130_fd_pr__nfet_01v8[cgb] 
save @m.xm1.msky130_fd_pr__nfet_01v8[csb]

save @m.xm2.msky130_fd_pr__pfet_01v8[cgg] 
save @m.xm2.msky130_fd_pr__pfet_01v8[cgs] 
save @m.xm2.msky130_fd_pr__pfet_01v8[cgd] 
save @m.xm2.msky130_fd_pr__pfet_01v8[cdd] 
save @m.xm2.msky130_fd_pr__pfet_01v8[cdb] 
save @m.xm2.msky130_fd_pr__pfet_01v8[cgb] 
save @m.xm2.msky130_fd_pr__pfet_01v8[csb]

save @m.xm3.msky130_fd_pr__nfet_01v8[cgg] 
save @m.xm3.msky130_fd_pr__nfet_01v8[cgs] 
save @m.xm3.msky130_fd_pr__nfet_01v8[cgd] 
save @m.xm3.msky130_fd_pr__nfet_01v8[cdd] 
save @m.xm3.msky130_fd_pr__nfet_01v8[cdb] 
save @m.xm3.msky130_fd_pr__nfet_01v8[cgb] 
save @m.xm3.msky130_fd_pr__nfet_01v8[csb]

save @m.xm4.msky130_fd_pr__pfet_01v8[cgg] 
save @m.xm4.msky130_fd_pr__pfet_01v8[cgs] 
save @m.xm4.msky130_fd_pr__pfet_01v8[cgd] 
save @m.xm4.msky130_fd_pr__pfet_01v8[cdd] 
save @m.xm4.msky130_fd_pr__pfet_01v8[cdb] 
save @m.xm4.msky130_fd_pr__pfet_01v8[cgb] 
save @m.xm4.msky130_fd_pr__pfet_01v8[csb]

DC V_tun $&v_min $&v_max $&v_step

let cgg1 = @m.xm1.msky130_fd_pr__nfet_01v8[cgg] 
let cgg2 = @m.xm2.msky130_fd_pr__pfet_01v8[cgg] 
let cgg3 = @m.xm3.msky130_fd_pr__nfet_01v8[cgg]
let cgg4 = @m.xm4.msky130_fd_pr__pfet_01v8[cgg] 

let cgs1 = @m.xm1.msky130_fd_pr__nfet_01v8[cgs] 
let cgs2 = @m.xm2.msky130_fd_pr__pfet_01v8[cgs] 
let cgs3 = @m.xm3.msky130_fd_pr__nfet_01v8[cgs]
let cgs4 = @m.xm4.msky130_fd_pr__pfet_01v8[cgs] 

let cgg1_deriv = deriv(cgg1)
let cgg2_deriv = deriv(cgg2)
let cgg3_deriv = deriv(cgg3)
let cgg4_deriv = deriv(cgg4)

let cgg1_deriv = deriv(cgg1_deriv)
let cgg2_deriv = deriv(cgg2_deriv)
let cgg3_deriv = deriv(cgg3_deriv)
let cgg4_deriv = deriv(cgg4_deriv)

meas dc v1 FIND cgg1 WHEN v-sweep=0.2 CROSS=LAST
meas dc v2 FIND cgg1 WHEN v-sweep=1.2 CROSS=LAST
print v1-v2

plot cgg1 cgg2 cgg3 cgg4 
plot cgs1 cgs2 cgs3 cgs4

*plot cgg1_deriv cgg2_deriv cgg3_deriv cgg4_deriv
*quit
.endc

.end
