**behaviour of the divider