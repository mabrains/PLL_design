** Test bench for ring

.include ../PEX/TOP_PEX.ext

.lib /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.temp 27.00
.options tnom=27.00
VDD VDD GND PWL(0 0 1u 1.8 0.8m 1.8)


xring Vin out VDD GND TOP

**** begin user architecture code

.control

    op 
    save all
        
    print all

    tran 5n 0.8m
    plot out
    meas tran tperiod TRIG out VAL=1.5 RISE=750 TARG out VAL=1.5 RISE=755
    let freq = 5/(tperiod*1000000)
    print freq
    
.endc

.GLOBAL GND
.GLOBAL VDD
.end
