* XCTL subckt

.PARAM main_freq = 10.0Meg
.PARAM cycle     = {1.0/main_freq}
.PARAM tpw       = {cycle / 2}
.PARAM t_rise    = {cycle / 50}
.PARAM t_fall    = {cycle / 50}
.PARAM t_delay   = {0}

.subckt xctl_behave REF VDD GND
+ trise={t_rise}   tfall={t_fall} T_cycle={cycle}
+ pulsewidth={tpw} delay={t_delay}

    Vref REF GND PULSE ( 0 1.8 delay trise t_fall pulsewidth T_cycle 0)

.ends