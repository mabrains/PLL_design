** sch_path: /home/ahmed/Mabrains_internship/VCO_Try1/VCO_try7.sch
**.subckt VCO_try7
XM11 vp net9 net1 net1 sky130_fd_pr__pfet_01v8 L=0.15 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
XM1 vn net8 net1 net1 sky130_fd_pr__pfet_01v8 L=0.15 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
XM2 vp net7 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
L1 vp net14 4n m=1
I0 net2 GND 5m
R1 net12 vn 1182 m=1
VDD VDD GND 1.8
R2 net13 vn 3 m=1
XM4 net1 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
XM5 net2 net5 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
XM7 vn net6 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
C1 vp vn 5f m=10
C3 vp GND 5f m=5
C2 vn GND 5f m=5
Vctrl net4 GND 1.7
XM10 net4 net10 net4 GND sky130_fd_pr__pfet_01v8_lvt L=1.3 W=12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
XM3 net4 net11 net4 GND sky130_fd_pr__pfet_01v8_lvt L=1.3 W=12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
C13 vp vn 10f m=10
V7 net6 vp DC 0 trnoise (0 0 0 0)
V2 net7 vn DC 0 trnoise (0 0 0 0)
V1 net8 vp DC 0 trnoise (0 0 0 0)
V11 net9 vn DC 0 trnoise (0 0 0 0)
V4 net3 net2 DC 0 trnoise (0 0 0 0)
V5 net5 net2 DC 0 trnoise (0 0 0 0)
V10 net10 vn DC 0 trnoise (0 0 0 0)
V3 net11 vp DC 0 trnoise (0 0 0 0)
VR1 net12 vp DC 0 trnoise (0 0 0 0)
VR2 net13 net14 DC 0 trnoise (0 0 0 0)
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


.tran 0.03n 20u
.save all
.control
  op
  save @m.xm1.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm11.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm2.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm4.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm5.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm7.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm10.msky130_fd_pr__pfet_01v8_lvt[gm]
  save @m.xm3.msky130_fd_pr__pfet_01v8_lvt[gm]

  run
  save @m.xm1.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm11.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm2.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm4.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm5.msky130_fd_pr__pfet_01v8[gm]
  save @m.xm7.msky130_fd_pr__nfet_01v8[gm]
  save @m.xm10.msky130_fd_pr__pfet_01v8_lvt[gm]
  save @m.xm3.msky130_fd_pr__pfet_01v8_lvt[gm]

 
  let vdiff = v(vp)-v(vn)
  save vdiff
  *plot vdiff
  linearize vdiff
  *save vdiff
  *fft (v(vp)-v(vn))
  fft vdiff
  *spec 0.5 1.5e9 210e3 vout
  
  
  wrdata gm1_no_noise.csv tran1.@m.xm1.msky130_fd_pr__pfet_01v8[gm]
  wrdata gm11_no_noise.csv tran1.@m.xm11.msky130_fd_pr__pfet_01v8[gm]
  wrdata gm2_no_noise.csv tran1.@m.xm2.msky130_fd_pr__nfet_01v8[gm]
  wrdata gm4_no_noise.csv tran1.@m.xm4.msky130_fd_pr__pfet_01v8[gm]
  wrdata gm5_no_noise.csv tran1.@m.xm5.msky130_fd_pr__pfet_01v8[gm]
  wrdata gm7_no_noise.csv tran1.@m.xm7.msky130_fd_pr__nfet_01v8[gm]
  wrdata gm10_no_noise.csv tran1.@m.xm10.msky130_fd_pr__pfet_01v8_lvt[gm]
  wrdata gm3_no_noise.csv tran1.@m.xm3.msky130_fd_pr__pfet_01v8_lvt[gm]
  

  plot mag(sp2.vdiff)
  
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
