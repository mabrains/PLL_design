* NGSPICE file created from CP.ext - technology: sky130A

.subckt CP UBP UP VBN DN DNB Nbais p_bais VBP net3 net5 net6 VOP net6_ota net5_ota
+ net3_ota net1_ota net1 net2 net4 net7 VON VDD GND
X0 net6.t6 UBP.t2 VOP.t0 VDD.t23 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1 VDD.t44 VDD.t45 VDD sky130_fd_pr__res_iso_pw w=2.65e+06u l=3e+07u
X2 w_4269_n7633# VBN.t1 VDD sky130_fd_pr__res_iso_pw w=2.65e+06u l=3e+07u
X3 VDD.t55 p_bais.t5 net1_ota.t2 VDD.t54 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=600000u
X4 net5.t10 VBN.t3 net4.t8 GND.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X5 VBP.t0 p_bais.t2 VDD sky130_fd_pr__res_iso_pw w=2.65e+06u l=3e+07u
X6 VDD.t57 p_bais.t6 net1_ota.t1 VDD.t56 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=600000u
X7 net3_ota.t3 VBP.t5 VON.t2 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VBP.t3 p_bais.t3 VDD sky130_fd_pr__res_iso_pw w=2.65e+06u l=3e+07u
X9 net4.t0 Nbais.t4 GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X10 DNB.t1 DN.t0 GND.t58 GND.t57 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VBP.t2 VBN.t4 net1.t1 GND.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X12 net4.t17 Nbais.t5 GND.t46 GND.t45 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X13 VDD.t3 VDD.t4 VDD sky130_fd_pr__res_iso_pw w=2.65e+06u l=3e+07u
X14 net5.t9 VBN.t5 net4.t12 GND.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X15 GND.t40 a_48058_n6837.t2 net5_ota.t1 GND.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.3e+06u l=1e+06u
X16 net4.t5 Nbais.t6 GND.t15 GND.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X17 net7.t9 p_bais.t7 VDD.t59 VDD.t58 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X18 VON.t1 DNB.t2 net5.t0 GND.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X19 w_4269_n7633# VBN.t0 VDD sky130_fd_pr__res_iso_pw w=2.65e+06u l=3e+07u
X20 net7.t8 p_bais.t8 VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X21 net5.t8 VBN.t6 net4.t7 GND.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X22 VOP.t1 DN.t1 net5.t11 GND.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X23 net6.t7 VBP.t6 net7.t19 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X24 UBP.t0 UP.t0 VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X25 a_16669_n8264.t1 VOP.t2 net1_ota.t3 GND.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 net4.t2 Nbais.t7 GND.t9 GND.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X27 net6.t8 VBP.t7 net7.t18 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X28 p_bais.t1 VBP.t8 net3.t3 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X29 net5.t7 VBN.t7 net4.t15 GND.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X30 net6_ota.t0 VON.t4 GND.t0 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X31 net4.t4 Nbais.t8 GND.t13 GND.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X32 net6.t0 VBP.t9 net7.t17 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X33 net7.t7 p_bais.t9 VDD.t49 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X34 net5.t6 VBN.t8 net4.t10 GND.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X35 a_16669_n8264.t3 Nbais.t9 GND.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X36 net1.t3 Nbais.t10 GND.t52 GND.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X37 net6.t1 VBP.t10 net7.t16 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X38 p_bais.t0 VBP.t11 net3.t2 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X39 w_4269_n7633# Nbais.t1 VDD sky130_fd_pr__res_iso_pw w=2.65e+06u l=3e+07u
X40 net7.t6 p_bais.t10 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X41 net4.t1 Nbais.t11 GND.t7 GND.t6 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X42 UBP.t1 UP.t1 GND.t21 GND.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 net5.t5 VBN.t9 net4.t13 GND.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X44 net1_ota.t0 VBP.t12 a_48058_n6837.t0 VDD.t27 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 net6_ota.t1 p_bais.t11 VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X46 VDD.t36 p_bais.t12 net3_ota.t2 VDD.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=600000u
X47 net3.t1 p_bais.t13 VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X48 VDD.t40 p_bais.t14 net3_ota.t1 VDD.t39 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=600000u
X49 w_4269_n7633# VBN.t2 VDD sky130_fd_pr__res_iso_pw w=2.65e+06u l=3e+07u
X50 VBP.t1 VBN.t10 net1.t0 GND.t30 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X51 net7.t5 p_bais.t15 VDD.t42 VDD.t41 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X52 Nbais.t0 VBN.t11 net2.t0 GND.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X53 DNB.t0 DN.t2 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X54 net7.t4 p_bais.t16 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X55 GND.t28 VBN.t12 VON.t3 GND.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X56 w_4269_n7633# Nbais.t3 VDD sky130_fd_pr__res_iso_pw w=2.65e+06u l=3e+07u
X57 net5.t4 VBN.t13 net4.t14 GND.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X58 net6.t5 UP.t2 VON.t0 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X59 net7.t3 p_bais.t17 VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X60 net5.t3 VBN.t14 net4.t9 GND.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X61 net7.t2 p_bais.t18 VDD.t16 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X62 a_16669_n8264.t2 Nbais.t12 GND.t48 GND.t47 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X63 net4.t16 Nbais.t13 GND.t44 GND.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X64 net1.t2 Nbais.t14 GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X65 net7.t1 p_bais.t19 VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X66 net5.t2 VBN.t15 net4.t11 GND.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X67 GND.t50 a_48058_n6837.t3 GND.t49 GND.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.3e+06u l=1e+06u
X68 net3.t0 p_bais.t20 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X69 a_16669_n8264.t0 VON.t5 net3_ota.t0 GND.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X70 net4.t3 Nbais.t15 GND.t11 GND.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X71 net2.t1 Nbais.t16 GND.t42 GND.t41 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X72 VBP.t4 p_bais.t4 VDD sky130_fd_pr__res_iso_pw w=2.65e+06u l=3e+07u
X73 net4.t18 Nbais.t17 GND.t54 GND.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X74 net6.t9 VBP.t13 net7.t15 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X75 net5.t1 VBN.t16 net4.t6 GND.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X76 net4.t19 Nbais.t18 GND.t56 GND.t55 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=600000u
X77 net6.t10 VBP.t14 net7.t14 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X78 net7.t0 p_bais.t21 VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X79 net6.t2 VBP.t15 net7.t13 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X80 w_4269_n7633# Nbais.t2 VDD sky130_fd_pr__res_iso_pw w=2.65e+06u l=3e+07u
X81 net6.t3 VBP.t16 net7.t12 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X82 net5_ota.t2 VBN.t17 a_48058_n6837.t1 GND.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X83 net6.t4 VBP.t17 net7.t11 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
X84 net6_ota.t2 VOP.t3 net5_ota.t0 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X85 net6.t11 VBP.t18 net7.t10 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6.66e+06u l=600000u
R0 UBP UBP.t2 1701.44
R1 UBP.n2 UBP.t0 232.401
R2 UBP.n8 UBP.n7 188.161
R3 UBP.n18 UBP.t1 23.416
R4 UBP.n2 UBP.n1 15.764
R5 UBP.n6 UBP.n5 9.3
R6 UBP.n10 UBP.n9 9.3
R7 UBP.n4 UBP.n3 9.3
R8 UBP UBP.n26 3.438
R9 UBP.n26 UBP.n17 2.255
R10 UBP.n26 UBP.n25 2.254
R11 UBP.n4 UBP.n2 1.248
R12 UBP.n23 UBP.n21 1.137
R13 UBP.n19 UBP.n18 1.065
R14 UBP.n12 UBP.n11 1.037
R15 UBP.n15 UBP.n14 0.853
R16 UBP.n9 UBP.n8 0.705
R17 UBP.n25 UBP.n24 0.7
R18 UBP.n17 UBP.n16 0.7
R19 UBP.n11 UBP.n10 0.127
R20 UBP.n14 UBP.n13 0.041
R21 UBP.n10 UBP.n6 0.04
R22 UBP.n21 UBP.n20 0.019
R23 UBP.n15 UBP.n0 0.013
R24 UBP.n14 UBP.n12 0.009
R25 UBP.n6 UBP.n4 0.005
R26 UBP.n21 UBP.n19 0.005
R27 UBP.n16 UBP.n15 0.004
R28 UBP.n24 UBP.n23 0.004
R29 UBP.n23 UBP.n22 0.001
R30 VOP.n753 VOP.t3 735.159
R31 VOP.n753 VOP.t2 238.945
R32 VOP.n108 VOP.n107 13.176
R33 VOP.n521 VOP.n520 13.176
R34 VOP.n90 VOP.n89 9.3
R35 VOP.n234 VOP.n233 9.3
R36 VOP.n312 VOP.n311 9.3
R37 VOP.n458 VOP.n457 9.3
R38 VOP.n460 VOP.n459 9.3
R39 VOP.n208 VOP.n207 9.3
R40 VOP.n101 VOP.n100 9.3
R41 VOP.n88 VOP.n87 9.3
R42 VOP.n220 VOP.n219 9.3
R43 VOP.n231 VOP.n230 9.3
R44 VOP.n326 VOP.n325 9.3
R45 VOP.n289 VOP.n288 9.3
R46 VOP.n314 VOP.n313 9.3
R47 VOP.n472 VOP.n471 9.3
R48 VOP.n484 VOP.n483 9.3
R49 VOP.n519 VOP.n518 9.3
R50 VOP.n669 VOP.n668 9.3
R51 VOP.n710 VOP.n709 9.3
R52 VOP.n607 VOP.n606 8.043
R53 VOP.n734 VOP.n733 7.029
R54 VOP.n752 VOP.n751 6.129
R55 VOP.n300 VOP.n299 5.417
R56 VOP.n457 VOP.n456 5.081
R57 VOP.n233 VOP.n232 4.704
R58 VOP.n19 VOP.n16 4.703
R59 VOP.n279 VOP.n278 4.65
R60 VOP.n511 VOP.n510 4.65
R61 VOP.n689 VOP.n688 4.65
R62 VOP.n594 VOP.n593 4.5
R63 VOP.n20 VOP.n19 4.5
R64 VOP.n11 VOP.n10 4.5
R65 VOP.n392 VOP.n391 4.5
R66 VOP.n384 VOP.n383 4.5
R67 VOP.n32 VOP.n28 4.5
R68 VOP.n120 VOP.n119 4.5
R69 VOP.n110 VOP.n109 4.5
R70 VOP.n94 VOP.n93 4.5
R71 VOP.n81 VOP.n80 4.5
R72 VOP.n75 VOP.n74 4.5
R73 VOP.n216 VOP.n215 4.5
R74 VOP.n228 VOP.n227 4.5
R75 VOP.n246 VOP.n245 4.5
R76 VOP.n266 VOP.n265 4.5
R77 VOP.n259 VOP.n258 4.5
R78 VOP.n252 VOP.n251 4.5
R79 VOP.n274 VOP.n273 4.5
R80 VOP.n330 VOP.n329 4.5
R81 VOP.n292 VOP.n291 4.5
R82 VOP.n319 VOP.n318 4.5
R83 VOP.n307 VOP.n303 4.5
R84 VOP.n422 VOP.n412 4.5
R85 VOP.n400 VOP.n399 4.5
R86 VOP.n417 VOP.n414 4.5
R87 VOP.n464 VOP.n463 4.5
R88 VOP.n489 VOP.n488 4.5
R89 VOP.n476 VOP.n475 4.5
R90 VOP.n559 VOP.n558 4.5
R91 VOP.n523 VOP.n522 4.5
R92 VOP.n567 VOP.n566 4.5
R93 VOP.n582 VOP.n581 4.5
R94 VOP.n574 VOP.n573 4.5
R95 VOP.n40 VOP.n39 4.5
R96 VOP.n745 VOP.n744 4.5
R97 VOP.n726 VOP.n725 4.5
R98 VOP.n716 VOP.n715 4.5
R99 VOP.n704 VOP.n703 4.5
R100 VOP.n655 VOP.n654 4.5
R101 VOP.n665 VOP.n664 4.5
R102 VOP.n697 VOP.n696 4.5
R103 VOP.n691 VOP.n690 4.5
R104 VOP.n687 VOP.n686 4.5
R105 VOP.n683 VOP.n682 4.5
R106 VOP.n677 VOP.n676 4.5
R107 VOP.n615 VOP.n614 4.5
R108 VOP.n617 VOP.n607 4.473
R109 VOP.n606 VOP.t1 4.35
R110 VOP.n74 VOP.n71 4.328
R111 VOP.n581 VOP.n580 4.326
R112 VOP.n654 VOP.n651 4.141
R113 VOP.n725 VOP.n724 4.141
R114 VOP.n566 VOP.n565 3.951
R115 VOP.n303 VOP.n301 3.946
R116 VOP.n18 VOP.n17 3.764
R117 VOP.n664 VOP.n661 3.764
R118 VOP.n703 VOP.n701 3.764
R119 VOP.n391 VOP.n388 3.572
R120 VOP.n273 VOP.n272 3.569
R121 VOP.n250 VOP.n249 3.388
R122 VOP.n614 VOP.n611 3.388
R123 VOP.n676 VOP.n675 3.388
R124 VOP.n715 VOP.n714 3.388
R125 VOP.n744 VOP.n743 3.388
R126 VOP.n412 VOP.n409 3.197
R127 VOP.n258 VOP.n257 3.195
R128 VOP.n238 VOP.n237 3.033
R129 VOP.n336 VOP.n300 3.033
R130 VOP.n283 VOP.n282 3.033
R131 VOP.n512 VOP.n508 3.033
R132 VOP.n600 VOP.n599 3.033
R133 VOP.n390 VOP.n389 3.011
R134 VOP.n614 VOP.n613 3.011
R135 VOP.n676 VOP.n673 3.011
R136 VOP.n682 VOP.n680 3.011
R137 VOP.n709 VOP.n708 3.011
R138 VOP.n715 VOP.n713 3.011
R139 VOP.n744 VOP.n742 3.011
R140 VOP.n298 VOP.t0 2.856
R141 VOP.n245 VOP.n244 2.82
R142 VOP.n752 VOP.n605 2.755
R143 VOP.n28 VOP.n27 2.635
R144 VOP.n572 VOP.n571 2.635
R145 VOP.n664 VOP.n663 2.635
R146 VOP.n668 VOP.n667 2.635
R147 VOP.n696 VOP.n695 2.635
R148 VOP.n703 VOP.n702 2.635
R149 VOP.n245 VOP.n243 2.258
R150 VOP.n593 VOP.n592 2.258
R151 VOP.n654 VOP.n653 2.258
R152 VOP.n725 VOP.n723 2.258
R153 VOP VOP.n754 2.234
R154 VOP.n10 VOP.n9 1.882
R155 VOP.n383 VOP.n382 1.882
R156 VOP.n412 VOP.n411 1.882
R157 VOP.n299 VOP.n298 1.844
R158 VOP.n73 VOP.n72 1.505
R159 VOP.n258 VOP.n256 1.505
R160 VOP.n265 VOP.n264 1.505
R161 VOP.n564 VOP.n563 1.505
R162 VOP.n566 VOP.n564 1.505
R163 VOP.n573 VOP.n572 1.505
R164 VOP.n696 VOP.n694 1.505
R165 VOP.n595 VOP.n594 1.5
R166 VOP.n33 VOP.n32 1.5
R167 VOP.n21 VOP.n20 1.5
R168 VOP.n121 VOP.n120 1.5
R169 VOP.n111 VOP.n110 1.5
R170 VOP.n423 VOP.n422 1.5
R171 VOP.n401 VOP.n400 1.5
R172 VOP.n490 VOP.n489 1.5
R173 VOP.n524 VOP.n523 1.5
R174 VOP.n601 VOP.n600 1.5
R175 VOP.n583 VOP.n582 1.5
R176 VOP.n41 VOP.n40 1.5
R177 VOP.n754 VOP.n752 1.249
R178 VOP.n74 VOP.n73 1.129
R179 VOP.n80 VOP.n79 1.129
R180 VOP.n215 VOP.n214 1.129
R181 VOP.n264 VOP.n263 1.129
R182 VOP.n382 VOP.n381 1.129
R183 VOP.n391 VOP.n390 1.129
R184 VOP.n399 VOP.n398 1.129
R185 VOP.n475 VOP.n474 1.129
R186 VOP.n682 VOP.n681 1.129
R187 VOP.n746 VOP.n745 1.125
R188 VOP.n346 VOP.n336 1.042
R189 VOP.n127 VOP.n126 0.853
R190 VOP.n172 VOP.n171 0.853
R191 VOP.n347 VOP.n346 0.853
R192 VOP.n426 VOP.n425 0.853
R193 VOP.n526 VOP.n525 0.853
R194 VOP.n604 VOP.n603 0.853
R195 VOP.n227 VOP.n226 0.752
R196 VOP.n243 VOP.n242 0.752
R197 VOP.n251 VOP.n250 0.752
R198 VOP.n273 VOP.n271 0.752
R199 VOP.n291 VOP.n290 0.752
R200 VOP.n329 VOP.n328 0.752
R201 VOP.n411 VOP.n410 0.752
R202 VOP.n558 VOP.n557 0.752
R203 VOP.n581 VOP.n579 0.752
R204 VOP.n618 VOP.n617 0.75
R205 VOP.n43 VOP.n42 0.704
R206 VOP.n733 VOP.n732 0.445
R207 VOP.n613 VOP.n612 0.414
R208 VOP.n742 VOP.n741 0.414
R209 VOP.n653 VOP.n652 0.382
R210 VOP.n723 VOP.n722 0.382
R211 VOP.n39 VOP.n38 0.376
R212 VOP.n27 VOP.n26 0.376
R213 VOP.n19 VOP.n18 0.376
R214 VOP.n93 VOP.n92 0.376
R215 VOP.n109 VOP.n108 0.376
R216 VOP.n119 VOP.n118 0.376
R217 VOP.n318 VOP.n317 0.376
R218 VOP.n303 VOP.n302 0.376
R219 VOP.n414 VOP.n413 0.376
R220 VOP.n463 VOP.n462 0.376
R221 VOP.n488 VOP.n487 0.376
R222 VOP.n522 VOP.n521 0.376
R223 VOP.n592 VOP.n591 0.376
R224 VOP.n100 VOP.n99 0.189
R225 VOP.n207 VOP.n206 0.189
R226 VOP.n483 VOP.n482 0.189
R227 VOP.n518 VOP.n517 0.189
R228 VOP.n87 VOP.n86 0.177
R229 VOP.n219 VOP.n218 0.177
R230 VOP.n471 VOP.n470 0.177
R231 VOP.n510 VOP.n509 0.177
R232 VOP.n754 VOP.n753 0.171
R233 VOP.n317 VOP.n316 0.121
R234 VOP.n282 VOP.n281 0.121
R235 VOP.n617 VOP.n616 0.113
R236 VOP.n328 VOP.n327 0.109
R237 VOP.n627 VOP.n626 0.1
R238 VOP.n641 VOP.n640 0.1
R239 VOP.n663 VOP.n662 0.072
R240 VOP.n713 VOP.n712 0.072
R241 VOP.n609 VOP.n608 0.06
R242 VOP.n658 VOP.n657 0.06
R243 VOP.n670 VOP.n669 0.06
R244 VOP.n710 VOP.n707 0.06
R245 VOP.n720 VOP.n719 0.06
R246 VOP.n730 VOP.n729 0.06
R247 VOP.n739 VOP.n738 0.06
R248 VOP.n620 VOP.n619 0.06
R249 VOP.n624 VOP.n623 0.06
R250 VOP.n644 VOP.n643 0.06
R251 VOP.n648 VOP.n647 0.06
R252 VOP.n748 VOP.n747 0.06
R253 VOP.n630 VOP.n629 0.055
R254 VOP.n634 VOP.n633 0.055
R255 VOP.n638 VOP.n637 0.055
R256 VOP.n619 VOP.n618 0.052
R257 VOP.n747 VOP.n746 0.052
R258 VOP.n687 VOP.n685 0.05
R259 VOP.n697 VOP.n693 0.05
R260 VOP.n633 VOP.n632 0.05
R261 VOP.n637 VOP.n636 0.05
R262 VOP.n746 VOP.n648 0.05
R263 VOP.n684 VOP.n683 0.048
R264 VOP.n692 VOP.n691 0.048
R265 VOP.n631 VOP.n630 0.048
R266 VOP.n635 VOP.n634 0.048
R267 VOP.n104 VOP.n103 0.047
R268 VOP.n235 VOP.n234 0.047
R269 VOP.n505 VOP.n504 0.047
R270 VOP.n202 VOP.n201 0.047
R271 VOP.n238 VOP.n236 0.045
R272 VOP.n295 VOP.n294 0.045
R273 VOP.n297 VOP.n296 0.045
R274 VOP.n469 VOP.n468 0.045
R275 VOP.n157 VOP.n156 0.045
R276 VOP.n342 VOP.n341 0.045
R277 VOP.n83 VOP.n82 0.043
R278 VOP.n222 VOP.n221 0.043
R279 VOP.n261 VOP.n260 0.043
R280 VOP.n335 VOP.n334 0.043
R281 VOP.n333 VOP.n332 0.043
R282 VOP.n387 VOP.n386 0.043
R283 VOP.n417 VOP.n416 0.043
R284 VOP.n556 VOP.n555 0.043
R285 VOP.n60 VOP.n59 0.043
R286 VOP.n167 VOP.n166 0.043
R287 VOP.n377 VOP.n376 0.043
R288 VOP.n406 VOP.n405 0.043
R289 VOP.n543 VOP.n542 0.043
R290 VOP.n623 VOP.n622 0.043
R291 VOP.n647 VOP.n646 0.043
R292 VOP.n751 VOP.n750 0.043
R293 VOP.n336 VOP.n335 0.041
R294 VOP.n467 VOP.n466 0.041
R295 VOP.n346 VOP.n345 0.041
R296 VOP.n443 VOP.n442 0.041
R297 VOP.n621 VOP.n620 0.04
R298 VOP.n629 VOP.n628 0.04
R299 VOP.n645 VOP.n644 0.04
R300 VOP.n749 VOP.n748 0.04
R301 VOP.n96 VOP.n95 0.039
R302 VOP.n224 VOP.n223 0.039
R303 VOP.n252 VOP.n248 0.039
R304 VOP.n336 VOP.n297 0.039
R305 VOP.n67 VOP.n66 0.039
R306 VOP.n150 VOP.n149 0.039
R307 VOP.n171 VOP.n170 0.039
R308 VOP.n346 VOP.n205 0.039
R309 VOP.n364 VOP.n363 0.039
R310 VOP.n424 VOP.n423 0.039
R311 VOP.n639 VOP.n638 0.038
R312 VOP.n98 VOP.n97 0.037
R313 VOP.n247 VOP.n246 0.037
R314 VOP.n279 VOP.n277 0.037
R315 VOP.n284 VOP.n283 0.037
R316 VOP.n321 VOP.n320 0.037
R317 VOP.n400 VOP.n397 0.037
R318 VOP.n481 VOP.n480 0.037
R319 VOP.n514 VOP.n513 0.037
R320 VOP.n161 VOP.n160 0.037
R321 VOP.n194 VOP.n193 0.037
R322 VOP.n425 VOP.n401 0.037
R323 VOP.n499 VOP.n498 0.037
R324 VOP.n675 VOP.n674 0.036
R325 VOP.n701 VOP.n700 0.036
R326 VOP.n729 VOP.n728 0.036
R327 VOP.n738 VOP.n737 0.036
R328 VOP.n210 VOP.n209 0.035
R329 VOP.n312 VOP.n310 0.035
R330 VOP.n516 VOP.n515 0.035
R331 VOP.n122 VOP.n121 0.035
R332 VOP.n491 VOP.n490 0.035
R333 VOP.n42 VOP.n41 0.035
R334 VOP.n105 VOP.n104 0.034
R335 VOP.n266 VOP.n262 0.034
R336 VOP.n276 VOP.n275 0.034
R337 VOP.n69 VOP.n68 0.034
R338 VOP.n126 VOP.n125 0.034
R339 VOP.n159 VOP.n158 0.034
R340 VOP.n189 VOP.n188 0.034
R341 VOP.n204 VOP.n203 0.034
R342 VOP.n344 VOP.n343 0.034
R343 VOP.n408 VOP.n407 0.034
R344 VOP.n524 VOP.n502 0.034
R345 VOP.n501 VOP.n500 0.034
R346 VOP.n610 VOP.n609 0.033
R347 VOP.n719 VOP.n718 0.033
R348 VOP.n643 VOP.n642 0.033
R349 VOP.n309 VOP.n308 0.032
R350 VOP.n385 VOP.n384 0.032
R351 VOP.n506 VOP.n505 0.032
R352 VOP.n512 VOP.n511 0.032
R353 VOP.n111 VOP.n70 0.032
R354 VOP.n148 VOP.n147 0.032
R355 VOP.n169 VOP.n168 0.032
R356 VOP.n191 VOP.n190 0.032
R357 VOP.n192 VOP.n191 0.032
R358 VOP.n366 VOP.n365 0.032
R359 VOP.n367 VOP.n366 0.032
R360 VOP.n369 VOP.n368 0.032
R361 VOP.n445 VOP.n444 0.032
R362 VOP.n525 VOP.n494 0.032
R363 VOP.n44 VOP.n43 0.031
R364 VOP.n55 VOP.n54 0.031
R365 VOP.n129 VOP.n128 0.031
R366 VOP.n140 VOP.n139 0.031
R367 VOP.n174 VOP.n173 0.031
R368 VOP.n185 VOP.n184 0.031
R369 VOP.n349 VOP.n348 0.031
R370 VOP.n360 VOP.n359 0.031
R371 VOP.n428 VOP.n427 0.031
R372 VOP.n439 VOP.n438 0.031
R373 VOP.n528 VOP.n527 0.031
R374 VOP.n539 VOP.n538 0.031
R375 VOP.n659 VOP.n658 0.031
R376 VOP.n731 VOP.n730 0.031
R377 VOP.n740 VOP.n739 0.031
R378 VOP.n625 VOP.n624 0.031
R379 VOP.n626 VOP.n625 0.031
R380 VOP.n91 VOP.n90 0.03
R381 VOP.n110 VOP.n101 0.03
R382 VOP.n287 VOP.n286 0.03
R383 VOP.n523 VOP.n519 0.03
R384 VOP.n600 VOP.n598 0.03
R385 VOP.n58 VOP.n57 0.03
R386 VOP.n64 VOP.n63 0.03
R387 VOP.n124 VOP.n123 0.03
R388 VOP.n144 VOP.n143 0.03
R389 VOP.n154 VOP.n153 0.03
R390 VOP.n379 VOP.n378 0.03
R391 VOP.n403 VOP.n402 0.03
R392 VOP.n449 VOP.n448 0.03
R393 VOP.n496 VOP.n495 0.03
R394 VOP.n603 VOP.n601 0.03
R395 VOP.n40 VOP.n37 0.028
R396 VOP.n31 VOP.n30 0.028
R397 VOP.n292 VOP.n289 0.028
R398 VOP.n330 VOP.n326 0.028
R399 VOP.n324 VOP.n323 0.028
R400 VOP.n590 VOP.n589 0.028
R401 VOP.n25 VOP.n24 0.028
R402 VOP.n493 VOP.n492 0.028
R403 VOP.n545 VOP.n544 0.028
R404 VOP.n587 VOP.n586 0.028
R405 VOP.n657 VOP.n656 0.028
R406 VOP.n691 VOP.n689 0.028
R407 VOP.n642 VOP.n641 0.028
R408 VOP.n48 VOP.n47 0.027
R409 VOP.n51 VOP.n50 0.027
R410 VOP.n133 VOP.n132 0.027
R411 VOP.n136 VOP.n135 0.027
R412 VOP.n178 VOP.n177 0.027
R413 VOP.n181 VOP.n180 0.027
R414 VOP.n353 VOP.n352 0.027
R415 VOP.n356 VOP.n355 0.027
R416 VOP.n432 VOP.n431 0.027
R417 VOP.n435 VOP.n434 0.027
R418 VOP.n532 VOP.n531 0.027
R419 VOP.n535 VOP.n534 0.027
R420 VOP.n280 VOP.n279 0.026
R421 VOP.n315 VOP.n314 0.026
R422 VOP.n554 VOP.n553 0.026
R423 VOP.n541 VOP.n540 0.026
R424 VOP.n689 VOP.n687 0.026
R425 VOP.n721 VOP.n720 0.026
R426 VOP.n78 VOP.n77 0.024
R427 VOP.n85 VOP.n84 0.024
R428 VOP.n213 VOP.n212 0.024
R429 VOP.n240 VOP.n239 0.024
R430 VOP.n420 VOP.n419 0.024
R431 VOP.n478 VOP.n477 0.024
R432 VOP.n561 VOP.n560 0.024
R433 VOP.n574 VOP.n570 0.024
R434 VOP.n34 VOP.n33 0.024
R435 VOP.n62 VOP.n61 0.024
R436 VOP.n550 VOP.n549 0.024
R437 VOP.n665 VOP.n660 0.024
R438 VOP.n669 VOP.n666 0.024
R439 VOP.n704 VOP.n699 0.024
R440 VOP.n707 VOP.n706 0.024
R441 VOP.n640 VOP.n639 0.024
R442 VOP.n11 VOP.n8 0.022
R443 VOP.n8 VOP.n7 0.022
R444 VOP.n570 VOP.n569 0.022
R445 VOP.n3 VOP.n2 0.022
R446 VOP.n2 VOP.n1 0.022
R447 VOP.n549 VOP.n548 0.022
R448 VOP.n583 VOP.n552 0.022
R449 VOP.n596 VOP.n595 0.022
R450 VOP.n616 VOP.n615 0.021
R451 VOP.n671 VOP.n670 0.021
R452 VOP.n672 VOP.n671 0.021
R453 VOP.n678 VOP.n677 0.021
R454 VOP.n706 VOP.n705 0.021
R455 VOP.n711 VOP.n710 0.021
R456 VOP.n717 VOP.n716 0.021
R457 VOP.n745 VOP.n740 0.021
R458 VOP.n628 VOP.n627 0.021
R459 VOP.n30 VOP.n29 0.02
R460 VOP.n7 VOP.n6 0.02
R461 VOP.n88 VOP.n85 0.02
R462 VOP.n464 VOP.n461 0.02
R463 VOP.n569 VOP.n568 0.02
R464 VOP.n589 VOP.n588 0.02
R465 VOP.n24 VOP.n23 0.02
R466 VOP.n21 VOP.n5 0.02
R467 VOP.n1 VOP.n0 0.02
R468 VOP.n146 VOP.n145 0.02
R469 VOP.n441 VOP.n440 0.02
R470 VOP.n453 VOP.n452 0.02
R471 VOP.n548 VOP.n547 0.02
R472 VOP.n586 VOP.n585 0.02
R473 VOP.n601 VOP.n596 0.02
R474 VOP.n127 VOP.n55 0.019
R475 VOP.n128 VOP.n127 0.019
R476 VOP.n172 VOP.n140 0.019
R477 VOP.n173 VOP.n172 0.019
R478 VOP.n347 VOP.n185 0.019
R479 VOP.n348 VOP.n347 0.019
R480 VOP.n426 VOP.n360 0.019
R481 VOP.n427 VOP.n426 0.019
R482 VOP.n526 VOP.n439 0.019
R483 VOP.n527 VOP.n526 0.019
R484 VOP.n615 VOP.n610 0.019
R485 VOP.n655 VOP.n650 0.019
R486 VOP.n677 VOP.n672 0.019
R487 VOP.n683 VOP.n679 0.019
R488 VOP.n716 VOP.n711 0.019
R489 VOP.n727 VOP.n726 0.019
R490 VOP.n745 VOP.n731 0.019
R491 VOP.n736 VOP.n735 0.019
R492 VOP.n622 VOP.n621 0.019
R493 VOP.n646 VOP.n645 0.019
R494 VOP.n750 VOP.n749 0.019
R495 VOP.n15 VOP.n14 0.018
R496 VOP.n229 VOP.n228 0.018
R497 VOP.n323 VOP.n322 0.018
R498 VOP.n479 VOP.n478 0.018
R499 VOP.n578 VOP.n577 0.018
R500 VOP.n41 VOP.n34 0.018
R501 VOP.n113 VOP.n112 0.018
R502 VOP.n152 VOP.n151 0.018
R503 VOP.n339 VOP.n338 0.018
R504 VOP.n362 VOP.n361 0.018
R505 VOP.n447 VOP.n446 0.018
R506 VOP.n450 VOP.n449 0.018
R507 VOP.n494 VOP.n493 0.018
R508 VOP.n212 VOP.n211 0.017
R509 VOP.n254 VOP.n253 0.017
R510 VOP.n269 VOP.n268 0.017
R511 VOP.n286 VOP.n285 0.017
R512 VOP.n308 VOP.n307 0.017
R513 VOP.n305 VOP.n304 0.017
R514 VOP.n395 VOP.n394 0.017
R515 VOP.n485 VOP.n484 0.017
R516 VOP.n568 VOP.n567 0.017
R517 VOP.n23 VOP.n22 0.017
R518 VOP.n5 VOP.n4 0.017
R519 VOP.n63 VOP.n62 0.017
R520 VOP.n125 VOP.n124 0.017
R521 VOP.n115 VOP.n114 0.017
R522 VOP.n143 VOP.n142 0.017
R523 VOP.n153 VOP.n152 0.017
R524 VOP.n165 VOP.n164 0.017
R525 VOP.n164 VOP.n163 0.017
R526 VOP.n196 VOP.n195 0.017
R527 VOP.n197 VOP.n196 0.017
R528 VOP.n199 VOP.n198 0.017
R529 VOP.n370 VOP.n369 0.017
R530 VOP.n372 VOP.n371 0.017
R531 VOP.n375 VOP.n374 0.017
R532 VOP.n452 VOP.n451 0.017
R533 VOP.n455 VOP.n454 0.017
R534 VOP.n547 VOP.n546 0.017
R535 VOP.n552 VOP.n551 0.017
R536 VOP.n585 VOP.n584 0.017
R537 VOP.n604 VOP.n539 0.016
R538 VOP.n666 VOP.n665 0.016
R539 VOP.n698 VOP.n697 0.016
R540 VOP.n705 VOP.n704 0.016
R541 VOP.n255 VOP.n254 0.015
R542 VOP.n275 VOP.n274 0.015
R543 VOP.n394 VOP.n393 0.015
R544 VOP.n126 VOP.n111 0.015
R545 VOP.n188 VOP.n187 0.015
R546 VOP.n200 VOP.n199 0.015
R547 VOP.n340 VOP.n339 0.015
R548 VOP.n373 VOP.n372 0.015
R549 VOP.n374 VOP.n373 0.015
R550 VOP.n525 VOP.n524 0.015
R551 VOP.n546 VOP.n545 0.015
R552 VOP.n605 VOP.n604 0.014
R553 VOP.n656 VOP.n655 0.014
R554 VOP.n679 VOP.n678 0.014
R555 VOP.n699 VOP.n698 0.014
R556 VOP.n726 VOP.n721 0.014
R557 VOP.n14 VOP.n13 0.013
R558 VOP.n106 VOP.n105 0.013
R559 VOP.n120 VOP.n117 0.013
R560 VOP.n217 VOP.n216 0.013
R561 VOP.n220 VOP.n217 0.013
R562 VOP.n473 VOP.n472 0.013
R563 VOP.n476 VOP.n473 0.013
R564 VOP.n489 VOP.n485 0.013
R565 VOP.n507 VOP.n506 0.013
R566 VOP.n577 VOP.n576 0.013
R567 VOP.n57 VOP.n56 0.013
R568 VOP.n121 VOP.n115 0.013
R569 VOP.n145 VOP.n144 0.013
R570 VOP.n155 VOP.n154 0.013
R571 VOP.n163 VOP.n162 0.013
R572 VOP.n187 VOP.n186 0.013
R573 VOP.n198 VOP.n197 0.013
R574 VOP.n401 VOP.n379 0.013
R575 VOP.n446 VOP.n445 0.013
R576 VOP.n448 VOP.n447 0.013
R577 VOP.n490 VOP.n455 0.013
R578 VOP.n49 VOP.n48 0.012
R579 VOP.n50 VOP.n49 0.012
R580 VOP.n134 VOP.n133 0.012
R581 VOP.n135 VOP.n134 0.012
R582 VOP.n179 VOP.n178 0.012
R583 VOP.n180 VOP.n179 0.012
R584 VOP.n354 VOP.n353 0.012
R585 VOP.n355 VOP.n354 0.012
R586 VOP.n433 VOP.n432 0.012
R587 VOP.n434 VOP.n433 0.012
R588 VOP.n533 VOP.n532 0.012
R589 VOP.n534 VOP.n533 0.012
R590 VOP.n209 VOP.n208 0.011
R591 VOP.n211 VOP.n210 0.011
R592 VOP.n246 VOP.n241 0.011
R593 VOP.n285 VOP.n284 0.011
R594 VOP.n310 VOP.n309 0.011
R595 VOP.n515 VOP.n514 0.011
R596 VOP.n513 VOP.n512 0.011
R597 VOP.n594 VOP.n590 0.011
R598 VOP.n114 VOP.n113 0.011
R599 VOP.n142 VOP.n141 0.011
R600 VOP.n147 VOP.n146 0.011
R601 VOP.n170 VOP.n169 0.011
R602 VOP.n195 VOP.n194 0.011
R603 VOP.n205 VOP.n204 0.011
R604 VOP.n338 VOP.n337 0.011
R605 VOP.n368 VOP.n367 0.011
R606 VOP.n371 VOP.n370 0.011
R607 VOP.n404 VOP.n403 0.011
R608 VOP.n500 VOP.n499 0.011
R609 VOP.n498 VOP.n497 0.011
R610 VOP.n595 VOP.n587 0.011
R611 VOP.n46 VOP.n45 0.011
R612 VOP.n53 VOP.n52 0.011
R613 VOP.n131 VOP.n130 0.011
R614 VOP.n138 VOP.n137 0.011
R615 VOP.n176 VOP.n175 0.011
R616 VOP.n183 VOP.n182 0.011
R617 VOP.n351 VOP.n350 0.011
R618 VOP.n358 VOP.n357 0.011
R619 VOP.n430 VOP.n429 0.011
R620 VOP.n437 VOP.n436 0.011
R621 VOP.n530 VOP.n529 0.011
R622 VOP.n537 VOP.n536 0.011
R623 VOP.n32 VOP.n31 0.009
R624 VOP.n95 VOP.n94 0.009
R625 VOP.n97 VOP.n96 0.009
R626 VOP.n231 VOP.n229 0.009
R627 VOP.n270 VOP.n269 0.009
R628 VOP.n277 VOP.n276 0.009
R629 VOP.n322 VOP.n321 0.009
R630 VOP.n306 VOP.n305 0.009
R631 VOP.n384 VOP.n380 0.009
R632 VOP.n422 VOP.n421 0.009
R633 VOP.n461 VOP.n460 0.009
R634 VOP.n480 VOP.n479 0.009
R635 VOP.n484 VOP.n481 0.009
R636 VOP.n33 VOP.n25 0.009
R637 VOP.n22 VOP.n21 0.009
R638 VOP.n66 VOP.n65 0.009
R639 VOP.n68 VOP.n67 0.009
R640 VOP.n151 VOP.n150 0.009
R641 VOP.n190 VOP.n189 0.009
R642 VOP.n345 VOP.n344 0.009
R643 VOP.n363 VOP.n362 0.009
R644 VOP.n451 VOP.n450 0.009
R645 VOP.n454 VOP.n453 0.009
R646 VOP.n685 VOP.n684 0.009
R647 VOP.n693 VOP.n692 0.009
R648 VOP.n632 VOP.n631 0.009
R649 VOP.n636 VOP.n635 0.009
R650 VOP.n603 VOP.n602 0.008
R651 VOP.n77 VOP.n76 0.007
R652 VOP.n221 VOP.n220 0.007
R653 VOP.n248 VOP.n247 0.007
R654 VOP.n259 VOP.n255 0.007
R655 VOP.n267 VOP.n266 0.007
R656 VOP.n397 VOP.n396 0.007
R657 VOP.n562 VOP.n561 0.007
R658 VOP.n567 VOP.n562 0.007
R659 VOP.n65 VOP.n64 0.007
R660 VOP.n171 VOP.n161 0.007
R661 VOP.n425 VOP.n424 0.007
R662 VOP.n442 VOP.n441 0.007
R663 VOP.n584 VOP.n583 0.007
R664 VOP.n650 VOP.n649 0.007
R665 VOP.n660 VOP.n659 0.007
R666 VOP.n718 VOP.n717 0.007
R667 VOP.n728 VOP.n727 0.007
R668 VOP.n45 VOP.n44 0.006
R669 VOP.n47 VOP.n46 0.006
R670 VOP.n52 VOP.n51 0.006
R671 VOP.n54 VOP.n53 0.006
R672 VOP.n130 VOP.n129 0.006
R673 VOP.n132 VOP.n131 0.006
R674 VOP.n137 VOP.n136 0.006
R675 VOP.n139 VOP.n138 0.006
R676 VOP.n175 VOP.n174 0.006
R677 VOP.n177 VOP.n176 0.006
R678 VOP.n182 VOP.n181 0.006
R679 VOP.n184 VOP.n183 0.006
R680 VOP.n350 VOP.n349 0.006
R681 VOP.n352 VOP.n351 0.006
R682 VOP.n357 VOP.n356 0.006
R683 VOP.n359 VOP.n358 0.006
R684 VOP.n429 VOP.n428 0.006
R685 VOP.n431 VOP.n430 0.006
R686 VOP.n436 VOP.n435 0.006
R687 VOP.n438 VOP.n437 0.006
R688 VOP.n529 VOP.n528 0.006
R689 VOP.n531 VOP.n530 0.006
R690 VOP.n536 VOP.n535 0.006
R691 VOP.n538 VOP.n537 0.006
R692 VOP.n12 VOP.n11 0.005
R693 VOP.n76 VOP.n75 0.005
R694 VOP.n81 VOP.n78 0.005
R695 VOP.n216 VOP.n213 0.005
R696 VOP.n225 VOP.n224 0.005
R697 VOP.n262 VOP.n261 0.005
R698 VOP.n268 VOP.n267 0.005
R699 VOP.n283 VOP.n280 0.005
R700 VOP.n326 VOP.n324 0.005
R701 VOP.n386 VOP.n385 0.005
R702 VOP.n393 VOP.n392 0.005
R703 VOP.n400 VOP.n395 0.005
R704 VOP.n416 VOP.n415 0.005
R705 VOP.n466 VOP.n465 0.005
R706 VOP.n472 VOP.n469 0.005
R707 VOP.n477 VOP.n476 0.005
R708 VOP.n504 VOP.n503 0.005
R709 VOP.n4 VOP.n3 0.005
R710 VOP.n160 VOP.n159 0.005
R711 VOP.n166 VOP.n165 0.005
R712 VOP.n193 VOP.n192 0.005
R713 VOP.n376 VOP.n375 0.005
R714 VOP.n407 VOP.n406 0.005
R715 VOP.n405 VOP.n404 0.005
R716 VOP.n492 VOP.n491 0.005
R717 VOP.n497 VOP.n496 0.005
R718 VOP.n735 VOP.n734 0.005
R719 VOP.n737 VOP.n736 0.004
R720 VOP.n13 VOP.n12 0.003
R721 VOP.n84 VOP.n83 0.003
R722 VOP.n103 VOP.n102 0.003
R723 VOP.n223 VOP.n222 0.003
R724 VOP.n228 VOP.n225 0.003
R725 VOP.n234 VOP.n231 0.003
R726 VOP.n236 VOP.n235 0.003
R727 VOP.n239 VOP.n238 0.003
R728 VOP.n241 VOP.n240 0.003
R729 VOP.n253 VOP.n252 0.003
R730 VOP.n274 VOP.n270 0.003
R731 VOP.n289 VOP.n287 0.003
R732 VOP.n334 VOP.n333 0.003
R733 VOP.n319 VOP.n315 0.003
R734 VOP.n392 VOP.n387 0.003
R735 VOP.n421 VOP.n420 0.003
R736 VOP.n419 VOP.n418 0.003
R737 VOP.n519 VOP.n516 0.003
R738 VOP.n559 VOP.n556 0.003
R739 VOP.n560 VOP.n559 0.003
R740 VOP.n575 VOP.n574 0.003
R741 VOP.n576 VOP.n575 0.003
R742 VOP.n582 VOP.n578 0.003
R743 VOP.n61 VOP.n60 0.003
R744 VOP.n70 VOP.n69 0.003
R745 VOP.n123 VOP.n122 0.003
R746 VOP.n149 VOP.n148 0.003
R747 VOP.n156 VOP.n155 0.003
R748 VOP.n158 VOP.n157 0.003
R749 VOP.n343 VOP.n342 0.003
R750 VOP.n365 VOP.n364 0.003
R751 VOP.n378 VOP.n377 0.003
R752 VOP.n423 VOP.n408 0.003
R753 VOP.n544 VOP.n543 0.003
R754 VOP.n551 VOP.n550 0.003
R755 VOP.n40 VOP.n35 0.001
R756 VOP.n37 VOP.n36 0.001
R757 VOP.n20 VOP.n15 0.001
R758 VOP.n82 VOP.n81 0.001
R759 VOP.n90 VOP.n88 0.001
R760 VOP.n94 VOP.n91 0.001
R761 VOP.n101 VOP.n98 0.001
R762 VOP.n110 VOP.n106 0.001
R763 VOP.n120 VOP.n116 0.001
R764 VOP.n260 VOP.n259 0.001
R765 VOP.n293 VOP.n292 0.001
R766 VOP.n294 VOP.n293 0.001
R767 VOP.n296 VOP.n295 0.001
R768 VOP.n332 VOP.n331 0.001
R769 VOP.n331 VOP.n330 0.001
R770 VOP.n320 VOP.n319 0.001
R771 VOP.n314 VOP.n312 0.001
R772 VOP.n307 VOP.n306 0.001
R773 VOP.n418 VOP.n417 0.001
R774 VOP.n460 VOP.n458 0.001
R775 VOP.n465 VOP.n464 0.001
R776 VOP.n468 VOP.n467 0.001
R777 VOP.n489 VOP.n486 0.001
R778 VOP.n523 VOP.n507 0.001
R779 VOP.n555 VOP.n554 0.001
R780 VOP.n598 VOP.n597 0.001
R781 VOP.n59 VOP.n58 0.001
R782 VOP.n168 VOP.n167 0.001
R783 VOP.n201 VOP.n200 0.001
R784 VOP.n203 VOP.n202 0.001
R785 VOP.n341 VOP.n340 0.001
R786 VOP.n444 VOP.n443 0.001
R787 VOP.n502 VOP.n501 0.001
R788 VOP.n542 VOP.n541 0.001
R789 net6.n3439 net6.n3438 13.176
R790 net6.n3078 net6.n3077 13.176
R791 net6.n2717 net6.n2716 13.176
R792 net6.n2356 net6.n2355 13.176
R793 net6.n1995 net6.n1994 13.176
R794 net6.n1633 net6.n1632 13.176
R795 net6.n1271 net6.n1270 13.176
R796 net6.n909 net6.n908 13.176
R797 net6.n547 net6.n546 13.176
R798 net6.n185 net6.n184 13.176
R799 net6.n3473 net6.n3472 9.3
R800 net6.n3599 net6.n3598 9.3
R801 net6.n3602 net6.n3601 9.3
R802 net6.n3610 net6.n3609 9.3
R803 net6.n3649 net6.n3648 9.3
R804 net6.n3660 net6.n3659 9.3
R805 net6.n3651 net6.n3650 9.3
R806 net6.n3639 net6.n3638 9.3
R807 net6.n3641 net6.n3640 9.3
R808 net6.n3613 net6.n3612 9.3
R809 net6.n3589 net6.n3588 9.3
R810 net6.n3444 net6.n3443 9.3
R811 net6.n3475 net6.n3474 9.3
R812 net6.n3360 net6.n3359 9.3
R813 net6.n3348 net6.n3347 9.3
R814 net6.n3346 net6.n3345 9.3
R815 net6.n3112 net6.n3111 9.3
R816 net6.n3238 net6.n3237 9.3
R817 net6.n3241 net6.n3240 9.3
R818 net6.n3249 net6.n3248 9.3
R819 net6.n3288 net6.n3287 9.3
R820 net6.n3299 net6.n3298 9.3
R821 net6.n3290 net6.n3289 9.3
R822 net6.n3278 net6.n3277 9.3
R823 net6.n3280 net6.n3279 9.3
R824 net6.n3252 net6.n3251 9.3
R825 net6.n3228 net6.n3227 9.3
R826 net6.n3083 net6.n3082 9.3
R827 net6.n3114 net6.n3113 9.3
R828 net6.n2999 net6.n2998 9.3
R829 net6.n2987 net6.n2986 9.3
R830 net6.n2985 net6.n2984 9.3
R831 net6.n2751 net6.n2750 9.3
R832 net6.n2877 net6.n2876 9.3
R833 net6.n2880 net6.n2879 9.3
R834 net6.n2888 net6.n2887 9.3
R835 net6.n2927 net6.n2926 9.3
R836 net6.n2938 net6.n2937 9.3
R837 net6.n2929 net6.n2928 9.3
R838 net6.n2917 net6.n2916 9.3
R839 net6.n2919 net6.n2918 9.3
R840 net6.n2891 net6.n2890 9.3
R841 net6.n2867 net6.n2866 9.3
R842 net6.n2722 net6.n2721 9.3
R843 net6.n2753 net6.n2752 9.3
R844 net6.n2638 net6.n2637 9.3
R845 net6.n2626 net6.n2625 9.3
R846 net6.n2624 net6.n2623 9.3
R847 net6.n2390 net6.n2389 9.3
R848 net6.n2516 net6.n2515 9.3
R849 net6.n2519 net6.n2518 9.3
R850 net6.n2527 net6.n2526 9.3
R851 net6.n2566 net6.n2565 9.3
R852 net6.n2577 net6.n2576 9.3
R853 net6.n2568 net6.n2567 9.3
R854 net6.n2556 net6.n2555 9.3
R855 net6.n2558 net6.n2557 9.3
R856 net6.n2530 net6.n2529 9.3
R857 net6.n2506 net6.n2505 9.3
R858 net6.n2361 net6.n2360 9.3
R859 net6.n2392 net6.n2391 9.3
R860 net6.n2277 net6.n2276 9.3
R861 net6.n2265 net6.n2264 9.3
R862 net6.n2263 net6.n2262 9.3
R863 net6.n2029 net6.n2028 9.3
R864 net6.n2155 net6.n2154 9.3
R865 net6.n2158 net6.n2157 9.3
R866 net6.n2166 net6.n2165 9.3
R867 net6.n2205 net6.n2204 9.3
R868 net6.n2216 net6.n2215 9.3
R869 net6.n2207 net6.n2206 9.3
R870 net6.n2195 net6.n2194 9.3
R871 net6.n2197 net6.n2196 9.3
R872 net6.n2169 net6.n2168 9.3
R873 net6.n2145 net6.n2144 9.3
R874 net6.n2000 net6.n1999 9.3
R875 net6.n2031 net6.n2030 9.3
R876 net6.n1916 net6.n1915 9.3
R877 net6.n1904 net6.n1903 9.3
R878 net6.n1902 net6.n1901 9.3
R879 net6.n1667 net6.n1666 9.3
R880 net6.n1793 net6.n1792 9.3
R881 net6.n1796 net6.n1795 9.3
R882 net6.n1804 net6.n1803 9.3
R883 net6.n1843 net6.n1842 9.3
R884 net6.n1854 net6.n1853 9.3
R885 net6.n1845 net6.n1844 9.3
R886 net6.n1833 net6.n1832 9.3
R887 net6.n1835 net6.n1834 9.3
R888 net6.n1807 net6.n1806 9.3
R889 net6.n1783 net6.n1782 9.3
R890 net6.n1638 net6.n1637 9.3
R891 net6.n1669 net6.n1668 9.3
R892 net6.n1554 net6.n1553 9.3
R893 net6.n1542 net6.n1541 9.3
R894 net6.n1540 net6.n1539 9.3
R895 net6.n1305 net6.n1304 9.3
R896 net6.n1431 net6.n1430 9.3
R897 net6.n1434 net6.n1433 9.3
R898 net6.n1442 net6.n1441 9.3
R899 net6.n1481 net6.n1480 9.3
R900 net6.n1492 net6.n1491 9.3
R901 net6.n1483 net6.n1482 9.3
R902 net6.n1471 net6.n1470 9.3
R903 net6.n1473 net6.n1472 9.3
R904 net6.n1445 net6.n1444 9.3
R905 net6.n1421 net6.n1420 9.3
R906 net6.n1276 net6.n1275 9.3
R907 net6.n1307 net6.n1306 9.3
R908 net6.n1192 net6.n1191 9.3
R909 net6.n1180 net6.n1179 9.3
R910 net6.n1178 net6.n1177 9.3
R911 net6.n943 net6.n942 9.3
R912 net6.n1069 net6.n1068 9.3
R913 net6.n1072 net6.n1071 9.3
R914 net6.n1080 net6.n1079 9.3
R915 net6.n1119 net6.n1118 9.3
R916 net6.n1130 net6.n1129 9.3
R917 net6.n1121 net6.n1120 9.3
R918 net6.n1109 net6.n1108 9.3
R919 net6.n1111 net6.n1110 9.3
R920 net6.n1083 net6.n1082 9.3
R921 net6.n1059 net6.n1058 9.3
R922 net6.n914 net6.n913 9.3
R923 net6.n945 net6.n944 9.3
R924 net6.n830 net6.n829 9.3
R925 net6.n818 net6.n817 9.3
R926 net6.n816 net6.n815 9.3
R927 net6.n581 net6.n580 9.3
R928 net6.n707 net6.n706 9.3
R929 net6.n710 net6.n709 9.3
R930 net6.n718 net6.n717 9.3
R931 net6.n757 net6.n756 9.3
R932 net6.n768 net6.n767 9.3
R933 net6.n759 net6.n758 9.3
R934 net6.n747 net6.n746 9.3
R935 net6.n749 net6.n748 9.3
R936 net6.n721 net6.n720 9.3
R937 net6.n697 net6.n696 9.3
R938 net6.n552 net6.n551 9.3
R939 net6.n583 net6.n582 9.3
R940 net6.n468 net6.n467 9.3
R941 net6.n456 net6.n455 9.3
R942 net6.n454 net6.n453 9.3
R943 net6.n219 net6.n218 9.3
R944 net6.n345 net6.n344 9.3
R945 net6.n348 net6.n347 9.3
R946 net6.n356 net6.n355 9.3
R947 net6.n395 net6.n394 9.3
R948 net6.n406 net6.n405 9.3
R949 net6.n397 net6.n396 9.3
R950 net6.n385 net6.n384 9.3
R951 net6.n387 net6.n386 9.3
R952 net6.n359 net6.n358 9.3
R953 net6.n335 net6.n334 9.3
R954 net6.n190 net6.n189 9.3
R955 net6.n221 net6.n220 9.3
R956 net6.n106 net6.n105 9.3
R957 net6.n94 net6.n93 9.3
R958 net6.n92 net6.n91 9.3
R959 net6.n3370 net6.n3369 8.454
R960 net6.n3009 net6.n3008 8.454
R961 net6.n2648 net6.n2647 8.454
R962 net6.n2287 net6.n2286 8.454
R963 net6.n1926 net6.n1925 8.454
R964 net6.n1564 net6.n1563 8.454
R965 net6.n1202 net6.n1201 8.454
R966 net6.n840 net6.n839 8.454
R967 net6.n478 net6.n477 8.454
R968 net6.n116 net6.n115 8.454
R969 net6.n3671 net6.n3670 8.454
R970 net6.n3310 net6.n3309 8.454
R971 net6.n2949 net6.n2948 8.454
R972 net6.n2588 net6.n2587 8.454
R973 net6.n2227 net6.n2226 8.454
R974 net6.n1865 net6.n1864 8.454
R975 net6.n1503 net6.n1502 8.454
R976 net6.n1141 net6.n1140 8.454
R977 net6.n779 net6.n778 8.454
R978 net6.n417 net6.n416 8.454
R979 net6.n28 net6.t6 6.137
R980 net6.n38 net6.t5 6.131
R981 net6.n3601 net6.n3600 5.458
R982 net6.n3240 net6.n3239 5.458
R983 net6.n2879 net6.n2878 5.458
R984 net6.n2518 net6.n2517 5.458
R985 net6.n2157 net6.n2156 5.458
R986 net6.n1795 net6.n1794 5.458
R987 net6.n1433 net6.n1432 5.458
R988 net6.n1071 net6.n1070 5.458
R989 net6.n709 net6.n708 5.458
R990 net6.n347 net6.n346 5.458
R991 net6.n3472 net6.n3471 5.081
R992 net6.n3111 net6.n3110 5.081
R993 net6.n2750 net6.n2749 5.081
R994 net6.n2389 net6.n2388 5.081
R995 net6.n2028 net6.n2027 5.081
R996 net6.n1666 net6.n1665 5.081
R997 net6.n1304 net6.n1303 5.081
R998 net6.n942 net6.n941 5.081
R999 net6.n580 net6.n579 5.081
R1000 net6.n218 net6.n217 5.081
R1001 net6.n3338 net6.n3337 4.65
R1002 net6.n3465 net6.n3464 4.65
R1003 net6.n2977 net6.n2976 4.65
R1004 net6.n3104 net6.n3103 4.65
R1005 net6.n2616 net6.n2615 4.65
R1006 net6.n2743 net6.n2742 4.65
R1007 net6.n2255 net6.n2254 4.65
R1008 net6.n2382 net6.n2381 4.65
R1009 net6.n1894 net6.n1893 4.65
R1010 net6.n2021 net6.n2020 4.65
R1011 net6.n1532 net6.n1531 4.65
R1012 net6.n1659 net6.n1658 4.65
R1013 net6.n1170 net6.n1169 4.65
R1014 net6.n1297 net6.n1296 4.65
R1015 net6.n808 net6.n807 4.65
R1016 net6.n935 net6.n934 4.65
R1017 net6.n446 net6.n445 4.65
R1018 net6.n573 net6.n572 4.65
R1019 net6.n84 net6.n83 4.65
R1020 net6.n211 net6.n210 4.65
R1021 net6.n3353 net6.n3352 4.5
R1022 net6.n3629 net6.n3628 4.5
R1023 net6.n3623 net6.n3580 4.5
R1024 net6.n3635 net6.n3576 4.5
R1025 net6.n3645 net6.n3644 4.5
R1026 net6.n3664 net6.n3663 4.5
R1027 net6.n3653 net6.n3573 4.5
R1028 net6.n3619 net6.n3618 4.5
R1029 net6.n3606 net6.n3582 4.5
R1030 net6.n3596 net6.n3595 4.5
R1031 net6.n3586 net6.n3584 4.5
R1032 net6.n3441 net6.n3440 4.5
R1033 net6.n3478 net6.n3477 4.5
R1034 net6.n3459 net6.n3450 4.5
R1035 net6.n3407 net6.n3404 4.5
R1036 net6.n3455 net6.n3454 4.5
R1037 net6.n3334 net6.n3333 4.5
R1038 net6.n3364 net6.n3363 4.5
R1039 net6.n2992 net6.n2991 4.5
R1040 net6.n3268 net6.n3267 4.5
R1041 net6.n3262 net6.n3219 4.5
R1042 net6.n3274 net6.n3215 4.5
R1043 net6.n3284 net6.n3283 4.5
R1044 net6.n3303 net6.n3302 4.5
R1045 net6.n3292 net6.n3212 4.5
R1046 net6.n3258 net6.n3257 4.5
R1047 net6.n3245 net6.n3221 4.5
R1048 net6.n3235 net6.n3234 4.5
R1049 net6.n3225 net6.n3223 4.5
R1050 net6.n3080 net6.n3079 4.5
R1051 net6.n3117 net6.n3116 4.5
R1052 net6.n3098 net6.n3089 4.5
R1053 net6.n3046 net6.n3043 4.5
R1054 net6.n3094 net6.n3093 4.5
R1055 net6.n2973 net6.n2972 4.5
R1056 net6.n3003 net6.n3002 4.5
R1057 net6.n2631 net6.n2630 4.5
R1058 net6.n2907 net6.n2906 4.5
R1059 net6.n2901 net6.n2858 4.5
R1060 net6.n2913 net6.n2854 4.5
R1061 net6.n2923 net6.n2922 4.5
R1062 net6.n2942 net6.n2941 4.5
R1063 net6.n2931 net6.n2851 4.5
R1064 net6.n2897 net6.n2896 4.5
R1065 net6.n2884 net6.n2860 4.5
R1066 net6.n2874 net6.n2873 4.5
R1067 net6.n2864 net6.n2862 4.5
R1068 net6.n2719 net6.n2718 4.5
R1069 net6.n2756 net6.n2755 4.5
R1070 net6.n2737 net6.n2728 4.5
R1071 net6.n2685 net6.n2682 4.5
R1072 net6.n2733 net6.n2732 4.5
R1073 net6.n2612 net6.n2611 4.5
R1074 net6.n2642 net6.n2641 4.5
R1075 net6.n2270 net6.n2269 4.5
R1076 net6.n2546 net6.n2545 4.5
R1077 net6.n2540 net6.n2497 4.5
R1078 net6.n2552 net6.n2493 4.5
R1079 net6.n2562 net6.n2561 4.5
R1080 net6.n2581 net6.n2580 4.5
R1081 net6.n2570 net6.n2490 4.5
R1082 net6.n2536 net6.n2535 4.5
R1083 net6.n2523 net6.n2499 4.5
R1084 net6.n2513 net6.n2512 4.5
R1085 net6.n2503 net6.n2501 4.5
R1086 net6.n2358 net6.n2357 4.5
R1087 net6.n2395 net6.n2394 4.5
R1088 net6.n2376 net6.n2367 4.5
R1089 net6.n2324 net6.n2321 4.5
R1090 net6.n2372 net6.n2371 4.5
R1091 net6.n2251 net6.n2250 4.5
R1092 net6.n2281 net6.n2280 4.5
R1093 net6.n1909 net6.n1908 4.5
R1094 net6.n2185 net6.n2184 4.5
R1095 net6.n2179 net6.n2136 4.5
R1096 net6.n2191 net6.n2132 4.5
R1097 net6.n2201 net6.n2200 4.5
R1098 net6.n2220 net6.n2219 4.5
R1099 net6.n2209 net6.n2129 4.5
R1100 net6.n2175 net6.n2174 4.5
R1101 net6.n2162 net6.n2138 4.5
R1102 net6.n2152 net6.n2151 4.5
R1103 net6.n2142 net6.n2140 4.5
R1104 net6.n1997 net6.n1996 4.5
R1105 net6.n2034 net6.n2033 4.5
R1106 net6.n2015 net6.n2006 4.5
R1107 net6.n1963 net6.n1960 4.5
R1108 net6.n2011 net6.n2010 4.5
R1109 net6.n1890 net6.n1889 4.5
R1110 net6.n1920 net6.n1919 4.5
R1111 net6.n1547 net6.n1546 4.5
R1112 net6.n1823 net6.n1822 4.5
R1113 net6.n1817 net6.n1774 4.5
R1114 net6.n1829 net6.n1770 4.5
R1115 net6.n1839 net6.n1838 4.5
R1116 net6.n1858 net6.n1857 4.5
R1117 net6.n1847 net6.n1767 4.5
R1118 net6.n1813 net6.n1812 4.5
R1119 net6.n1800 net6.n1776 4.5
R1120 net6.n1790 net6.n1789 4.5
R1121 net6.n1780 net6.n1778 4.5
R1122 net6.n1635 net6.n1634 4.5
R1123 net6.n1672 net6.n1671 4.5
R1124 net6.n1653 net6.n1644 4.5
R1125 net6.n1601 net6.n1598 4.5
R1126 net6.n1649 net6.n1648 4.5
R1127 net6.n1528 net6.n1527 4.5
R1128 net6.n1558 net6.n1557 4.5
R1129 net6.n1185 net6.n1184 4.5
R1130 net6.n1461 net6.n1460 4.5
R1131 net6.n1455 net6.n1412 4.5
R1132 net6.n1467 net6.n1408 4.5
R1133 net6.n1477 net6.n1476 4.5
R1134 net6.n1496 net6.n1495 4.5
R1135 net6.n1485 net6.n1405 4.5
R1136 net6.n1451 net6.n1450 4.5
R1137 net6.n1438 net6.n1414 4.5
R1138 net6.n1428 net6.n1427 4.5
R1139 net6.n1418 net6.n1416 4.5
R1140 net6.n1273 net6.n1272 4.5
R1141 net6.n1310 net6.n1309 4.5
R1142 net6.n1291 net6.n1282 4.5
R1143 net6.n1239 net6.n1236 4.5
R1144 net6.n1287 net6.n1286 4.5
R1145 net6.n1166 net6.n1165 4.5
R1146 net6.n1196 net6.n1195 4.5
R1147 net6.n823 net6.n822 4.5
R1148 net6.n1099 net6.n1098 4.5
R1149 net6.n1093 net6.n1050 4.5
R1150 net6.n1105 net6.n1046 4.5
R1151 net6.n1115 net6.n1114 4.5
R1152 net6.n1134 net6.n1133 4.5
R1153 net6.n1123 net6.n1043 4.5
R1154 net6.n1089 net6.n1088 4.5
R1155 net6.n1076 net6.n1052 4.5
R1156 net6.n1066 net6.n1065 4.5
R1157 net6.n1056 net6.n1054 4.5
R1158 net6.n911 net6.n910 4.5
R1159 net6.n948 net6.n947 4.5
R1160 net6.n929 net6.n920 4.5
R1161 net6.n877 net6.n874 4.5
R1162 net6.n925 net6.n924 4.5
R1163 net6.n804 net6.n803 4.5
R1164 net6.n834 net6.n833 4.5
R1165 net6.n461 net6.n460 4.5
R1166 net6.n737 net6.n736 4.5
R1167 net6.n731 net6.n688 4.5
R1168 net6.n743 net6.n684 4.5
R1169 net6.n753 net6.n752 4.5
R1170 net6.n772 net6.n771 4.5
R1171 net6.n761 net6.n681 4.5
R1172 net6.n727 net6.n726 4.5
R1173 net6.n714 net6.n690 4.5
R1174 net6.n704 net6.n703 4.5
R1175 net6.n694 net6.n692 4.5
R1176 net6.n549 net6.n548 4.5
R1177 net6.n586 net6.n585 4.5
R1178 net6.n567 net6.n558 4.5
R1179 net6.n515 net6.n512 4.5
R1180 net6.n563 net6.n562 4.5
R1181 net6.n442 net6.n441 4.5
R1182 net6.n472 net6.n471 4.5
R1183 net6.n99 net6.n98 4.5
R1184 net6.n375 net6.n374 4.5
R1185 net6.n369 net6.n326 4.5
R1186 net6.n381 net6.n322 4.5
R1187 net6.n391 net6.n390 4.5
R1188 net6.n410 net6.n409 4.5
R1189 net6.n399 net6.n319 4.5
R1190 net6.n365 net6.n364 4.5
R1191 net6.n352 net6.n328 4.5
R1192 net6.n342 net6.n341 4.5
R1193 net6.n332 net6.n330 4.5
R1194 net6.n187 net6.n186 4.5
R1195 net6.n224 net6.n223 4.5
R1196 net6.n205 net6.n196 4.5
R1197 net6.n153 net6.n150 4.5
R1198 net6.n201 net6.n200 4.5
R1199 net6.n80 net6.n79 4.5
R1200 net6.n110 net6.n109 4.5
R1201 net6.n3576 net6.n3574 4.325
R1202 net6.n3215 net6.n3213 4.325
R1203 net6.n2854 net6.n2852 4.325
R1204 net6.n2493 net6.n2491 4.325
R1205 net6.n2132 net6.n2130 4.325
R1206 net6.n1770 net6.n1768 4.325
R1207 net6.n1408 net6.n1406 4.325
R1208 net6.n1046 net6.n1044 4.325
R1209 net6.n684 net6.n682 4.325
R1210 net6.n322 net6.n320 4.325
R1211 net6.n3669 net6.t11 4.289
R1212 net6.n3308 net6.t1 4.289
R1213 net6.n2947 net6.t4 4.289
R1214 net6.n2586 net6.t3 4.289
R1215 net6.n2225 net6.t0 4.289
R1216 net6.n1863 net6.t8 4.289
R1217 net6.n1501 net6.t2 4.289
R1218 net6.n1139 net6.t10 4.289
R1219 net6.n777 net6.t7 4.289
R1220 net6.n415 net6.t9 4.289
R1221 net6.n3580 net6.n3577 3.95
R1222 net6.n3219 net6.n3216 3.95
R1223 net6.n2858 net6.n2855 3.95
R1224 net6.n2497 net6.n2494 3.95
R1225 net6.n2136 net6.n2133 3.95
R1226 net6.n1774 net6.n1771 3.95
R1227 net6.n1412 net6.n1409 3.95
R1228 net6.n1050 net6.n1047 3.95
R1229 net6.n688 net6.n685 3.95
R1230 net6.n326 net6.n323 3.95
R1231 net6.n3333 net6.n3332 3.948
R1232 net6.n2972 net6.n2971 3.948
R1233 net6.n2611 net6.n2610 3.948
R1234 net6.n2250 net6.n2249 3.948
R1235 net6.n1889 net6.n1888 3.948
R1236 net6.n1527 net6.n1526 3.948
R1237 net6.n1165 net6.n1164 3.948
R1238 net6.n803 net6.n802 3.948
R1239 net6.n441 net6.n440 3.948
R1240 net6.n79 net6.n78 3.948
R1241 net6.n3454 net6.n3453 3.573
R1242 net6.n3093 net6.n3092 3.573
R1243 net6.n2732 net6.n2731 3.573
R1244 net6.n2371 net6.n2370 3.573
R1245 net6.n2010 net6.n2009 3.573
R1246 net6.n1648 net6.n1647 3.573
R1247 net6.n1286 net6.n1285 3.573
R1248 net6.n924 net6.n923 3.573
R1249 net6.n562 net6.n561 3.573
R1250 net6.n200 net6.n199 3.573
R1251 net6.n3467 net6.n3448 3.033
R1252 net6.n3342 net6.n3341 3.033
R1253 net6.n3106 net6.n3087 3.033
R1254 net6.n2981 net6.n2980 3.033
R1255 net6.n2745 net6.n2726 3.033
R1256 net6.n2620 net6.n2619 3.033
R1257 net6.n2384 net6.n2365 3.033
R1258 net6.n2259 net6.n2258 3.033
R1259 net6.n2023 net6.n2004 3.033
R1260 net6.n1898 net6.n1897 3.033
R1261 net6.n1661 net6.n1642 3.033
R1262 net6.n1536 net6.n1535 3.033
R1263 net6.n1299 net6.n1280 3.033
R1264 net6.n1174 net6.n1173 3.033
R1265 net6.n937 net6.n918 3.033
R1266 net6.n812 net6.n811 3.033
R1267 net6.n575 net6.n556 3.033
R1268 net6.n450 net6.n449 3.033
R1269 net6.n213 net6.n194 3.033
R1270 net6.n88 net6.n87 3.033
R1271 net6.n3579 net6.n3578 2.258
R1272 net6.n3452 net6.n3451 2.258
R1273 net6.n3218 net6.n3217 2.258
R1274 net6.n3091 net6.n3090 2.258
R1275 net6.n2857 net6.n2856 2.258
R1276 net6.n2730 net6.n2729 2.258
R1277 net6.n2496 net6.n2495 2.258
R1278 net6.n2369 net6.n2368 2.258
R1279 net6.n2135 net6.n2134 2.258
R1280 net6.n2008 net6.n2007 2.258
R1281 net6.n1773 net6.n1772 2.258
R1282 net6.n1646 net6.n1645 2.258
R1283 net6.n1411 net6.n1410 2.258
R1284 net6.n1284 net6.n1283 2.258
R1285 net6.n1049 net6.n1048 2.258
R1286 net6.n922 net6.n921 2.258
R1287 net6.n687 net6.n686 2.258
R1288 net6.n560 net6.n559 2.258
R1289 net6.n325 net6.n324 2.258
R1290 net6.n198 net6.n197 2.258
R1291 net6.n49 net6.n48 2.25
R1292 net6.n3679 net6.n3678 2.07
R1293 net6.n3679 net6.n3317 2.014
R1294 net6.n3681 net6.n2595 2.014
R1295 net6.n1873 net6.n1872 2.014
R1296 net6.n1149 net6.n1148 2.014
R1297 net6.n425 net6.n424 2.014
R1298 net6.n787 net6.n786 2.014
R1299 net6.n1511 net6.n1510 2.014
R1300 net6.n3682 net6.n2234 2.014
R1301 net6.n3680 net6.n2956 2.014
R1302 net6.n3627 net6.n3626 1.882
R1303 net6.n3628 net6.n3627 1.882
R1304 net6.n3403 net6.n3402 1.882
R1305 net6.n3266 net6.n3265 1.882
R1306 net6.n3267 net6.n3266 1.882
R1307 net6.n3042 net6.n3041 1.882
R1308 net6.n2905 net6.n2904 1.882
R1309 net6.n2906 net6.n2905 1.882
R1310 net6.n2681 net6.n2680 1.882
R1311 net6.n2544 net6.n2543 1.882
R1312 net6.n2545 net6.n2544 1.882
R1313 net6.n2320 net6.n2319 1.882
R1314 net6.n2183 net6.n2182 1.882
R1315 net6.n2184 net6.n2183 1.882
R1316 net6.n1959 net6.n1958 1.882
R1317 net6.n1821 net6.n1820 1.882
R1318 net6.n1822 net6.n1821 1.882
R1319 net6.n1597 net6.n1596 1.882
R1320 net6.n1459 net6.n1458 1.882
R1321 net6.n1460 net6.n1459 1.882
R1322 net6.n1235 net6.n1234 1.882
R1323 net6.n1097 net6.n1096 1.882
R1324 net6.n1098 net6.n1097 1.882
R1325 net6.n873 net6.n872 1.882
R1326 net6.n735 net6.n734 1.882
R1327 net6.n736 net6.n735 1.882
R1328 net6.n511 net6.n510 1.882
R1329 net6.n373 net6.n372 1.882
R1330 net6.n374 net6.n373 1.882
R1331 net6.n149 net6.n148 1.882
R1332 net6.n3670 net6.n3669 1.844
R1333 net6.n3309 net6.n3308 1.844
R1334 net6.n2948 net6.n2947 1.844
R1335 net6.n2587 net6.n2586 1.844
R1336 net6.n2226 net6.n2225 1.844
R1337 net6.n1864 net6.n1863 1.844
R1338 net6.n1502 net6.n1501 1.844
R1339 net6.n1140 net6.n1139 1.844
R1340 net6.n778 net6.n777 1.844
R1341 net6.n416 net6.n415 1.844
R1342 net6.n59 net6.n22 1.712
R1343 net6.n12 net6.n11 1.706
R1344 net6.n59 net6.n58 1.701
R1345 net6.n59 net6.n51 1.701
R1346 net6.n3454 net6.n3452 1.505
R1347 net6.n3404 net6.n3403 1.505
R1348 net6.n3093 net6.n3091 1.505
R1349 net6.n3043 net6.n3042 1.505
R1350 net6.n2732 net6.n2730 1.505
R1351 net6.n2682 net6.n2681 1.505
R1352 net6.n2371 net6.n2369 1.505
R1353 net6.n2321 net6.n2320 1.505
R1354 net6.n2010 net6.n2008 1.505
R1355 net6.n1960 net6.n1959 1.505
R1356 net6.n1648 net6.n1646 1.505
R1357 net6.n1598 net6.n1597 1.505
R1358 net6.n1286 net6.n1284 1.505
R1359 net6.n1236 net6.n1235 1.505
R1360 net6.n924 net6.n922 1.505
R1361 net6.n874 net6.n873 1.505
R1362 net6.n562 net6.n560 1.505
R1363 net6.n512 net6.n511 1.505
R1364 net6.n200 net6.n198 1.505
R1365 net6.n150 net6.n149 1.505
R1366 net6.n3430 net6.n3429 1.137
R1367 net6.n3508 net6.n3507 1.137
R1368 net6.n3515 net6.n3514 1.137
R1369 net6.n3519 net6.n3518 1.137
R1370 net6.n3526 net6.n3525 1.137
R1371 net6.n3544 net6.n3543 1.137
R1372 net6.n3561 net6.n3560 1.137
R1373 net6.n3568 net6.n3567 1.137
R1374 net6.n3557 net6.n3556 1.137
R1375 net6.n3550 net6.n3549 1.137
R1376 net6.n3536 net6.n3535 1.137
R1377 net6.n3500 net6.n3499 1.137
R1378 net6.n3491 net6.n3490 1.137
R1379 net6.n3482 net6.n3481 1.137
R1380 net6.n3419 net6.n3418 1.137
R1381 net6.n3426 net6.n3425 1.137
R1382 net6.n3411 net6.n3410 1.137
R1383 net6.n3396 net6.n3395 1.137
R1384 net6.n3380 net6.n3379 1.137
R1385 net6.n3387 net6.n3386 1.137
R1386 net6.n3678 net6.n3677 1.137
R1387 net6.n3069 net6.n3068 1.137
R1388 net6.n3147 net6.n3146 1.137
R1389 net6.n3154 net6.n3153 1.137
R1390 net6.n3158 net6.n3157 1.137
R1391 net6.n3165 net6.n3164 1.137
R1392 net6.n3183 net6.n3182 1.137
R1393 net6.n3200 net6.n3199 1.137
R1394 net6.n3207 net6.n3206 1.137
R1395 net6.n3196 net6.n3195 1.137
R1396 net6.n3189 net6.n3188 1.137
R1397 net6.n3175 net6.n3174 1.137
R1398 net6.n3139 net6.n3138 1.137
R1399 net6.n3130 net6.n3129 1.137
R1400 net6.n3121 net6.n3120 1.137
R1401 net6.n3058 net6.n3057 1.137
R1402 net6.n3065 net6.n3064 1.137
R1403 net6.n3050 net6.n3049 1.137
R1404 net6.n3035 net6.n3034 1.137
R1405 net6.n3019 net6.n3018 1.137
R1406 net6.n3026 net6.n3025 1.137
R1407 net6.n3317 net6.n3316 1.137
R1408 net6.n2708 net6.n2707 1.137
R1409 net6.n2786 net6.n2785 1.137
R1410 net6.n2793 net6.n2792 1.137
R1411 net6.n2797 net6.n2796 1.137
R1412 net6.n2804 net6.n2803 1.137
R1413 net6.n2822 net6.n2821 1.137
R1414 net6.n2839 net6.n2838 1.137
R1415 net6.n2846 net6.n2845 1.137
R1416 net6.n2835 net6.n2834 1.137
R1417 net6.n2828 net6.n2827 1.137
R1418 net6.n2814 net6.n2813 1.137
R1419 net6.n2778 net6.n2777 1.137
R1420 net6.n2769 net6.n2768 1.137
R1421 net6.n2760 net6.n2759 1.137
R1422 net6.n2697 net6.n2696 1.137
R1423 net6.n2704 net6.n2703 1.137
R1424 net6.n2689 net6.n2688 1.137
R1425 net6.n2674 net6.n2673 1.137
R1426 net6.n2658 net6.n2657 1.137
R1427 net6.n2665 net6.n2664 1.137
R1428 net6.n2956 net6.n2955 1.137
R1429 net6.n2347 net6.n2346 1.137
R1430 net6.n2425 net6.n2424 1.137
R1431 net6.n2432 net6.n2431 1.137
R1432 net6.n2436 net6.n2435 1.137
R1433 net6.n2443 net6.n2442 1.137
R1434 net6.n2461 net6.n2460 1.137
R1435 net6.n2478 net6.n2477 1.137
R1436 net6.n2485 net6.n2484 1.137
R1437 net6.n2474 net6.n2473 1.137
R1438 net6.n2467 net6.n2466 1.137
R1439 net6.n2453 net6.n2452 1.137
R1440 net6.n2417 net6.n2416 1.137
R1441 net6.n2408 net6.n2407 1.137
R1442 net6.n2399 net6.n2398 1.137
R1443 net6.n2336 net6.n2335 1.137
R1444 net6.n2343 net6.n2342 1.137
R1445 net6.n2328 net6.n2327 1.137
R1446 net6.n2313 net6.n2312 1.137
R1447 net6.n2297 net6.n2296 1.137
R1448 net6.n2304 net6.n2303 1.137
R1449 net6.n2595 net6.n2594 1.137
R1450 net6.n1986 net6.n1985 1.137
R1451 net6.n2064 net6.n2063 1.137
R1452 net6.n2071 net6.n2070 1.137
R1453 net6.n2075 net6.n2074 1.137
R1454 net6.n2082 net6.n2081 1.137
R1455 net6.n2100 net6.n2099 1.137
R1456 net6.n2117 net6.n2116 1.137
R1457 net6.n2124 net6.n2123 1.137
R1458 net6.n2113 net6.n2112 1.137
R1459 net6.n2106 net6.n2105 1.137
R1460 net6.n2092 net6.n2091 1.137
R1461 net6.n2056 net6.n2055 1.137
R1462 net6.n2047 net6.n2046 1.137
R1463 net6.n2038 net6.n2037 1.137
R1464 net6.n1975 net6.n1974 1.137
R1465 net6.n1982 net6.n1981 1.137
R1466 net6.n1967 net6.n1966 1.137
R1467 net6.n1952 net6.n1951 1.137
R1468 net6.n1936 net6.n1935 1.137
R1469 net6.n1943 net6.n1942 1.137
R1470 net6.n2234 net6.n2233 1.137
R1471 net6.n1624 net6.n1623 1.137
R1472 net6.n1702 net6.n1701 1.137
R1473 net6.n1709 net6.n1708 1.137
R1474 net6.n1713 net6.n1712 1.137
R1475 net6.n1720 net6.n1719 1.137
R1476 net6.n1738 net6.n1737 1.137
R1477 net6.n1755 net6.n1754 1.137
R1478 net6.n1762 net6.n1761 1.137
R1479 net6.n1751 net6.n1750 1.137
R1480 net6.n1744 net6.n1743 1.137
R1481 net6.n1730 net6.n1729 1.137
R1482 net6.n1694 net6.n1693 1.137
R1483 net6.n1685 net6.n1684 1.137
R1484 net6.n1676 net6.n1675 1.137
R1485 net6.n1613 net6.n1612 1.137
R1486 net6.n1620 net6.n1619 1.137
R1487 net6.n1605 net6.n1604 1.137
R1488 net6.n1590 net6.n1589 1.137
R1489 net6.n1574 net6.n1573 1.137
R1490 net6.n1581 net6.n1580 1.137
R1491 net6.n1872 net6.n1871 1.137
R1492 net6.n1262 net6.n1261 1.137
R1493 net6.n1340 net6.n1339 1.137
R1494 net6.n1347 net6.n1346 1.137
R1495 net6.n1351 net6.n1350 1.137
R1496 net6.n1358 net6.n1357 1.137
R1497 net6.n1376 net6.n1375 1.137
R1498 net6.n1393 net6.n1392 1.137
R1499 net6.n1400 net6.n1399 1.137
R1500 net6.n1389 net6.n1388 1.137
R1501 net6.n1382 net6.n1381 1.137
R1502 net6.n1368 net6.n1367 1.137
R1503 net6.n1332 net6.n1331 1.137
R1504 net6.n1323 net6.n1322 1.137
R1505 net6.n1314 net6.n1313 1.137
R1506 net6.n1251 net6.n1250 1.137
R1507 net6.n1258 net6.n1257 1.137
R1508 net6.n1243 net6.n1242 1.137
R1509 net6.n1228 net6.n1227 1.137
R1510 net6.n1212 net6.n1211 1.137
R1511 net6.n1219 net6.n1218 1.137
R1512 net6.n1510 net6.n1509 1.137
R1513 net6.n900 net6.n899 1.137
R1514 net6.n978 net6.n977 1.137
R1515 net6.n985 net6.n984 1.137
R1516 net6.n989 net6.n988 1.137
R1517 net6.n996 net6.n995 1.137
R1518 net6.n1014 net6.n1013 1.137
R1519 net6.n1031 net6.n1030 1.137
R1520 net6.n1038 net6.n1037 1.137
R1521 net6.n1027 net6.n1026 1.137
R1522 net6.n1020 net6.n1019 1.137
R1523 net6.n1006 net6.n1005 1.137
R1524 net6.n970 net6.n969 1.137
R1525 net6.n961 net6.n960 1.137
R1526 net6.n952 net6.n951 1.137
R1527 net6.n889 net6.n888 1.137
R1528 net6.n896 net6.n895 1.137
R1529 net6.n881 net6.n880 1.137
R1530 net6.n866 net6.n865 1.137
R1531 net6.n850 net6.n849 1.137
R1532 net6.n857 net6.n856 1.137
R1533 net6.n1148 net6.n1147 1.137
R1534 net6.n538 net6.n537 1.137
R1535 net6.n616 net6.n615 1.137
R1536 net6.n623 net6.n622 1.137
R1537 net6.n627 net6.n626 1.137
R1538 net6.n634 net6.n633 1.137
R1539 net6.n652 net6.n651 1.137
R1540 net6.n669 net6.n668 1.137
R1541 net6.n676 net6.n675 1.137
R1542 net6.n665 net6.n664 1.137
R1543 net6.n658 net6.n657 1.137
R1544 net6.n644 net6.n643 1.137
R1545 net6.n608 net6.n607 1.137
R1546 net6.n599 net6.n598 1.137
R1547 net6.n590 net6.n589 1.137
R1548 net6.n527 net6.n526 1.137
R1549 net6.n534 net6.n533 1.137
R1550 net6.n519 net6.n518 1.137
R1551 net6.n504 net6.n503 1.137
R1552 net6.n488 net6.n487 1.137
R1553 net6.n495 net6.n494 1.137
R1554 net6.n786 net6.n785 1.137
R1555 net6.n176 net6.n175 1.137
R1556 net6.n254 net6.n253 1.137
R1557 net6.n261 net6.n260 1.137
R1558 net6.n265 net6.n264 1.137
R1559 net6.n272 net6.n271 1.137
R1560 net6.n290 net6.n289 1.137
R1561 net6.n307 net6.n306 1.137
R1562 net6.n314 net6.n313 1.137
R1563 net6.n303 net6.n302 1.137
R1564 net6.n296 net6.n295 1.137
R1565 net6.n282 net6.n281 1.137
R1566 net6.n246 net6.n245 1.137
R1567 net6.n237 net6.n236 1.137
R1568 net6.n228 net6.n227 1.137
R1569 net6.n165 net6.n164 1.137
R1570 net6.n172 net6.n171 1.137
R1571 net6.n157 net6.n156 1.137
R1572 net6.n142 net6.n141 1.137
R1573 net6.n126 net6.n125 1.137
R1574 net6.n133 net6.n132 1.137
R1575 net6.n424 net6.n423 1.137
R1576 net6.n3573 net6.n3572 1.129
R1577 net6.n3580 net6.n3579 1.129
R1578 net6.n3618 net6.n3617 1.129
R1579 net6.n3212 net6.n3211 1.129
R1580 net6.n3219 net6.n3218 1.129
R1581 net6.n3257 net6.n3256 1.129
R1582 net6.n2851 net6.n2850 1.129
R1583 net6.n2858 net6.n2857 1.129
R1584 net6.n2896 net6.n2895 1.129
R1585 net6.n2490 net6.n2489 1.129
R1586 net6.n2497 net6.n2496 1.129
R1587 net6.n2535 net6.n2534 1.129
R1588 net6.n2129 net6.n2128 1.129
R1589 net6.n2136 net6.n2135 1.129
R1590 net6.n2174 net6.n2173 1.129
R1591 net6.n1767 net6.n1766 1.129
R1592 net6.n1774 net6.n1773 1.129
R1593 net6.n1812 net6.n1811 1.129
R1594 net6.n1405 net6.n1404 1.129
R1595 net6.n1412 net6.n1411 1.129
R1596 net6.n1450 net6.n1449 1.129
R1597 net6.n1043 net6.n1042 1.129
R1598 net6.n1050 net6.n1049 1.129
R1599 net6.n1088 net6.n1087 1.129
R1600 net6.n681 net6.n680 1.129
R1601 net6.n688 net6.n687 1.129
R1602 net6.n726 net6.n725 1.129
R1603 net6.n319 net6.n318 1.129
R1604 net6.n326 net6.n325 1.129
R1605 net6.n364 net6.n363 1.129
R1606 net6.n3408 net6.n3407 1.125
R1607 net6.n3047 net6.n3046 1.125
R1608 net6.n2686 net6.n2685 1.125
R1609 net6.n2325 net6.n2324 1.125
R1610 net6.n1964 net6.n1963 1.125
R1611 net6.n1602 net6.n1601 1.125
R1612 net6.n1240 net6.n1239 1.125
R1613 net6.n878 net6.n877 1.125
R1614 net6.n516 net6.n515 1.125
R1615 net6.n154 net6.n153 1.125
R1616 net6.n425 net6.n63 1.079
R1617 net6.n3481 net6.n3478 1.042
R1618 net6.n3120 net6.n3117 1.042
R1619 net6.n2759 net6.n2756 1.042
R1620 net6.n2398 net6.n2395 1.042
R1621 net6.n2037 net6.n2034 1.042
R1622 net6.n1675 net6.n1672 1.042
R1623 net6.n1313 net6.n1310 1.042
R1624 net6.n951 net6.n948 1.042
R1625 net6.n589 net6.n586 1.042
R1626 net6.n227 net6.n224 1.042
R1627 net6.n3372 net6.n3371 0.869
R1628 net6.n3011 net6.n3010 0.869
R1629 net6.n2650 net6.n2649 0.869
R1630 net6.n2289 net6.n2288 0.869
R1631 net6.n1928 net6.n1927 0.869
R1632 net6.n1566 net6.n1565 0.869
R1633 net6.n1204 net6.n1203 0.869
R1634 net6.n842 net6.n841 0.869
R1635 net6.n480 net6.n479 0.869
R1636 net6.n118 net6.n117 0.869
R1637 net6.n3663 net6.n3662 0.752
R1638 net6.n3477 net6.n3476 0.752
R1639 net6.n3450 net6.n3449 0.752
R1640 net6.n3333 net6.n3331 0.752
R1641 net6.n3352 net6.n3351 0.752
R1642 net6.n3363 net6.n3362 0.752
R1643 net6.n3302 net6.n3301 0.752
R1644 net6.n3116 net6.n3115 0.752
R1645 net6.n3089 net6.n3088 0.752
R1646 net6.n2972 net6.n2970 0.752
R1647 net6.n2991 net6.n2990 0.752
R1648 net6.n3002 net6.n3001 0.752
R1649 net6.n2941 net6.n2940 0.752
R1650 net6.n2755 net6.n2754 0.752
R1651 net6.n2728 net6.n2727 0.752
R1652 net6.n2611 net6.n2609 0.752
R1653 net6.n2630 net6.n2629 0.752
R1654 net6.n2641 net6.n2640 0.752
R1655 net6.n2580 net6.n2579 0.752
R1656 net6.n2394 net6.n2393 0.752
R1657 net6.n2367 net6.n2366 0.752
R1658 net6.n2250 net6.n2248 0.752
R1659 net6.n2269 net6.n2268 0.752
R1660 net6.n2280 net6.n2279 0.752
R1661 net6.n2219 net6.n2218 0.752
R1662 net6.n2033 net6.n2032 0.752
R1663 net6.n2006 net6.n2005 0.752
R1664 net6.n1889 net6.n1887 0.752
R1665 net6.n1908 net6.n1907 0.752
R1666 net6.n1919 net6.n1918 0.752
R1667 net6.n1857 net6.n1856 0.752
R1668 net6.n1671 net6.n1670 0.752
R1669 net6.n1644 net6.n1643 0.752
R1670 net6.n1527 net6.n1525 0.752
R1671 net6.n1546 net6.n1545 0.752
R1672 net6.n1557 net6.n1556 0.752
R1673 net6.n1495 net6.n1494 0.752
R1674 net6.n1309 net6.n1308 0.752
R1675 net6.n1282 net6.n1281 0.752
R1676 net6.n1165 net6.n1163 0.752
R1677 net6.n1184 net6.n1183 0.752
R1678 net6.n1195 net6.n1194 0.752
R1679 net6.n1133 net6.n1132 0.752
R1680 net6.n947 net6.n946 0.752
R1681 net6.n920 net6.n919 0.752
R1682 net6.n803 net6.n801 0.752
R1683 net6.n822 net6.n821 0.752
R1684 net6.n833 net6.n832 0.752
R1685 net6.n771 net6.n770 0.752
R1686 net6.n585 net6.n584 0.752
R1687 net6.n558 net6.n557 0.752
R1688 net6.n441 net6.n439 0.752
R1689 net6.n460 net6.n459 0.752
R1690 net6.n471 net6.n470 0.752
R1691 net6.n409 net6.n408 0.752
R1692 net6.n223 net6.n222 0.752
R1693 net6.n196 net6.n195 0.752
R1694 net6.n79 net6.n77 0.752
R1695 net6.n98 net6.n97 0.752
R1696 net6.n109 net6.n108 0.752
R1697 net6.n3371 net6.n3370 0.728
R1698 net6.n3010 net6.n3009 0.728
R1699 net6.n2649 net6.n2648 0.728
R1700 net6.n2288 net6.n2287 0.728
R1701 net6.n1927 net6.n1926 0.728
R1702 net6.n1565 net6.n1564 0.728
R1703 net6.n1203 net6.n1202 0.728
R1704 net6.n841 net6.n840 0.728
R1705 net6.n479 net6.n478 0.728
R1706 net6.n117 net6.n116 0.728
R1707 net6.n3677 net6.n3671 0.725
R1708 net6.n3316 net6.n3310 0.725
R1709 net6.n2955 net6.n2949 0.725
R1710 net6.n2594 net6.n2588 0.725
R1711 net6.n2233 net6.n2227 0.725
R1712 net6.n1871 net6.n1865 0.725
R1713 net6.n1509 net6.n1503 0.725
R1714 net6.n1147 net6.n1141 0.725
R1715 net6.n785 net6.n779 0.725
R1716 net6.n423 net6.n417 0.725
R1717 net6.n3644 net6.n3643 0.376
R1718 net6.n3576 net6.n3575 0.376
R1719 net6.n3582 net6.n3581 0.376
R1720 net6.n3595 net6.n3594 0.376
R1721 net6.n3584 net6.n3583 0.376
R1722 net6.n3440 net6.n3439 0.376
R1723 net6.n3283 net6.n3282 0.376
R1724 net6.n3215 net6.n3214 0.376
R1725 net6.n3221 net6.n3220 0.376
R1726 net6.n3234 net6.n3233 0.376
R1727 net6.n3223 net6.n3222 0.376
R1728 net6.n3079 net6.n3078 0.376
R1729 net6.n2922 net6.n2921 0.376
R1730 net6.n2854 net6.n2853 0.376
R1731 net6.n2860 net6.n2859 0.376
R1732 net6.n2873 net6.n2872 0.376
R1733 net6.n2862 net6.n2861 0.376
R1734 net6.n2718 net6.n2717 0.376
R1735 net6.n2561 net6.n2560 0.376
R1736 net6.n2493 net6.n2492 0.376
R1737 net6.n2499 net6.n2498 0.376
R1738 net6.n2512 net6.n2511 0.376
R1739 net6.n2501 net6.n2500 0.376
R1740 net6.n2357 net6.n2356 0.376
R1741 net6.n2200 net6.n2199 0.376
R1742 net6.n2132 net6.n2131 0.376
R1743 net6.n2138 net6.n2137 0.376
R1744 net6.n2151 net6.n2150 0.376
R1745 net6.n2140 net6.n2139 0.376
R1746 net6.n1996 net6.n1995 0.376
R1747 net6.n1838 net6.n1837 0.376
R1748 net6.n1770 net6.n1769 0.376
R1749 net6.n1776 net6.n1775 0.376
R1750 net6.n1789 net6.n1788 0.376
R1751 net6.n1778 net6.n1777 0.376
R1752 net6.n1634 net6.n1633 0.376
R1753 net6.n1476 net6.n1475 0.376
R1754 net6.n1408 net6.n1407 0.376
R1755 net6.n1414 net6.n1413 0.376
R1756 net6.n1427 net6.n1426 0.376
R1757 net6.n1416 net6.n1415 0.376
R1758 net6.n1272 net6.n1271 0.376
R1759 net6.n1114 net6.n1113 0.376
R1760 net6.n1046 net6.n1045 0.376
R1761 net6.n1052 net6.n1051 0.376
R1762 net6.n1065 net6.n1064 0.376
R1763 net6.n1054 net6.n1053 0.376
R1764 net6.n910 net6.n909 0.376
R1765 net6.n752 net6.n751 0.376
R1766 net6.n684 net6.n683 0.376
R1767 net6.n690 net6.n689 0.376
R1768 net6.n703 net6.n702 0.376
R1769 net6.n692 net6.n691 0.376
R1770 net6.n548 net6.n547 0.376
R1771 net6.n390 net6.n389 0.376
R1772 net6.n322 net6.n321 0.376
R1773 net6.n328 net6.n327 0.376
R1774 net6.n341 net6.n340 0.376
R1775 net6.n330 net6.n329 0.376
R1776 net6.n186 net6.n185 0.376
R1777 net6.n3443 net6.n3442 0.189
R1778 net6.n3082 net6.n3081 0.189
R1779 net6.n2721 net6.n2720 0.189
R1780 net6.n2360 net6.n2359 0.189
R1781 net6.n1999 net6.n1998 0.189
R1782 net6.n1637 net6.n1636 0.189
R1783 net6.n1275 net6.n1274 0.189
R1784 net6.n913 net6.n912 0.189
R1785 net6.n551 net6.n550 0.189
R1786 net6.n189 net6.n188 0.189
R1787 net6.n3588 net6.n3587 0.188
R1788 net6.n3227 net6.n3226 0.188
R1789 net6.n2866 net6.n2865 0.188
R1790 net6.n2505 net6.n2504 0.188
R1791 net6.n2144 net6.n2143 0.188
R1792 net6.n1782 net6.n1781 0.188
R1793 net6.n1420 net6.n1419 0.188
R1794 net6.n1058 net6.n1057 0.188
R1795 net6.n696 net6.n695 0.188
R1796 net6.n334 net6.n333 0.188
R1797 net6.n61 net6.n2 0.182
R1798 net6.n3464 net6.n3463 0.166
R1799 net6.n3103 net6.n3102 0.166
R1800 net6.n2742 net6.n2741 0.166
R1801 net6.n2381 net6.n2380 0.166
R1802 net6.n2020 net6.n2019 0.166
R1803 net6.n1658 net6.n1657 0.166
R1804 net6.n1296 net6.n1295 0.166
R1805 net6.n934 net6.n933 0.166
R1806 net6.n572 net6.n571 0.166
R1807 net6.n210 net6.n209 0.166
R1808 net6.n3612 net6.n3611 0.166
R1809 net6.n3251 net6.n3250 0.166
R1810 net6.n2890 net6.n2889 0.166
R1811 net6.n2529 net6.n2528 0.166
R1812 net6.n2168 net6.n2167 0.166
R1813 net6.n1806 net6.n1805 0.166
R1814 net6.n1444 net6.n1443 0.166
R1815 net6.n1082 net6.n1081 0.166
R1816 net6.n720 net6.n719 0.166
R1817 net6.n358 net6.n357 0.166
R1818 net6.n3341 net6.n3340 0.133
R1819 net6.n2980 net6.n2979 0.133
R1820 net6.n2619 net6.n2618 0.133
R1821 net6.n2258 net6.n2257 0.133
R1822 net6.n1897 net6.n1896 0.133
R1823 net6.n1535 net6.n1534 0.133
R1824 net6.n1173 net6.n1172 0.133
R1825 net6.n811 net6.n810 0.133
R1826 net6.n449 net6.n448 0.133
R1827 net6.n87 net6.n86 0.133
R1828 net6.n3643 net6.n3642 0.132
R1829 net6.n3282 net6.n3281 0.132
R1830 net6.n2921 net6.n2920 0.132
R1831 net6.n2560 net6.n2559 0.132
R1832 net6.n2199 net6.n2198 0.132
R1833 net6.n1837 net6.n1836 0.132
R1834 net6.n1475 net6.n1474 0.132
R1835 net6.n1113 net6.n1112 0.132
R1836 net6.n751 net6.n750 0.132
R1837 net6.n389 net6.n388 0.132
R1838 net6.n3351 net6.n3350 0.121
R1839 net6.n2990 net6.n2989 0.121
R1840 net6.n2629 net6.n2628 0.121
R1841 net6.n2268 net6.n2267 0.121
R1842 net6.n1907 net6.n1906 0.121
R1843 net6.n1545 net6.n1544 0.121
R1844 net6.n1183 net6.n1182 0.121
R1845 net6.n821 net6.n820 0.121
R1846 net6.n459 net6.n458 0.121
R1847 net6.n97 net6.n96 0.121
R1848 net6.n3572 net6.n3571 0.121
R1849 net6.n3211 net6.n3210 0.121
R1850 net6.n2850 net6.n2849 0.121
R1851 net6.n2489 net6.n2488 0.121
R1852 net6.n2128 net6.n2127 0.121
R1853 net6.n1766 net6.n1765 0.121
R1854 net6.n1404 net6.n1403 0.121
R1855 net6.n1042 net6.n1041 0.121
R1856 net6.n680 net6.n679 0.121
R1857 net6.n318 net6.n317 0.121
R1858 net6.n1511 net6.n1149 0.116
R1859 net6.n3681 net6.n3680 0.116
R1860 net6 net6.n1873 0.097
R1861 net6.n2 net6.n1 0.089
R1862 net6.n34 net6.n33 0.071
R1863 net6.n44 net6.n43 0.071
R1864 net6.n787 net6.n425 0.058
R1865 net6.n1149 net6.n787 0.058
R1866 net6.n1873 net6.n1511 0.058
R1867 net6.n3682 net6.n3681 0.058
R1868 net6.n3680 net6.n3679 0.058
R1869 net6.n37 net6.n36 0.053
R1870 net6.n47 net6.n46 0.053
R1871 net6.n3549 net6.n3548 0.049
R1872 net6.n3544 net6.n3536 0.049
R1873 net6.n3500 net6.n3491 0.049
R1874 net6.n3411 net6.n3396 0.049
R1875 net6.n3188 net6.n3187 0.049
R1876 net6.n3183 net6.n3175 0.049
R1877 net6.n3139 net6.n3130 0.049
R1878 net6.n3050 net6.n3035 0.049
R1879 net6.n2827 net6.n2826 0.049
R1880 net6.n2822 net6.n2814 0.049
R1881 net6.n2778 net6.n2769 0.049
R1882 net6.n2689 net6.n2674 0.049
R1883 net6.n2466 net6.n2465 0.049
R1884 net6.n2461 net6.n2453 0.049
R1885 net6.n2417 net6.n2408 0.049
R1886 net6.n2328 net6.n2313 0.049
R1887 net6.n2105 net6.n2104 0.049
R1888 net6.n2100 net6.n2092 0.049
R1889 net6.n2056 net6.n2047 0.049
R1890 net6.n1967 net6.n1952 0.049
R1891 net6.n1743 net6.n1742 0.049
R1892 net6.n1738 net6.n1730 0.049
R1893 net6.n1694 net6.n1685 0.049
R1894 net6.n1605 net6.n1590 0.049
R1895 net6.n1381 net6.n1380 0.049
R1896 net6.n1376 net6.n1368 0.049
R1897 net6.n1332 net6.n1323 0.049
R1898 net6.n1243 net6.n1228 0.049
R1899 net6.n1019 net6.n1018 0.049
R1900 net6.n1014 net6.n1006 0.049
R1901 net6.n970 net6.n961 0.049
R1902 net6.n881 net6.n866 0.049
R1903 net6.n657 net6.n656 0.049
R1904 net6.n652 net6.n644 0.049
R1905 net6.n608 net6.n599 0.049
R1906 net6.n519 net6.n504 0.049
R1907 net6.n295 net6.n294 0.049
R1908 net6.n290 net6.n282 0.049
R1909 net6.n246 net6.n237 0.049
R1910 net6.n157 net6.n142 0.049
R1911 net6.n3668 net6.n3667 0.047
R1912 net6.n3649 net6.n3647 0.047
R1913 net6.n3647 net6.n3646 0.047
R1914 net6.n3639 net6.n3637 0.047
R1915 net6.n3591 net6.n3590 0.047
R1916 net6.n3446 net6.n3445 0.047
R1917 net6.n3338 net6.n3336 0.047
R1918 net6.n3343 net6.n3342 0.047
R1919 net6.n3346 net6.n3344 0.047
R1920 net6.n3368 net6.n3367 0.047
R1921 net6.n3506 net6.n3505 0.047
R1922 net6.n3307 net6.n3306 0.047
R1923 net6.n3288 net6.n3286 0.047
R1924 net6.n3286 net6.n3285 0.047
R1925 net6.n3278 net6.n3276 0.047
R1926 net6.n3230 net6.n3229 0.047
R1927 net6.n3085 net6.n3084 0.047
R1928 net6.n2977 net6.n2975 0.047
R1929 net6.n2982 net6.n2981 0.047
R1930 net6.n2985 net6.n2983 0.047
R1931 net6.n3007 net6.n3006 0.047
R1932 net6.n3145 net6.n3144 0.047
R1933 net6.n2946 net6.n2945 0.047
R1934 net6.n2927 net6.n2925 0.047
R1935 net6.n2925 net6.n2924 0.047
R1936 net6.n2917 net6.n2915 0.047
R1937 net6.n2869 net6.n2868 0.047
R1938 net6.n2724 net6.n2723 0.047
R1939 net6.n2616 net6.n2614 0.047
R1940 net6.n2621 net6.n2620 0.047
R1941 net6.n2624 net6.n2622 0.047
R1942 net6.n2646 net6.n2645 0.047
R1943 net6.n2784 net6.n2783 0.047
R1944 net6.n2585 net6.n2584 0.047
R1945 net6.n2566 net6.n2564 0.047
R1946 net6.n2564 net6.n2563 0.047
R1947 net6.n2556 net6.n2554 0.047
R1948 net6.n2508 net6.n2507 0.047
R1949 net6.n2363 net6.n2362 0.047
R1950 net6.n2255 net6.n2253 0.047
R1951 net6.n2260 net6.n2259 0.047
R1952 net6.n2263 net6.n2261 0.047
R1953 net6.n2285 net6.n2284 0.047
R1954 net6.n2423 net6.n2422 0.047
R1955 net6.n2224 net6.n2223 0.047
R1956 net6.n2205 net6.n2203 0.047
R1957 net6.n2203 net6.n2202 0.047
R1958 net6.n2195 net6.n2193 0.047
R1959 net6.n2147 net6.n2146 0.047
R1960 net6.n2002 net6.n2001 0.047
R1961 net6.n1894 net6.n1892 0.047
R1962 net6.n1899 net6.n1898 0.047
R1963 net6.n1902 net6.n1900 0.047
R1964 net6.n1924 net6.n1923 0.047
R1965 net6.n2062 net6.n2061 0.047
R1966 net6.n1862 net6.n1861 0.047
R1967 net6.n1843 net6.n1841 0.047
R1968 net6.n1841 net6.n1840 0.047
R1969 net6.n1833 net6.n1831 0.047
R1970 net6.n1785 net6.n1784 0.047
R1971 net6.n1640 net6.n1639 0.047
R1972 net6.n1532 net6.n1530 0.047
R1973 net6.n1537 net6.n1536 0.047
R1974 net6.n1540 net6.n1538 0.047
R1975 net6.n1562 net6.n1561 0.047
R1976 net6.n1700 net6.n1699 0.047
R1977 net6.n1500 net6.n1499 0.047
R1978 net6.n1481 net6.n1479 0.047
R1979 net6.n1479 net6.n1478 0.047
R1980 net6.n1471 net6.n1469 0.047
R1981 net6.n1423 net6.n1422 0.047
R1982 net6.n1278 net6.n1277 0.047
R1983 net6.n1170 net6.n1168 0.047
R1984 net6.n1175 net6.n1174 0.047
R1985 net6.n1178 net6.n1176 0.047
R1986 net6.n1200 net6.n1199 0.047
R1987 net6.n1338 net6.n1337 0.047
R1988 net6.n1138 net6.n1137 0.047
R1989 net6.n1119 net6.n1117 0.047
R1990 net6.n1117 net6.n1116 0.047
R1991 net6.n1109 net6.n1107 0.047
R1992 net6.n1061 net6.n1060 0.047
R1993 net6.n916 net6.n915 0.047
R1994 net6.n808 net6.n806 0.047
R1995 net6.n813 net6.n812 0.047
R1996 net6.n816 net6.n814 0.047
R1997 net6.n838 net6.n837 0.047
R1998 net6.n976 net6.n975 0.047
R1999 net6.n776 net6.n775 0.047
R2000 net6.n757 net6.n755 0.047
R2001 net6.n755 net6.n754 0.047
R2002 net6.n747 net6.n745 0.047
R2003 net6.n699 net6.n698 0.047
R2004 net6.n554 net6.n553 0.047
R2005 net6.n446 net6.n444 0.047
R2006 net6.n451 net6.n450 0.047
R2007 net6.n454 net6.n452 0.047
R2008 net6.n476 net6.n475 0.047
R2009 net6.n614 net6.n613 0.047
R2010 net6.n414 net6.n413 0.047
R2011 net6.n395 net6.n393 0.047
R2012 net6.n393 net6.n392 0.047
R2013 net6.n385 net6.n383 0.047
R2014 net6.n337 net6.n336 0.047
R2015 net6.n192 net6.n191 0.047
R2016 net6.n84 net6.n82 0.047
R2017 net6.n89 net6.n88 0.047
R2018 net6.n92 net6.n90 0.047
R2019 net6.n114 net6.n113 0.047
R2020 net6.n252 net6.n251 0.047
R2021 net6.n1 net6.n0 0.045
R2022 net6.n3593 net6.n3592 0.045
R2023 net6.n3447 net6.n3446 0.045
R2024 net6.n3232 net6.n3231 0.045
R2025 net6.n3086 net6.n3085 0.045
R2026 net6.n2871 net6.n2870 0.045
R2027 net6.n2725 net6.n2724 0.045
R2028 net6.n2510 net6.n2509 0.045
R2029 net6.n2364 net6.n2363 0.045
R2030 net6.n2149 net6.n2148 0.045
R2031 net6.n2003 net6.n2002 0.045
R2032 net6.n1787 net6.n1786 0.045
R2033 net6.n1641 net6.n1640 0.045
R2034 net6.n1425 net6.n1424 0.045
R2035 net6.n1279 net6.n1278 0.045
R2036 net6.n1063 net6.n1062 0.045
R2037 net6.n917 net6.n916 0.045
R2038 net6.n701 net6.n700 0.045
R2039 net6.n555 net6.n554 0.045
R2040 net6.n339 net6.n338 0.045
R2041 net6.n193 net6.n192 0.045
R2042 net6.n3616 net6.n3615 0.043
R2043 net6.n3407 net6.n3401 0.043
R2044 net6.n3499 net6.n3498 0.043
R2045 net6.n3409 net6.n3408 0.043
R2046 net6.n3394 net6.n3393 0.043
R2047 net6.n3255 net6.n3254 0.043
R2048 net6.n3046 net6.n3040 0.043
R2049 net6.n3138 net6.n3137 0.043
R2050 net6.n3048 net6.n3047 0.043
R2051 net6.n3033 net6.n3032 0.043
R2052 net6.n2894 net6.n2893 0.043
R2053 net6.n2685 net6.n2679 0.043
R2054 net6.n2777 net6.n2776 0.043
R2055 net6.n2687 net6.n2686 0.043
R2056 net6.n2672 net6.n2671 0.043
R2057 net6.n2533 net6.n2532 0.043
R2058 net6.n2324 net6.n2318 0.043
R2059 net6.n2416 net6.n2415 0.043
R2060 net6.n2326 net6.n2325 0.043
R2061 net6.n2311 net6.n2310 0.043
R2062 net6.n2172 net6.n2171 0.043
R2063 net6.n1963 net6.n1957 0.043
R2064 net6.n2055 net6.n2054 0.043
R2065 net6.n1965 net6.n1964 0.043
R2066 net6.n1950 net6.n1949 0.043
R2067 net6.n1810 net6.n1809 0.043
R2068 net6.n1601 net6.n1595 0.043
R2069 net6.n1693 net6.n1692 0.043
R2070 net6.n1603 net6.n1602 0.043
R2071 net6.n1588 net6.n1587 0.043
R2072 net6.n1448 net6.n1447 0.043
R2073 net6.n1239 net6.n1233 0.043
R2074 net6.n1331 net6.n1330 0.043
R2075 net6.n1241 net6.n1240 0.043
R2076 net6.n1226 net6.n1225 0.043
R2077 net6.n1086 net6.n1085 0.043
R2078 net6.n877 net6.n871 0.043
R2079 net6.n969 net6.n968 0.043
R2080 net6.n879 net6.n878 0.043
R2081 net6.n864 net6.n863 0.043
R2082 net6.n724 net6.n723 0.043
R2083 net6.n515 net6.n509 0.043
R2084 net6.n607 net6.n606 0.043
R2085 net6.n517 net6.n516 0.043
R2086 net6.n502 net6.n501 0.043
R2087 net6.n362 net6.n361 0.043
R2088 net6.n153 net6.n147 0.043
R2089 net6.n245 net6.n244 0.043
R2090 net6.n155 net6.n154 0.043
R2091 net6.n140 net6.n139 0.043
R2092 net6.n3671 net6.n3668 0.043
R2093 net6.n3310 net6.n3307 0.043
R2094 net6.n2949 net6.n2946 0.043
R2095 net6.n2588 net6.n2585 0.043
R2096 net6.n2227 net6.n2224 0.043
R2097 net6.n1865 net6.n1862 0.043
R2098 net6.n1503 net6.n1500 0.043
R2099 net6.n1141 net6.n1138 0.043
R2100 net6.n779 net6.n776 0.043
R2101 net6.n417 net6.n414 0.043
R2102 net6.n3636 net6.n3635 0.041
R2103 net6.n3629 net6.n3625 0.041
R2104 net6.n3437 net6.n3436 0.041
R2105 net6.n3461 net6.n3460 0.041
R2106 net6.n3358 net6.n3357 0.041
R2107 net6.n3543 net6.n3542 0.041
R2108 net6.n3417 net6.n3416 0.041
R2109 net6.n3275 net6.n3274 0.041
R2110 net6.n3268 net6.n3264 0.041
R2111 net6.n3076 net6.n3075 0.041
R2112 net6.n3100 net6.n3099 0.041
R2113 net6.n2997 net6.n2996 0.041
R2114 net6.n3182 net6.n3181 0.041
R2115 net6.n3056 net6.n3055 0.041
R2116 net6.n2914 net6.n2913 0.041
R2117 net6.n2907 net6.n2903 0.041
R2118 net6.n2715 net6.n2714 0.041
R2119 net6.n2739 net6.n2738 0.041
R2120 net6.n2636 net6.n2635 0.041
R2121 net6.n2821 net6.n2820 0.041
R2122 net6.n2695 net6.n2694 0.041
R2123 net6.n2553 net6.n2552 0.041
R2124 net6.n2546 net6.n2542 0.041
R2125 net6.n2354 net6.n2353 0.041
R2126 net6.n2378 net6.n2377 0.041
R2127 net6.n2275 net6.n2274 0.041
R2128 net6.n2460 net6.n2459 0.041
R2129 net6.n2334 net6.n2333 0.041
R2130 net6.n2192 net6.n2191 0.041
R2131 net6.n2185 net6.n2181 0.041
R2132 net6.n1993 net6.n1992 0.041
R2133 net6.n2017 net6.n2016 0.041
R2134 net6.n1914 net6.n1913 0.041
R2135 net6.n2099 net6.n2098 0.041
R2136 net6.n1973 net6.n1972 0.041
R2137 net6.n1830 net6.n1829 0.041
R2138 net6.n1823 net6.n1819 0.041
R2139 net6.n1631 net6.n1630 0.041
R2140 net6.n1655 net6.n1654 0.041
R2141 net6.n1552 net6.n1551 0.041
R2142 net6.n1737 net6.n1736 0.041
R2143 net6.n1611 net6.n1610 0.041
R2144 net6.n1468 net6.n1467 0.041
R2145 net6.n1461 net6.n1457 0.041
R2146 net6.n1269 net6.n1268 0.041
R2147 net6.n1293 net6.n1292 0.041
R2148 net6.n1190 net6.n1189 0.041
R2149 net6.n1375 net6.n1374 0.041
R2150 net6.n1249 net6.n1248 0.041
R2151 net6.n1106 net6.n1105 0.041
R2152 net6.n1099 net6.n1095 0.041
R2153 net6.n907 net6.n906 0.041
R2154 net6.n931 net6.n930 0.041
R2155 net6.n828 net6.n827 0.041
R2156 net6.n1013 net6.n1012 0.041
R2157 net6.n887 net6.n886 0.041
R2158 net6.n744 net6.n743 0.041
R2159 net6.n737 net6.n733 0.041
R2160 net6.n545 net6.n544 0.041
R2161 net6.n569 net6.n568 0.041
R2162 net6.n466 net6.n465 0.041
R2163 net6.n651 net6.n650 0.041
R2164 net6.n525 net6.n524 0.041
R2165 net6.n382 net6.n381 0.041
R2166 net6.n375 net6.n371 0.041
R2167 net6.n183 net6.n182 0.041
R2168 net6.n207 net6.n206 0.041
R2169 net6.n104 net6.n103 0.041
R2170 net6.n289 net6.n288 0.041
R2171 net6.n163 net6.n162 0.041
R2172 net6.n3370 net6.n3368 0.041
R2173 net6.n3009 net6.n3007 0.041
R2174 net6.n2648 net6.n2646 0.041
R2175 net6.n2287 net6.n2285 0.041
R2176 net6.n1926 net6.n1924 0.041
R2177 net6.n1564 net6.n1562 0.041
R2178 net6.n1202 net6.n1200 0.041
R2179 net6.n840 net6.n838 0.041
R2180 net6.n478 net6.n476 0.041
R2181 net6.n116 net6.n114 0.041
R2182 net6.n3658 net6.n3657 0.039
R2183 net6.n3614 net6.n3613 0.039
R2184 net6.n3465 net6.n3462 0.039
R2185 net6.n3335 net6.n3334 0.039
R2186 net6.n3395 net6.n3390 0.039
R2187 net6.n3297 net6.n3296 0.039
R2188 net6.n3253 net6.n3252 0.039
R2189 net6.n3104 net6.n3101 0.039
R2190 net6.n2974 net6.n2973 0.039
R2191 net6.n3034 net6.n3029 0.039
R2192 net6.n2936 net6.n2935 0.039
R2193 net6.n2892 net6.n2891 0.039
R2194 net6.n2743 net6.n2740 0.039
R2195 net6.n2613 net6.n2612 0.039
R2196 net6.n2673 net6.n2668 0.039
R2197 net6.n2575 net6.n2574 0.039
R2198 net6.n2531 net6.n2530 0.039
R2199 net6.n2382 net6.n2379 0.039
R2200 net6.n2252 net6.n2251 0.039
R2201 net6.n2312 net6.n2307 0.039
R2202 net6.n2214 net6.n2213 0.039
R2203 net6.n2170 net6.n2169 0.039
R2204 net6.n2021 net6.n2018 0.039
R2205 net6.n1891 net6.n1890 0.039
R2206 net6.n1951 net6.n1946 0.039
R2207 net6.n1852 net6.n1851 0.039
R2208 net6.n1808 net6.n1807 0.039
R2209 net6.n1659 net6.n1656 0.039
R2210 net6.n1529 net6.n1528 0.039
R2211 net6.n1589 net6.n1584 0.039
R2212 net6.n1490 net6.n1489 0.039
R2213 net6.n1446 net6.n1445 0.039
R2214 net6.n1297 net6.n1294 0.039
R2215 net6.n1167 net6.n1166 0.039
R2216 net6.n1227 net6.n1222 0.039
R2217 net6.n1128 net6.n1127 0.039
R2218 net6.n1084 net6.n1083 0.039
R2219 net6.n935 net6.n932 0.039
R2220 net6.n805 net6.n804 0.039
R2221 net6.n865 net6.n860 0.039
R2222 net6.n766 net6.n765 0.039
R2223 net6.n722 net6.n721 0.039
R2224 net6.n573 net6.n570 0.039
R2225 net6.n443 net6.n442 0.039
R2226 net6.n503 net6.n498 0.039
R2227 net6.n404 net6.n403 0.039
R2228 net6.n360 net6.n359 0.039
R2229 net6.n211 net6.n208 0.039
R2230 net6.n81 net6.n80 0.039
R2231 net6.n141 net6.n136 0.039
R2232 net6.n3624 net6.n3623 0.037
R2233 net6.n3263 net6.n3262 0.037
R2234 net6.n2902 net6.n2901 0.037
R2235 net6.n2541 net6.n2540 0.037
R2236 net6.n2180 net6.n2179 0.037
R2237 net6.n1818 net6.n1817 0.037
R2238 net6.n1456 net6.n1455 0.037
R2239 net6.n1094 net6.n1093 0.037
R2240 net6.n732 net6.n731 0.037
R2241 net6.n370 net6.n369 0.037
R2242 net6.n30 net6.n29 0.035
R2243 net6.n32 net6.n31 0.035
R2244 net6.n42 net6.n41 0.035
R2245 net6.n40 net6.n39 0.035
R2246 net6.n9 net6.n8 0.035
R2247 net6.n7 net6.n6 0.035
R2248 net6.n17 net6.n16 0.035
R2249 net6.n19 net6.n18 0.035
R2250 net6.n3325 net6.n3324 0.035
R2251 net6.n2964 net6.n2963 0.035
R2252 net6.n2603 net6.n2602 0.035
R2253 net6.n2242 net6.n2241 0.035
R2254 net6.n1881 net6.n1880 0.035
R2255 net6.n1519 net6.n1518 0.035
R2256 net6.n1157 net6.n1156 0.035
R2257 net6.n795 net6.n794 0.035
R2258 net6.n433 net6.n432 0.035
R2259 net6.n71 net6.n70 0.035
R2260 net6.n3603 net6.n3602 0.034
R2261 net6.n3435 net6.n3434 0.034
R2262 net6.n3548 net6.n3547 0.034
R2263 net6.n3541 net6.n3540 0.034
R2264 net6.n3497 net6.n3496 0.034
R2265 net6.n3486 net6.n3485 0.034
R2266 net6.n3408 net6.n3399 0.034
R2267 net6.n3393 net6.n3392 0.034
R2268 net6.n3242 net6.n3241 0.034
R2269 net6.n3074 net6.n3073 0.034
R2270 net6.n3187 net6.n3186 0.034
R2271 net6.n3180 net6.n3179 0.034
R2272 net6.n3136 net6.n3135 0.034
R2273 net6.n3125 net6.n3124 0.034
R2274 net6.n3047 net6.n3038 0.034
R2275 net6.n3032 net6.n3031 0.034
R2276 net6.n2881 net6.n2880 0.034
R2277 net6.n2713 net6.n2712 0.034
R2278 net6.n2826 net6.n2825 0.034
R2279 net6.n2819 net6.n2818 0.034
R2280 net6.n2775 net6.n2774 0.034
R2281 net6.n2764 net6.n2763 0.034
R2282 net6.n2686 net6.n2677 0.034
R2283 net6.n2671 net6.n2670 0.034
R2284 net6.n2520 net6.n2519 0.034
R2285 net6.n2352 net6.n2351 0.034
R2286 net6.n2465 net6.n2464 0.034
R2287 net6.n2458 net6.n2457 0.034
R2288 net6.n2414 net6.n2413 0.034
R2289 net6.n2403 net6.n2402 0.034
R2290 net6.n2325 net6.n2316 0.034
R2291 net6.n2310 net6.n2309 0.034
R2292 net6.n2159 net6.n2158 0.034
R2293 net6.n1991 net6.n1990 0.034
R2294 net6.n2104 net6.n2103 0.034
R2295 net6.n2097 net6.n2096 0.034
R2296 net6.n2053 net6.n2052 0.034
R2297 net6.n2042 net6.n2041 0.034
R2298 net6.n1964 net6.n1955 0.034
R2299 net6.n1949 net6.n1948 0.034
R2300 net6.n1797 net6.n1796 0.034
R2301 net6.n1629 net6.n1628 0.034
R2302 net6.n1742 net6.n1741 0.034
R2303 net6.n1735 net6.n1734 0.034
R2304 net6.n1691 net6.n1690 0.034
R2305 net6.n1680 net6.n1679 0.034
R2306 net6.n1602 net6.n1593 0.034
R2307 net6.n1587 net6.n1586 0.034
R2308 net6.n1435 net6.n1434 0.034
R2309 net6.n1267 net6.n1266 0.034
R2310 net6.n1380 net6.n1379 0.034
R2311 net6.n1373 net6.n1372 0.034
R2312 net6.n1329 net6.n1328 0.034
R2313 net6.n1318 net6.n1317 0.034
R2314 net6.n1240 net6.n1231 0.034
R2315 net6.n1225 net6.n1224 0.034
R2316 net6.n1073 net6.n1072 0.034
R2317 net6.n905 net6.n904 0.034
R2318 net6.n1018 net6.n1017 0.034
R2319 net6.n1011 net6.n1010 0.034
R2320 net6.n967 net6.n966 0.034
R2321 net6.n956 net6.n955 0.034
R2322 net6.n878 net6.n869 0.034
R2323 net6.n863 net6.n862 0.034
R2324 net6.n711 net6.n710 0.034
R2325 net6.n543 net6.n542 0.034
R2326 net6.n656 net6.n655 0.034
R2327 net6.n649 net6.n648 0.034
R2328 net6.n605 net6.n604 0.034
R2329 net6.n594 net6.n593 0.034
R2330 net6.n516 net6.n507 0.034
R2331 net6.n501 net6.n500 0.034
R2332 net6.n349 net6.n348 0.034
R2333 net6.n181 net6.n180 0.034
R2334 net6.n294 net6.n293 0.034
R2335 net6.n287 net6.n286 0.034
R2336 net6.n243 net6.n242 0.034
R2337 net6.n232 net6.n231 0.034
R2338 net6.n154 net6.n145 0.034
R2339 net6.n139 net6.n138 0.034
R2340 net6.n3666 net6.n3665 0.032
R2341 net6.n3473 net6.n3470 0.032
R2342 net6.n3366 net6.n3365 0.032
R2343 net6.n3504 net6.n3503 0.032
R2344 net6.n3305 net6.n3304 0.032
R2345 net6.n3112 net6.n3109 0.032
R2346 net6.n3005 net6.n3004 0.032
R2347 net6.n3143 net6.n3142 0.032
R2348 net6.n2944 net6.n2943 0.032
R2349 net6.n2751 net6.n2748 0.032
R2350 net6.n2644 net6.n2643 0.032
R2351 net6.n2782 net6.n2781 0.032
R2352 net6.n2583 net6.n2582 0.032
R2353 net6.n2390 net6.n2387 0.032
R2354 net6.n2283 net6.n2282 0.032
R2355 net6.n2421 net6.n2420 0.032
R2356 net6.n2222 net6.n2221 0.032
R2357 net6.n2029 net6.n2026 0.032
R2358 net6.n1922 net6.n1921 0.032
R2359 net6.n2060 net6.n2059 0.032
R2360 net6.n1860 net6.n1859 0.032
R2361 net6.n1667 net6.n1664 0.032
R2362 net6.n1560 net6.n1559 0.032
R2363 net6.n1698 net6.n1697 0.032
R2364 net6.n1498 net6.n1497 0.032
R2365 net6.n1305 net6.n1302 0.032
R2366 net6.n1198 net6.n1197 0.032
R2367 net6.n1336 net6.n1335 0.032
R2368 net6.n1136 net6.n1135 0.032
R2369 net6.n943 net6.n940 0.032
R2370 net6.n836 net6.n835 0.032
R2371 net6.n974 net6.n973 0.032
R2372 net6.n774 net6.n773 0.032
R2373 net6.n581 net6.n578 0.032
R2374 net6.n474 net6.n473 0.032
R2375 net6.n612 net6.n611 0.032
R2376 net6.n412 net6.n411 0.032
R2377 net6.n219 net6.n216 0.032
R2378 net6.n112 net6.n111 0.032
R2379 net6.n250 net6.n249 0.032
R2380 net6.n3569 net6.n3568 0.031
R2381 net6.n3550 net6.n3546 0.031
R2382 net6.n3527 net6.n3526 0.031
R2383 net6.n3508 net6.n3502 0.031
R2384 net6.n3483 net6.n3482 0.031
R2385 net6.n3419 net6.n3413 0.031
R2386 net6.n3388 net6.n3387 0.031
R2387 net6.n3373 net6.n3372 0.031
R2388 net6.n3208 net6.n3207 0.031
R2389 net6.n3189 net6.n3185 0.031
R2390 net6.n3166 net6.n3165 0.031
R2391 net6.n3147 net6.n3141 0.031
R2392 net6.n3122 net6.n3121 0.031
R2393 net6.n3058 net6.n3052 0.031
R2394 net6.n3027 net6.n3026 0.031
R2395 net6.n3012 net6.n3011 0.031
R2396 net6.n2847 net6.n2846 0.031
R2397 net6.n2828 net6.n2824 0.031
R2398 net6.n2805 net6.n2804 0.031
R2399 net6.n2786 net6.n2780 0.031
R2400 net6.n2761 net6.n2760 0.031
R2401 net6.n2697 net6.n2691 0.031
R2402 net6.n2666 net6.n2665 0.031
R2403 net6.n2651 net6.n2650 0.031
R2404 net6.n2486 net6.n2485 0.031
R2405 net6.n2467 net6.n2463 0.031
R2406 net6.n2444 net6.n2443 0.031
R2407 net6.n2425 net6.n2419 0.031
R2408 net6.n2400 net6.n2399 0.031
R2409 net6.n2336 net6.n2330 0.031
R2410 net6.n2305 net6.n2304 0.031
R2411 net6.n2290 net6.n2289 0.031
R2412 net6.n2125 net6.n2124 0.031
R2413 net6.n2106 net6.n2102 0.031
R2414 net6.n2083 net6.n2082 0.031
R2415 net6.n2064 net6.n2058 0.031
R2416 net6.n2039 net6.n2038 0.031
R2417 net6.n1975 net6.n1969 0.031
R2418 net6.n1944 net6.n1943 0.031
R2419 net6.n1929 net6.n1928 0.031
R2420 net6.n1763 net6.n1762 0.031
R2421 net6.n1744 net6.n1740 0.031
R2422 net6.n1721 net6.n1720 0.031
R2423 net6.n1702 net6.n1696 0.031
R2424 net6.n1677 net6.n1676 0.031
R2425 net6.n1613 net6.n1607 0.031
R2426 net6.n1582 net6.n1581 0.031
R2427 net6.n1567 net6.n1566 0.031
R2428 net6.n1401 net6.n1400 0.031
R2429 net6.n1382 net6.n1378 0.031
R2430 net6.n1359 net6.n1358 0.031
R2431 net6.n1340 net6.n1334 0.031
R2432 net6.n1315 net6.n1314 0.031
R2433 net6.n1251 net6.n1245 0.031
R2434 net6.n1220 net6.n1219 0.031
R2435 net6.n1205 net6.n1204 0.031
R2436 net6.n1039 net6.n1038 0.031
R2437 net6.n1020 net6.n1016 0.031
R2438 net6.n997 net6.n996 0.031
R2439 net6.n978 net6.n972 0.031
R2440 net6.n953 net6.n952 0.031
R2441 net6.n889 net6.n883 0.031
R2442 net6.n858 net6.n857 0.031
R2443 net6.n843 net6.n842 0.031
R2444 net6.n677 net6.n676 0.031
R2445 net6.n658 net6.n654 0.031
R2446 net6.n635 net6.n634 0.031
R2447 net6.n616 net6.n610 0.031
R2448 net6.n591 net6.n590 0.031
R2449 net6.n527 net6.n521 0.031
R2450 net6.n496 net6.n495 0.031
R2451 net6.n481 net6.n480 0.031
R2452 net6.n315 net6.n314 0.031
R2453 net6.n296 net6.n292 0.031
R2454 net6.n273 net6.n272 0.031
R2455 net6.n254 net6.n248 0.031
R2456 net6.n229 net6.n228 0.031
R2457 net6.n165 net6.n159 0.031
R2458 net6.n134 net6.n133 0.031
R2459 net6.n119 net6.n118 0.031
R2460 net6.n3645 net6.n3641 0.03
R2461 net6.n3589 net6.n3586 0.03
R2462 net6.n3444 net6.n3441 0.03
R2463 net6.n3339 net6.n3338 0.03
R2464 net6.n3356 net6.n3355 0.03
R2465 net6.n3488 net6.n3487 0.03
R2466 net6.n3284 net6.n3280 0.03
R2467 net6.n3228 net6.n3225 0.03
R2468 net6.n3083 net6.n3080 0.03
R2469 net6.n2978 net6.n2977 0.03
R2470 net6.n2995 net6.n2994 0.03
R2471 net6.n3127 net6.n3126 0.03
R2472 net6.n2923 net6.n2919 0.03
R2473 net6.n2867 net6.n2864 0.03
R2474 net6.n2722 net6.n2719 0.03
R2475 net6.n2617 net6.n2616 0.03
R2476 net6.n2634 net6.n2633 0.03
R2477 net6.n2766 net6.n2765 0.03
R2478 net6.n2562 net6.n2558 0.03
R2479 net6.n2506 net6.n2503 0.03
R2480 net6.n2361 net6.n2358 0.03
R2481 net6.n2256 net6.n2255 0.03
R2482 net6.n2273 net6.n2272 0.03
R2483 net6.n2405 net6.n2404 0.03
R2484 net6.n2201 net6.n2197 0.03
R2485 net6.n2145 net6.n2142 0.03
R2486 net6.n2000 net6.n1997 0.03
R2487 net6.n1895 net6.n1894 0.03
R2488 net6.n1912 net6.n1911 0.03
R2489 net6.n2044 net6.n2043 0.03
R2490 net6.n1839 net6.n1835 0.03
R2491 net6.n1783 net6.n1780 0.03
R2492 net6.n1638 net6.n1635 0.03
R2493 net6.n1533 net6.n1532 0.03
R2494 net6.n1550 net6.n1549 0.03
R2495 net6.n1682 net6.n1681 0.03
R2496 net6.n1477 net6.n1473 0.03
R2497 net6.n1421 net6.n1418 0.03
R2498 net6.n1276 net6.n1273 0.03
R2499 net6.n1171 net6.n1170 0.03
R2500 net6.n1188 net6.n1187 0.03
R2501 net6.n1320 net6.n1319 0.03
R2502 net6.n1115 net6.n1111 0.03
R2503 net6.n1059 net6.n1056 0.03
R2504 net6.n914 net6.n911 0.03
R2505 net6.n809 net6.n808 0.03
R2506 net6.n826 net6.n825 0.03
R2507 net6.n958 net6.n957 0.03
R2508 net6.n753 net6.n749 0.03
R2509 net6.n697 net6.n694 0.03
R2510 net6.n552 net6.n549 0.03
R2511 net6.n447 net6.n446 0.03
R2512 net6.n464 net6.n463 0.03
R2513 net6.n596 net6.n595 0.03
R2514 net6.n391 net6.n387 0.03
R2515 net6.n335 net6.n332 0.03
R2516 net6.n190 net6.n187 0.03
R2517 net6.n85 net6.n84 0.03
R2518 net6.n102 net6.n101 0.03
R2519 net6.n234 net6.n233 0.03
R2520 net6.n48 net6.n37 0.029
R2521 net6.n48 net6.n47 0.029
R2522 net6.n50 net6.n49 0.029
R2523 net6.n31 net6.n30 0.028
R2524 net6.n41 net6.n40 0.028
R2525 net6.n8 net6.n7 0.028
R2526 net6.n54 net6.n53 0.028
R2527 net6.n24 net6.n23 0.028
R2528 net6.n18 net6.n17 0.028
R2529 net6.n3656 net6.n3655 0.028
R2530 net6.n3599 net6.n3597 0.028
R2531 net6.n3478 net6.n3475 0.028
R2532 net6.n3468 net6.n3467 0.028
R2533 net6.n3559 net6.n3558 0.028
R2534 net6.n3534 net6.n3533 0.028
R2535 net6.n3532 net6.n3531 0.028
R2536 net6.n3493 net6.n3492 0.028
R2537 net6.n3295 net6.n3294 0.028
R2538 net6.n3238 net6.n3236 0.028
R2539 net6.n3117 net6.n3114 0.028
R2540 net6.n3107 net6.n3106 0.028
R2541 net6.n3198 net6.n3197 0.028
R2542 net6.n3173 net6.n3172 0.028
R2543 net6.n3171 net6.n3170 0.028
R2544 net6.n3132 net6.n3131 0.028
R2545 net6.n2934 net6.n2933 0.028
R2546 net6.n2877 net6.n2875 0.028
R2547 net6.n2756 net6.n2753 0.028
R2548 net6.n2746 net6.n2745 0.028
R2549 net6.n2837 net6.n2836 0.028
R2550 net6.n2812 net6.n2811 0.028
R2551 net6.n2810 net6.n2809 0.028
R2552 net6.n2771 net6.n2770 0.028
R2553 net6.n2573 net6.n2572 0.028
R2554 net6.n2516 net6.n2514 0.028
R2555 net6.n2395 net6.n2392 0.028
R2556 net6.n2385 net6.n2384 0.028
R2557 net6.n2476 net6.n2475 0.028
R2558 net6.n2451 net6.n2450 0.028
R2559 net6.n2449 net6.n2448 0.028
R2560 net6.n2410 net6.n2409 0.028
R2561 net6.n2212 net6.n2211 0.028
R2562 net6.n2155 net6.n2153 0.028
R2563 net6.n2034 net6.n2031 0.028
R2564 net6.n2024 net6.n2023 0.028
R2565 net6.n2115 net6.n2114 0.028
R2566 net6.n2090 net6.n2089 0.028
R2567 net6.n2088 net6.n2087 0.028
R2568 net6.n2049 net6.n2048 0.028
R2569 net6.n1850 net6.n1849 0.028
R2570 net6.n1793 net6.n1791 0.028
R2571 net6.n1672 net6.n1669 0.028
R2572 net6.n1662 net6.n1661 0.028
R2573 net6.n1753 net6.n1752 0.028
R2574 net6.n1728 net6.n1727 0.028
R2575 net6.n1726 net6.n1725 0.028
R2576 net6.n1687 net6.n1686 0.028
R2577 net6.n1488 net6.n1487 0.028
R2578 net6.n1431 net6.n1429 0.028
R2579 net6.n1310 net6.n1307 0.028
R2580 net6.n1300 net6.n1299 0.028
R2581 net6.n1391 net6.n1390 0.028
R2582 net6.n1366 net6.n1365 0.028
R2583 net6.n1364 net6.n1363 0.028
R2584 net6.n1325 net6.n1324 0.028
R2585 net6.n1126 net6.n1125 0.028
R2586 net6.n1069 net6.n1067 0.028
R2587 net6.n948 net6.n945 0.028
R2588 net6.n938 net6.n937 0.028
R2589 net6.n1029 net6.n1028 0.028
R2590 net6.n1004 net6.n1003 0.028
R2591 net6.n1002 net6.n1001 0.028
R2592 net6.n963 net6.n962 0.028
R2593 net6.n764 net6.n763 0.028
R2594 net6.n707 net6.n705 0.028
R2595 net6.n586 net6.n583 0.028
R2596 net6.n576 net6.n575 0.028
R2597 net6.n667 net6.n666 0.028
R2598 net6.n642 net6.n641 0.028
R2599 net6.n640 net6.n639 0.028
R2600 net6.n601 net6.n600 0.028
R2601 net6.n402 net6.n401 0.028
R2602 net6.n345 net6.n343 0.028
R2603 net6.n224 net6.n221 0.028
R2604 net6.n214 net6.n213 0.028
R2605 net6.n305 net6.n304 0.028
R2606 net6.n280 net6.n279 0.028
R2607 net6.n278 net6.n277 0.028
R2608 net6.n239 net6.n238 0.028
R2609 net6.n3371 net6.n3328 0.027
R2610 net6.n3010 net6.n2967 0.027
R2611 net6.n2649 net6.n2606 0.027
R2612 net6.n2288 net6.n2245 0.027
R2613 net6.n1927 net6.n1884 0.027
R2614 net6.n1565 net6.n1522 0.027
R2615 net6.n1203 net6.n1160 0.027
R2616 net6.n841 net6.n798 0.027
R2617 net6.n479 net6.n436 0.027
R2618 net6.n117 net6.n74 0.027
R2619 net6.n3561 net6.n3557 0.027
R2620 net6.n3519 net6.n3515 0.027
R2621 net6.n3430 net6.n3426 0.027
R2622 net6.n3380 net6.n3376 0.027
R2623 net6.n3200 net6.n3196 0.027
R2624 net6.n3158 net6.n3154 0.027
R2625 net6.n3069 net6.n3065 0.027
R2626 net6.n3019 net6.n3015 0.027
R2627 net6.n2839 net6.n2835 0.027
R2628 net6.n2797 net6.n2793 0.027
R2629 net6.n2708 net6.n2704 0.027
R2630 net6.n2658 net6.n2654 0.027
R2631 net6.n2478 net6.n2474 0.027
R2632 net6.n2436 net6.n2432 0.027
R2633 net6.n2347 net6.n2343 0.027
R2634 net6.n2297 net6.n2293 0.027
R2635 net6.n2117 net6.n2113 0.027
R2636 net6.n2075 net6.n2071 0.027
R2637 net6.n1986 net6.n1982 0.027
R2638 net6.n1936 net6.n1932 0.027
R2639 net6.n1755 net6.n1751 0.027
R2640 net6.n1713 net6.n1709 0.027
R2641 net6.n1624 net6.n1620 0.027
R2642 net6.n1574 net6.n1570 0.027
R2643 net6.n1393 net6.n1389 0.027
R2644 net6.n1351 net6.n1347 0.027
R2645 net6.n1262 net6.n1258 0.027
R2646 net6.n1212 net6.n1208 0.027
R2647 net6.n1031 net6.n1027 0.027
R2648 net6.n989 net6.n985 0.027
R2649 net6.n900 net6.n896 0.027
R2650 net6.n850 net6.n846 0.027
R2651 net6.n669 net6.n665 0.027
R2652 net6.n627 net6.n623 0.027
R2653 net6.n538 net6.n534 0.027
R2654 net6.n488 net6.n484 0.027
R2655 net6.n307 net6.n303 0.027
R2656 net6.n265 net6.n261 0.027
R2657 net6.n176 net6.n172 0.027
R2658 net6.n126 net6.n122 0.027
R2659 net6.n3606 net6.n3605 0.026
R2660 net6.n3674 net6.n3673 0.026
R2661 net6.n3517 net6.n3516 0.026
R2662 net6.n3415 net6.n3414 0.026
R2663 net6.n3398 net6.n3397 0.026
R2664 net6.n3245 net6.n3244 0.026
R2665 net6.n3313 net6.n3312 0.026
R2666 net6.n3156 net6.n3155 0.026
R2667 net6.n3054 net6.n3053 0.026
R2668 net6.n3037 net6.n3036 0.026
R2669 net6.n2884 net6.n2883 0.026
R2670 net6.n2952 net6.n2951 0.026
R2671 net6.n2795 net6.n2794 0.026
R2672 net6.n2693 net6.n2692 0.026
R2673 net6.n2676 net6.n2675 0.026
R2674 net6.n2523 net6.n2522 0.026
R2675 net6.n2591 net6.n2590 0.026
R2676 net6.n2434 net6.n2433 0.026
R2677 net6.n2332 net6.n2331 0.026
R2678 net6.n2315 net6.n2314 0.026
R2679 net6.n2162 net6.n2161 0.026
R2680 net6.n2230 net6.n2229 0.026
R2681 net6.n2073 net6.n2072 0.026
R2682 net6.n1971 net6.n1970 0.026
R2683 net6.n1954 net6.n1953 0.026
R2684 net6.n1800 net6.n1799 0.026
R2685 net6.n1868 net6.n1867 0.026
R2686 net6.n1711 net6.n1710 0.026
R2687 net6.n1609 net6.n1608 0.026
R2688 net6.n1592 net6.n1591 0.026
R2689 net6.n1438 net6.n1437 0.026
R2690 net6.n1506 net6.n1505 0.026
R2691 net6.n1349 net6.n1348 0.026
R2692 net6.n1247 net6.n1246 0.026
R2693 net6.n1230 net6.n1229 0.026
R2694 net6.n1076 net6.n1075 0.026
R2695 net6.n1144 net6.n1143 0.026
R2696 net6.n987 net6.n986 0.026
R2697 net6.n885 net6.n884 0.026
R2698 net6.n868 net6.n867 0.026
R2699 net6.n714 net6.n713 0.026
R2700 net6.n782 net6.n781 0.026
R2701 net6.n625 net6.n624 0.026
R2702 net6.n523 net6.n522 0.026
R2703 net6.n506 net6.n505 0.026
R2704 net6.n352 net6.n351 0.026
R2705 net6.n420 net6.n419 0.026
R2706 net6.n263 net6.n262 0.026
R2707 net6.n161 net6.n160 0.026
R2708 net6.n144 net6.n143 0.026
R2709 net6.n3466 net6.n3465 0.024
R2710 net6.n3567 net6.n3566 0.024
R2711 net6.n3556 net6.n3555 0.024
R2712 net6.n3525 net6.n3524 0.024
R2713 net6.n3514 net6.n3513 0.024
R2714 net6.n3481 net6.n3480 0.024
R2715 net6.n3425 net6.n3424 0.024
R2716 net6.n3320 net6.n3319 0.024
R2717 net6.n3327 net6.n3326 0.024
R2718 net6.n3105 net6.n3104 0.024
R2719 net6.n3206 net6.n3205 0.024
R2720 net6.n3195 net6.n3194 0.024
R2721 net6.n3164 net6.n3163 0.024
R2722 net6.n3153 net6.n3152 0.024
R2723 net6.n3120 net6.n3119 0.024
R2724 net6.n3064 net6.n3063 0.024
R2725 net6.n2959 net6.n2958 0.024
R2726 net6.n2966 net6.n2965 0.024
R2727 net6.n2744 net6.n2743 0.024
R2728 net6.n2845 net6.n2844 0.024
R2729 net6.n2834 net6.n2833 0.024
R2730 net6.n2803 net6.n2802 0.024
R2731 net6.n2792 net6.n2791 0.024
R2732 net6.n2759 net6.n2758 0.024
R2733 net6.n2703 net6.n2702 0.024
R2734 net6.n2598 net6.n2597 0.024
R2735 net6.n2605 net6.n2604 0.024
R2736 net6.n2383 net6.n2382 0.024
R2737 net6.n2484 net6.n2483 0.024
R2738 net6.n2473 net6.n2472 0.024
R2739 net6.n2442 net6.n2441 0.024
R2740 net6.n2431 net6.n2430 0.024
R2741 net6.n2398 net6.n2397 0.024
R2742 net6.n2342 net6.n2341 0.024
R2743 net6.n2237 net6.n2236 0.024
R2744 net6.n2244 net6.n2243 0.024
R2745 net6.n2022 net6.n2021 0.024
R2746 net6.n2123 net6.n2122 0.024
R2747 net6.n2112 net6.n2111 0.024
R2748 net6.n2081 net6.n2080 0.024
R2749 net6.n2070 net6.n2069 0.024
R2750 net6.n2037 net6.n2036 0.024
R2751 net6.n1981 net6.n1980 0.024
R2752 net6.n1876 net6.n1875 0.024
R2753 net6.n1883 net6.n1882 0.024
R2754 net6.n1660 net6.n1659 0.024
R2755 net6.n1761 net6.n1760 0.024
R2756 net6.n1750 net6.n1749 0.024
R2757 net6.n1719 net6.n1718 0.024
R2758 net6.n1708 net6.n1707 0.024
R2759 net6.n1675 net6.n1674 0.024
R2760 net6.n1619 net6.n1618 0.024
R2761 net6.n1514 net6.n1513 0.024
R2762 net6.n1521 net6.n1520 0.024
R2763 net6.n1298 net6.n1297 0.024
R2764 net6.n1399 net6.n1398 0.024
R2765 net6.n1388 net6.n1387 0.024
R2766 net6.n1357 net6.n1356 0.024
R2767 net6.n1346 net6.n1345 0.024
R2768 net6.n1313 net6.n1312 0.024
R2769 net6.n1257 net6.n1256 0.024
R2770 net6.n1152 net6.n1151 0.024
R2771 net6.n1159 net6.n1158 0.024
R2772 net6.n936 net6.n935 0.024
R2773 net6.n1037 net6.n1036 0.024
R2774 net6.n1026 net6.n1025 0.024
R2775 net6.n995 net6.n994 0.024
R2776 net6.n984 net6.n983 0.024
R2777 net6.n951 net6.n950 0.024
R2778 net6.n895 net6.n894 0.024
R2779 net6.n790 net6.n789 0.024
R2780 net6.n797 net6.n796 0.024
R2781 net6.n574 net6.n573 0.024
R2782 net6.n675 net6.n674 0.024
R2783 net6.n664 net6.n663 0.024
R2784 net6.n633 net6.n632 0.024
R2785 net6.n622 net6.n621 0.024
R2786 net6.n589 net6.n588 0.024
R2787 net6.n533 net6.n532 0.024
R2788 net6.n428 net6.n427 0.024
R2789 net6.n435 net6.n434 0.024
R2790 net6.n212 net6.n211 0.024
R2791 net6.n313 net6.n312 0.024
R2792 net6.n302 net6.n301 0.024
R2793 net6.n271 net6.n270 0.024
R2794 net6.n260 net6.n259 0.024
R2795 net6.n227 net6.n226 0.024
R2796 net6.n171 net6.n170 0.024
R2797 net6.n66 net6.n65 0.024
R2798 net6.n73 net6.n72 0.024
R2799 net6.n35 net6.n34 0.023
R2800 net6.n45 net6.n44 0.023
R2801 net6.n55 net6.n54 0.023
R2802 net6.n25 net6.n24 0.023
R2803 net6.n58 net6.n57 0.022
R2804 net6.n51 net6.n27 0.022
R2805 net6.n3610 net6.n3608 0.022
R2806 net6.n3605 net6.n3604 0.022
R2807 net6.n3676 net6.n3675 0.022
R2808 net6.n3385 net6.n3384 0.022
R2809 net6.n3323 net6.n3322 0.022
R2810 net6.n3328 net6.n3327 0.022
R2811 net6.n3249 net6.n3247 0.022
R2812 net6.n3244 net6.n3243 0.022
R2813 net6.n3315 net6.n3314 0.022
R2814 net6.n3024 net6.n3023 0.022
R2815 net6.n2962 net6.n2961 0.022
R2816 net6.n2967 net6.n2966 0.022
R2817 net6.n2888 net6.n2886 0.022
R2818 net6.n2883 net6.n2882 0.022
R2819 net6.n2954 net6.n2953 0.022
R2820 net6.n2663 net6.n2662 0.022
R2821 net6.n2601 net6.n2600 0.022
R2822 net6.n2606 net6.n2605 0.022
R2823 net6.n2527 net6.n2525 0.022
R2824 net6.n2522 net6.n2521 0.022
R2825 net6.n2593 net6.n2592 0.022
R2826 net6.n2302 net6.n2301 0.022
R2827 net6.n2240 net6.n2239 0.022
R2828 net6.n2245 net6.n2244 0.022
R2829 net6.n2166 net6.n2164 0.022
R2830 net6.n2161 net6.n2160 0.022
R2831 net6.n2232 net6.n2231 0.022
R2832 net6.n1941 net6.n1940 0.022
R2833 net6.n1879 net6.n1878 0.022
R2834 net6.n1884 net6.n1883 0.022
R2835 net6.n1804 net6.n1802 0.022
R2836 net6.n1799 net6.n1798 0.022
R2837 net6.n1870 net6.n1869 0.022
R2838 net6.n1579 net6.n1578 0.022
R2839 net6.n1517 net6.n1516 0.022
R2840 net6.n1522 net6.n1521 0.022
R2841 net6.n1442 net6.n1440 0.022
R2842 net6.n1437 net6.n1436 0.022
R2843 net6.n1508 net6.n1507 0.022
R2844 net6.n1217 net6.n1216 0.022
R2845 net6.n1155 net6.n1154 0.022
R2846 net6.n1160 net6.n1159 0.022
R2847 net6.n1080 net6.n1078 0.022
R2848 net6.n1075 net6.n1074 0.022
R2849 net6.n1146 net6.n1145 0.022
R2850 net6.n855 net6.n854 0.022
R2851 net6.n793 net6.n792 0.022
R2852 net6.n798 net6.n797 0.022
R2853 net6.n718 net6.n716 0.022
R2854 net6.n713 net6.n712 0.022
R2855 net6.n784 net6.n783 0.022
R2856 net6.n493 net6.n492 0.022
R2857 net6.n431 net6.n430 0.022
R2858 net6.n436 net6.n435 0.022
R2859 net6.n356 net6.n354 0.022
R2860 net6.n351 net6.n350 0.022
R2861 net6.n422 net6.n421 0.022
R2862 net6.n131 net6.n130 0.022
R2863 net6.n69 net6.n68 0.022
R2864 net6.n74 net6.n73 0.022
R2865 net6.n57 net6.n56 0.02
R2866 net6.n27 net6.n26 0.02
R2867 net6.n3621 net6.n3620 0.02
R2868 net6.n3469 net6.n3468 0.02
R2869 net6.n3458 net6.n3457 0.02
R2870 net6.n3675 net6.n3674 0.02
R2871 net6.n3428 net6.n3427 0.02
R2872 net6.n3260 net6.n3259 0.02
R2873 net6.n3108 net6.n3107 0.02
R2874 net6.n3097 net6.n3096 0.02
R2875 net6.n3314 net6.n3313 0.02
R2876 net6.n3067 net6.n3066 0.02
R2877 net6.n2899 net6.n2898 0.02
R2878 net6.n2747 net6.n2746 0.02
R2879 net6.n2736 net6.n2735 0.02
R2880 net6.n2953 net6.n2952 0.02
R2881 net6.n2706 net6.n2705 0.02
R2882 net6.n2538 net6.n2537 0.02
R2883 net6.n2386 net6.n2385 0.02
R2884 net6.n2375 net6.n2374 0.02
R2885 net6.n2592 net6.n2591 0.02
R2886 net6.n2345 net6.n2344 0.02
R2887 net6.n2177 net6.n2176 0.02
R2888 net6.n2025 net6.n2024 0.02
R2889 net6.n2014 net6.n2013 0.02
R2890 net6.n2231 net6.n2230 0.02
R2891 net6.n1984 net6.n1983 0.02
R2892 net6.n1815 net6.n1814 0.02
R2893 net6.n1663 net6.n1662 0.02
R2894 net6.n1652 net6.n1651 0.02
R2895 net6.n1869 net6.n1868 0.02
R2896 net6.n1622 net6.n1621 0.02
R2897 net6.n1453 net6.n1452 0.02
R2898 net6.n1301 net6.n1300 0.02
R2899 net6.n1290 net6.n1289 0.02
R2900 net6.n1507 net6.n1506 0.02
R2901 net6.n1260 net6.n1259 0.02
R2902 net6.n1091 net6.n1090 0.02
R2903 net6.n939 net6.n938 0.02
R2904 net6.n928 net6.n927 0.02
R2905 net6.n1145 net6.n1144 0.02
R2906 net6.n898 net6.n897 0.02
R2907 net6.n729 net6.n728 0.02
R2908 net6.n577 net6.n576 0.02
R2909 net6.n566 net6.n565 0.02
R2910 net6.n783 net6.n782 0.02
R2911 net6.n536 net6.n535 0.02
R2912 net6.n367 net6.n366 0.02
R2913 net6.n215 net6.n214 0.02
R2914 net6.n204 net6.n203 0.02
R2915 net6.n421 net6.n420 0.02
R2916 net6.n174 net6.n173 0.02
R2917 net6.n3378 net6.n3377 0.018
R2918 net6.n3017 net6.n3016 0.018
R2919 net6.n2656 net6.n2655 0.018
R2920 net6.n2295 net6.n2294 0.018
R2921 net6.n1934 net6.n1933 0.018
R2922 net6.n1572 net6.n1571 0.018
R2923 net6.n1210 net6.n1209 0.018
R2924 net6.n848 net6.n847 0.018
R2925 net6.n486 net6.n485 0.018
R2926 net6.n124 net6.n123 0.018
R2927 net6 net6.n3682 0.018
R2928 net6.n36 net6.n35 0.017
R2929 net6.n46 net6.n45 0.017
R2930 net6.n56 net6.n55 0.017
R2931 net6.n26 net6.n25 0.017
R2932 net6.n3633 net6.n3632 0.017
R2933 net6.n3353 net6.n3349 0.017
R2934 net6.n3379 net6.n3378 0.017
R2935 net6.n3272 net6.n3271 0.017
R2936 net6.n2992 net6.n2988 0.017
R2937 net6.n3018 net6.n3017 0.017
R2938 net6.n2911 net6.n2910 0.017
R2939 net6.n2631 net6.n2627 0.017
R2940 net6.n2657 net6.n2656 0.017
R2941 net6.n2550 net6.n2549 0.017
R2942 net6.n2270 net6.n2266 0.017
R2943 net6.n2296 net6.n2295 0.017
R2944 net6.n2189 net6.n2188 0.017
R2945 net6.n1909 net6.n1905 0.017
R2946 net6.n1935 net6.n1934 0.017
R2947 net6.n1827 net6.n1826 0.017
R2948 net6.n1547 net6.n1543 0.017
R2949 net6.n1573 net6.n1572 0.017
R2950 net6.n1465 net6.n1464 0.017
R2951 net6.n1185 net6.n1181 0.017
R2952 net6.n1211 net6.n1210 0.017
R2953 net6.n1103 net6.n1102 0.017
R2954 net6.n823 net6.n819 0.017
R2955 net6.n849 net6.n848 0.017
R2956 net6.n741 net6.n740 0.017
R2957 net6.n461 net6.n457 0.017
R2958 net6.n487 net6.n486 0.017
R2959 net6.n379 net6.n378 0.017
R2960 net6.n99 net6.n95 0.017
R2961 net6.n125 net6.n124 0.017
R2962 net6.n3570 net6.n3569 0.016
R2963 net6.n3546 net6.n3545 0.016
R2964 net6.n3528 net6.n3527 0.016
R2965 net6.n3502 net6.n3501 0.016
R2966 net6.n3484 net6.n3483 0.016
R2967 net6.n3413 net6.n3412 0.016
R2968 net6.n3389 net6.n3388 0.016
R2969 net6.n3209 net6.n3208 0.016
R2970 net6.n3185 net6.n3184 0.016
R2971 net6.n3167 net6.n3166 0.016
R2972 net6.n3141 net6.n3140 0.016
R2973 net6.n3123 net6.n3122 0.016
R2974 net6.n3052 net6.n3051 0.016
R2975 net6.n3028 net6.n3027 0.016
R2976 net6.n2848 net6.n2847 0.016
R2977 net6.n2824 net6.n2823 0.016
R2978 net6.n2806 net6.n2805 0.016
R2979 net6.n2780 net6.n2779 0.016
R2980 net6.n2762 net6.n2761 0.016
R2981 net6.n2691 net6.n2690 0.016
R2982 net6.n2667 net6.n2666 0.016
R2983 net6.n2487 net6.n2486 0.016
R2984 net6.n2463 net6.n2462 0.016
R2985 net6.n2445 net6.n2444 0.016
R2986 net6.n2419 net6.n2418 0.016
R2987 net6.n2401 net6.n2400 0.016
R2988 net6.n2330 net6.n2329 0.016
R2989 net6.n2306 net6.n2305 0.016
R2990 net6.n2126 net6.n2125 0.016
R2991 net6.n2102 net6.n2101 0.016
R2992 net6.n2084 net6.n2083 0.016
R2993 net6.n2058 net6.n2057 0.016
R2994 net6.n2040 net6.n2039 0.016
R2995 net6.n1969 net6.n1968 0.016
R2996 net6.n1945 net6.n1944 0.016
R2997 net6.n1764 net6.n1763 0.016
R2998 net6.n1740 net6.n1739 0.016
R2999 net6.n1722 net6.n1721 0.016
R3000 net6.n1696 net6.n1695 0.016
R3001 net6.n1678 net6.n1677 0.016
R3002 net6.n1607 net6.n1606 0.016
R3003 net6.n1583 net6.n1582 0.016
R3004 net6.n1402 net6.n1401 0.016
R3005 net6.n1378 net6.n1377 0.016
R3006 net6.n1360 net6.n1359 0.016
R3007 net6.n1334 net6.n1333 0.016
R3008 net6.n1316 net6.n1315 0.016
R3009 net6.n1245 net6.n1244 0.016
R3010 net6.n1221 net6.n1220 0.016
R3011 net6.n1040 net6.n1039 0.016
R3012 net6.n1016 net6.n1015 0.016
R3013 net6.n998 net6.n997 0.016
R3014 net6.n972 net6.n971 0.016
R3015 net6.n954 net6.n953 0.016
R3016 net6.n883 net6.n882 0.016
R3017 net6.n859 net6.n858 0.016
R3018 net6.n678 net6.n677 0.016
R3019 net6.n654 net6.n653 0.016
R3020 net6.n636 net6.n635 0.016
R3021 net6.n610 net6.n609 0.016
R3022 net6.n592 net6.n591 0.016
R3023 net6.n521 net6.n520 0.016
R3024 net6.n497 net6.n496 0.016
R3025 net6.n316 net6.n315 0.016
R3026 net6.n292 net6.n291 0.016
R3027 net6.n274 net6.n273 0.016
R3028 net6.n248 net6.n247 0.016
R3029 net6.n230 net6.n229 0.016
R3030 net6.n159 net6.n158 0.016
R3031 net6.n135 net6.n134 0.016
R3032 net6.n3661 net6.n3660 0.015
R3033 net6.n3655 net6.n3654 0.015
R3034 net6.n3653 net6.n3652 0.015
R3035 net6.n3470 net6.n3469 0.015
R3036 net6.n3355 net6.n3354 0.015
R3037 net6.n3361 net6.n3360 0.015
R3038 net6.n3566 net6.n3565 0.015
R3039 net6.n3556 net6.n3553 0.015
R3040 net6.n3555 net6.n3554 0.015
R3041 net6.n3533 net6.n3532 0.015
R3042 net6.n3524 net6.n3523 0.015
R3043 net6.n3513 net6.n3512 0.015
R3044 net6.n3480 net6.n3479 0.015
R3045 net6.n3429 net6.n3428 0.015
R3046 net6.n3424 net6.n3423 0.015
R3047 net6.n3384 net6.n3383 0.015
R3048 net6.n3321 net6.n3320 0.015
R3049 net6.n3300 net6.n3299 0.015
R3050 net6.n3294 net6.n3293 0.015
R3051 net6.n3292 net6.n3291 0.015
R3052 net6.n3109 net6.n3108 0.015
R3053 net6.n2994 net6.n2993 0.015
R3054 net6.n3000 net6.n2999 0.015
R3055 net6.n3205 net6.n3204 0.015
R3056 net6.n3195 net6.n3192 0.015
R3057 net6.n3194 net6.n3193 0.015
R3058 net6.n3172 net6.n3171 0.015
R3059 net6.n3163 net6.n3162 0.015
R3060 net6.n3152 net6.n3151 0.015
R3061 net6.n3119 net6.n3118 0.015
R3062 net6.n3068 net6.n3067 0.015
R3063 net6.n3063 net6.n3062 0.015
R3064 net6.n3023 net6.n3022 0.015
R3065 net6.n2960 net6.n2959 0.015
R3066 net6.n2939 net6.n2938 0.015
R3067 net6.n2933 net6.n2932 0.015
R3068 net6.n2931 net6.n2930 0.015
R3069 net6.n2748 net6.n2747 0.015
R3070 net6.n2633 net6.n2632 0.015
R3071 net6.n2639 net6.n2638 0.015
R3072 net6.n2844 net6.n2843 0.015
R3073 net6.n2834 net6.n2831 0.015
R3074 net6.n2833 net6.n2832 0.015
R3075 net6.n2811 net6.n2810 0.015
R3076 net6.n2802 net6.n2801 0.015
R3077 net6.n2791 net6.n2790 0.015
R3078 net6.n2758 net6.n2757 0.015
R3079 net6.n2707 net6.n2706 0.015
R3080 net6.n2702 net6.n2701 0.015
R3081 net6.n2662 net6.n2661 0.015
R3082 net6.n2599 net6.n2598 0.015
R3083 net6.n2578 net6.n2577 0.015
R3084 net6.n2572 net6.n2571 0.015
R3085 net6.n2570 net6.n2569 0.015
R3086 net6.n2387 net6.n2386 0.015
R3087 net6.n2272 net6.n2271 0.015
R3088 net6.n2278 net6.n2277 0.015
R3089 net6.n2483 net6.n2482 0.015
R3090 net6.n2473 net6.n2470 0.015
R3091 net6.n2472 net6.n2471 0.015
R3092 net6.n2450 net6.n2449 0.015
R3093 net6.n2441 net6.n2440 0.015
R3094 net6.n2430 net6.n2429 0.015
R3095 net6.n2397 net6.n2396 0.015
R3096 net6.n2346 net6.n2345 0.015
R3097 net6.n2341 net6.n2340 0.015
R3098 net6.n2301 net6.n2300 0.015
R3099 net6.n2238 net6.n2237 0.015
R3100 net6.n2217 net6.n2216 0.015
R3101 net6.n2211 net6.n2210 0.015
R3102 net6.n2209 net6.n2208 0.015
R3103 net6.n2026 net6.n2025 0.015
R3104 net6.n1911 net6.n1910 0.015
R3105 net6.n1917 net6.n1916 0.015
R3106 net6.n2122 net6.n2121 0.015
R3107 net6.n2112 net6.n2109 0.015
R3108 net6.n2111 net6.n2110 0.015
R3109 net6.n2089 net6.n2088 0.015
R3110 net6.n2080 net6.n2079 0.015
R3111 net6.n2069 net6.n2068 0.015
R3112 net6.n2036 net6.n2035 0.015
R3113 net6.n1985 net6.n1984 0.015
R3114 net6.n1980 net6.n1979 0.015
R3115 net6.n1940 net6.n1939 0.015
R3116 net6.n1877 net6.n1876 0.015
R3117 net6.n1855 net6.n1854 0.015
R3118 net6.n1849 net6.n1848 0.015
R3119 net6.n1847 net6.n1846 0.015
R3120 net6.n1664 net6.n1663 0.015
R3121 net6.n1549 net6.n1548 0.015
R3122 net6.n1555 net6.n1554 0.015
R3123 net6.n1760 net6.n1759 0.015
R3124 net6.n1750 net6.n1747 0.015
R3125 net6.n1749 net6.n1748 0.015
R3126 net6.n1727 net6.n1726 0.015
R3127 net6.n1718 net6.n1717 0.015
R3128 net6.n1707 net6.n1706 0.015
R3129 net6.n1674 net6.n1673 0.015
R3130 net6.n1623 net6.n1622 0.015
R3131 net6.n1618 net6.n1617 0.015
R3132 net6.n1578 net6.n1577 0.015
R3133 net6.n1515 net6.n1514 0.015
R3134 net6.n1493 net6.n1492 0.015
R3135 net6.n1487 net6.n1486 0.015
R3136 net6.n1485 net6.n1484 0.015
R3137 net6.n1302 net6.n1301 0.015
R3138 net6.n1187 net6.n1186 0.015
R3139 net6.n1193 net6.n1192 0.015
R3140 net6.n1398 net6.n1397 0.015
R3141 net6.n1388 net6.n1385 0.015
R3142 net6.n1387 net6.n1386 0.015
R3143 net6.n1365 net6.n1364 0.015
R3144 net6.n1356 net6.n1355 0.015
R3145 net6.n1345 net6.n1344 0.015
R3146 net6.n1312 net6.n1311 0.015
R3147 net6.n1261 net6.n1260 0.015
R3148 net6.n1256 net6.n1255 0.015
R3149 net6.n1216 net6.n1215 0.015
R3150 net6.n1153 net6.n1152 0.015
R3151 net6.n1131 net6.n1130 0.015
R3152 net6.n1125 net6.n1124 0.015
R3153 net6.n1123 net6.n1122 0.015
R3154 net6.n940 net6.n939 0.015
R3155 net6.n825 net6.n824 0.015
R3156 net6.n831 net6.n830 0.015
R3157 net6.n1036 net6.n1035 0.015
R3158 net6.n1026 net6.n1023 0.015
R3159 net6.n1025 net6.n1024 0.015
R3160 net6.n1003 net6.n1002 0.015
R3161 net6.n994 net6.n993 0.015
R3162 net6.n983 net6.n982 0.015
R3163 net6.n950 net6.n949 0.015
R3164 net6.n899 net6.n898 0.015
R3165 net6.n894 net6.n893 0.015
R3166 net6.n854 net6.n853 0.015
R3167 net6.n791 net6.n790 0.015
R3168 net6.n769 net6.n768 0.015
R3169 net6.n763 net6.n762 0.015
R3170 net6.n761 net6.n760 0.015
R3171 net6.n578 net6.n577 0.015
R3172 net6.n463 net6.n462 0.015
R3173 net6.n469 net6.n468 0.015
R3174 net6.n674 net6.n673 0.015
R3175 net6.n664 net6.n661 0.015
R3176 net6.n663 net6.n662 0.015
R3177 net6.n641 net6.n640 0.015
R3178 net6.n632 net6.n631 0.015
R3179 net6.n621 net6.n620 0.015
R3180 net6.n588 net6.n587 0.015
R3181 net6.n537 net6.n536 0.015
R3182 net6.n532 net6.n531 0.015
R3183 net6.n492 net6.n491 0.015
R3184 net6.n429 net6.n428 0.015
R3185 net6.n407 net6.n406 0.015
R3186 net6.n401 net6.n400 0.015
R3187 net6.n399 net6.n398 0.015
R3188 net6.n216 net6.n215 0.015
R3189 net6.n101 net6.n100 0.015
R3190 net6.n107 net6.n106 0.015
R3191 net6.n312 net6.n311 0.015
R3192 net6.n302 net6.n299 0.015
R3193 net6.n301 net6.n300 0.015
R3194 net6.n279 net6.n278 0.015
R3195 net6.n270 net6.n269 0.015
R3196 net6.n259 net6.n258 0.015
R3197 net6.n226 net6.n225 0.015
R3198 net6.n175 net6.n174 0.015
R3199 net6.n170 net6.n169 0.015
R3200 net6.n130 net6.n129 0.015
R3201 net6.n67 net6.n66 0.015
R3202 net6.n3664 net6.n3661 0.013
R3203 net6.n3604 net6.n3603 0.013
R3204 net6.n3364 net6.n3361 0.013
R3205 net6.n3567 net6.n3564 0.013
R3206 net6.n3514 net6.n3511 0.013
R3207 net6.n3487 net6.n3486 0.013
R3208 net6.n3324 net6.n3323 0.013
R3209 net6.n3303 net6.n3300 0.013
R3210 net6.n3243 net6.n3242 0.013
R3211 net6.n3003 net6.n3000 0.013
R3212 net6.n3206 net6.n3203 0.013
R3213 net6.n3153 net6.n3150 0.013
R3214 net6.n3126 net6.n3125 0.013
R3215 net6.n2963 net6.n2962 0.013
R3216 net6.n2942 net6.n2939 0.013
R3217 net6.n2882 net6.n2881 0.013
R3218 net6.n2642 net6.n2639 0.013
R3219 net6.n2845 net6.n2842 0.013
R3220 net6.n2792 net6.n2789 0.013
R3221 net6.n2765 net6.n2764 0.013
R3222 net6.n2602 net6.n2601 0.013
R3223 net6.n2581 net6.n2578 0.013
R3224 net6.n2521 net6.n2520 0.013
R3225 net6.n2281 net6.n2278 0.013
R3226 net6.n2484 net6.n2481 0.013
R3227 net6.n2431 net6.n2428 0.013
R3228 net6.n2404 net6.n2403 0.013
R3229 net6.n2241 net6.n2240 0.013
R3230 net6.n2220 net6.n2217 0.013
R3231 net6.n2160 net6.n2159 0.013
R3232 net6.n1920 net6.n1917 0.013
R3233 net6.n2123 net6.n2120 0.013
R3234 net6.n2070 net6.n2067 0.013
R3235 net6.n2043 net6.n2042 0.013
R3236 net6.n1880 net6.n1879 0.013
R3237 net6.n1858 net6.n1855 0.013
R3238 net6.n1798 net6.n1797 0.013
R3239 net6.n1558 net6.n1555 0.013
R3240 net6.n1761 net6.n1758 0.013
R3241 net6.n1708 net6.n1705 0.013
R3242 net6.n1681 net6.n1680 0.013
R3243 net6.n1518 net6.n1517 0.013
R3244 net6.n1496 net6.n1493 0.013
R3245 net6.n1436 net6.n1435 0.013
R3246 net6.n1196 net6.n1193 0.013
R3247 net6.n1399 net6.n1396 0.013
R3248 net6.n1346 net6.n1343 0.013
R3249 net6.n1319 net6.n1318 0.013
R3250 net6.n1156 net6.n1155 0.013
R3251 net6.n1134 net6.n1131 0.013
R3252 net6.n1074 net6.n1073 0.013
R3253 net6.n834 net6.n831 0.013
R3254 net6.n1037 net6.n1034 0.013
R3255 net6.n984 net6.n981 0.013
R3256 net6.n957 net6.n956 0.013
R3257 net6.n794 net6.n793 0.013
R3258 net6.n772 net6.n769 0.013
R3259 net6.n712 net6.n711 0.013
R3260 net6.n472 net6.n469 0.013
R3261 net6.n675 net6.n672 0.013
R3262 net6.n622 net6.n619 0.013
R3263 net6.n595 net6.n594 0.013
R3264 net6.n432 net6.n431 0.013
R3265 net6.n410 net6.n407 0.013
R3266 net6.n350 net6.n349 0.013
R3267 net6.n110 net6.n107 0.013
R3268 net6.n313 net6.n310 0.013
R3269 net6.n260 net6.n257 0.013
R3270 net6.n233 net6.n232 0.013
R3271 net6.n70 net6.n69 0.013
R3272 net6.n3652 net6.n3651 0.011
R3273 net6.n3622 net6.n3621 0.011
R3274 net6.n3457 net6.n3456 0.011
R3275 net6.n3349 net6.n3348 0.011
R3276 net6.n3291 net6.n3290 0.011
R3277 net6.n3261 net6.n3260 0.011
R3278 net6.n3096 net6.n3095 0.011
R3279 net6.n2988 net6.n2987 0.011
R3280 net6.n2930 net6.n2929 0.011
R3281 net6.n2900 net6.n2899 0.011
R3282 net6.n2735 net6.n2734 0.011
R3283 net6.n2627 net6.n2626 0.011
R3284 net6.n2569 net6.n2568 0.011
R3285 net6.n2539 net6.n2538 0.011
R3286 net6.n2374 net6.n2373 0.011
R3287 net6.n2266 net6.n2265 0.011
R3288 net6.n2208 net6.n2207 0.011
R3289 net6.n2178 net6.n2177 0.011
R3290 net6.n2013 net6.n2012 0.011
R3291 net6.n1905 net6.n1904 0.011
R3292 net6.n1846 net6.n1845 0.011
R3293 net6.n1816 net6.n1815 0.011
R3294 net6.n1651 net6.n1650 0.011
R3295 net6.n1543 net6.n1542 0.011
R3296 net6.n1484 net6.n1483 0.011
R3297 net6.n1454 net6.n1453 0.011
R3298 net6.n1289 net6.n1288 0.011
R3299 net6.n1181 net6.n1180 0.011
R3300 net6.n1122 net6.n1121 0.011
R3301 net6.n1092 net6.n1091 0.011
R3302 net6.n927 net6.n926 0.011
R3303 net6.n819 net6.n818 0.011
R3304 net6.n760 net6.n759 0.011
R3305 net6.n730 net6.n729 0.011
R3306 net6.n565 net6.n564 0.011
R3307 net6.n457 net6.n456 0.011
R3308 net6.n398 net6.n397 0.011
R3309 net6.n368 net6.n367 0.011
R3310 net6.n203 net6.n202 0.011
R3311 net6.n95 net6.n94 0.011
R3312 net6.n51 net6.n50 0.01
R3313 net6.n58 net6.n52 0.01
R3314 net6.n3660 net6.n3658 0.009
R3315 net6.n3632 net6.n3631 0.009
R3316 net6.n3406 net6.n3405 0.009
R3317 net6.n3336 net6.n3335 0.009
R3318 net6.n3367 net6.n3366 0.009
R3319 net6.n3677 net6.n3676 0.009
R3320 net6.n3535 net6.n3534 0.009
R3321 net6.n3518 net6.n3517 0.009
R3322 net6.n3410 net6.n3398 0.009
R3323 net6.n3395 net6.n3394 0.009
R3324 net6.n3326 net6.n3325 0.009
R3325 net6.n3568 net6.n3563 0.009
R3326 net6.n3562 net6.n3561 0.009
R3327 net6.n3557 net6.n3552 0.009
R3328 net6.n3551 net6.n3550 0.009
R3329 net6.n3526 net6.n3521 0.009
R3330 net6.n3520 net6.n3519 0.009
R3331 net6.n3515 net6.n3510 0.009
R3332 net6.n3509 net6.n3508 0.009
R3333 net6.n3482 net6.n3432 0.009
R3334 net6.n3431 net6.n3430 0.009
R3335 net6.n3426 net6.n3421 0.009
R3336 net6.n3420 net6.n3419 0.009
R3337 net6.n3387 net6.n3382 0.009
R3338 net6.n3381 net6.n3380 0.009
R3339 net6.n3376 net6.n3375 0.009
R3340 net6.n3374 net6.n3373 0.009
R3341 net6.n3299 net6.n3297 0.009
R3342 net6.n3271 net6.n3270 0.009
R3343 net6.n3045 net6.n3044 0.009
R3344 net6.n2975 net6.n2974 0.009
R3345 net6.n3006 net6.n3005 0.009
R3346 net6.n3316 net6.n3315 0.009
R3347 net6.n3174 net6.n3173 0.009
R3348 net6.n3157 net6.n3156 0.009
R3349 net6.n3049 net6.n3037 0.009
R3350 net6.n3034 net6.n3033 0.009
R3351 net6.n2965 net6.n2964 0.009
R3352 net6.n3207 net6.n3202 0.009
R3353 net6.n3201 net6.n3200 0.009
R3354 net6.n3196 net6.n3191 0.009
R3355 net6.n3190 net6.n3189 0.009
R3356 net6.n3165 net6.n3160 0.009
R3357 net6.n3159 net6.n3158 0.009
R3358 net6.n3154 net6.n3149 0.009
R3359 net6.n3148 net6.n3147 0.009
R3360 net6.n3121 net6.n3071 0.009
R3361 net6.n3070 net6.n3069 0.009
R3362 net6.n3065 net6.n3060 0.009
R3363 net6.n3059 net6.n3058 0.009
R3364 net6.n3026 net6.n3021 0.009
R3365 net6.n3020 net6.n3019 0.009
R3366 net6.n3015 net6.n3014 0.009
R3367 net6.n3013 net6.n3012 0.009
R3368 net6.n2938 net6.n2936 0.009
R3369 net6.n2910 net6.n2909 0.009
R3370 net6.n2684 net6.n2683 0.009
R3371 net6.n2614 net6.n2613 0.009
R3372 net6.n2645 net6.n2644 0.009
R3373 net6.n2955 net6.n2954 0.009
R3374 net6.n2813 net6.n2812 0.009
R3375 net6.n2796 net6.n2795 0.009
R3376 net6.n2688 net6.n2676 0.009
R3377 net6.n2673 net6.n2672 0.009
R3378 net6.n2604 net6.n2603 0.009
R3379 net6.n2846 net6.n2841 0.009
R3380 net6.n2840 net6.n2839 0.009
R3381 net6.n2835 net6.n2830 0.009
R3382 net6.n2829 net6.n2828 0.009
R3383 net6.n2804 net6.n2799 0.009
R3384 net6.n2798 net6.n2797 0.009
R3385 net6.n2793 net6.n2788 0.009
R3386 net6.n2787 net6.n2786 0.009
R3387 net6.n2760 net6.n2710 0.009
R3388 net6.n2709 net6.n2708 0.009
R3389 net6.n2704 net6.n2699 0.009
R3390 net6.n2698 net6.n2697 0.009
R3391 net6.n2665 net6.n2660 0.009
R3392 net6.n2659 net6.n2658 0.009
R3393 net6.n2654 net6.n2653 0.009
R3394 net6.n2652 net6.n2651 0.009
R3395 net6.n2577 net6.n2575 0.009
R3396 net6.n2549 net6.n2548 0.009
R3397 net6.n2323 net6.n2322 0.009
R3398 net6.n2253 net6.n2252 0.009
R3399 net6.n2284 net6.n2283 0.009
R3400 net6.n2594 net6.n2593 0.009
R3401 net6.n2452 net6.n2451 0.009
R3402 net6.n2435 net6.n2434 0.009
R3403 net6.n2327 net6.n2315 0.009
R3404 net6.n2312 net6.n2311 0.009
R3405 net6.n2243 net6.n2242 0.009
R3406 net6.n2485 net6.n2480 0.009
R3407 net6.n2479 net6.n2478 0.009
R3408 net6.n2474 net6.n2469 0.009
R3409 net6.n2468 net6.n2467 0.009
R3410 net6.n2443 net6.n2438 0.009
R3411 net6.n2437 net6.n2436 0.009
R3412 net6.n2432 net6.n2427 0.009
R3413 net6.n2426 net6.n2425 0.009
R3414 net6.n2399 net6.n2349 0.009
R3415 net6.n2348 net6.n2347 0.009
R3416 net6.n2343 net6.n2338 0.009
R3417 net6.n2337 net6.n2336 0.009
R3418 net6.n2304 net6.n2299 0.009
R3419 net6.n2298 net6.n2297 0.009
R3420 net6.n2293 net6.n2292 0.009
R3421 net6.n2291 net6.n2290 0.009
R3422 net6.n2216 net6.n2214 0.009
R3423 net6.n2188 net6.n2187 0.009
R3424 net6.n1962 net6.n1961 0.009
R3425 net6.n1892 net6.n1891 0.009
R3426 net6.n1923 net6.n1922 0.009
R3427 net6.n2233 net6.n2232 0.009
R3428 net6.n2091 net6.n2090 0.009
R3429 net6.n2074 net6.n2073 0.009
R3430 net6.n1966 net6.n1954 0.009
R3431 net6.n1951 net6.n1950 0.009
R3432 net6.n1882 net6.n1881 0.009
R3433 net6.n2124 net6.n2119 0.009
R3434 net6.n2118 net6.n2117 0.009
R3435 net6.n2113 net6.n2108 0.009
R3436 net6.n2107 net6.n2106 0.009
R3437 net6.n2082 net6.n2077 0.009
R3438 net6.n2076 net6.n2075 0.009
R3439 net6.n2071 net6.n2066 0.009
R3440 net6.n2065 net6.n2064 0.009
R3441 net6.n2038 net6.n1988 0.009
R3442 net6.n1987 net6.n1986 0.009
R3443 net6.n1982 net6.n1977 0.009
R3444 net6.n1976 net6.n1975 0.009
R3445 net6.n1943 net6.n1938 0.009
R3446 net6.n1937 net6.n1936 0.009
R3447 net6.n1932 net6.n1931 0.009
R3448 net6.n1930 net6.n1929 0.009
R3449 net6.n1854 net6.n1852 0.009
R3450 net6.n1826 net6.n1825 0.009
R3451 net6.n1600 net6.n1599 0.009
R3452 net6.n1530 net6.n1529 0.009
R3453 net6.n1561 net6.n1560 0.009
R3454 net6.n1871 net6.n1870 0.009
R3455 net6.n1729 net6.n1728 0.009
R3456 net6.n1712 net6.n1711 0.009
R3457 net6.n1604 net6.n1592 0.009
R3458 net6.n1589 net6.n1588 0.009
R3459 net6.n1520 net6.n1519 0.009
R3460 net6.n1762 net6.n1757 0.009
R3461 net6.n1756 net6.n1755 0.009
R3462 net6.n1751 net6.n1746 0.009
R3463 net6.n1745 net6.n1744 0.009
R3464 net6.n1720 net6.n1715 0.009
R3465 net6.n1714 net6.n1713 0.009
R3466 net6.n1709 net6.n1704 0.009
R3467 net6.n1703 net6.n1702 0.009
R3468 net6.n1676 net6.n1626 0.009
R3469 net6.n1625 net6.n1624 0.009
R3470 net6.n1620 net6.n1615 0.009
R3471 net6.n1614 net6.n1613 0.009
R3472 net6.n1581 net6.n1576 0.009
R3473 net6.n1575 net6.n1574 0.009
R3474 net6.n1570 net6.n1569 0.009
R3475 net6.n1568 net6.n1567 0.009
R3476 net6.n1492 net6.n1490 0.009
R3477 net6.n1464 net6.n1463 0.009
R3478 net6.n1238 net6.n1237 0.009
R3479 net6.n1168 net6.n1167 0.009
R3480 net6.n1199 net6.n1198 0.009
R3481 net6.n1509 net6.n1508 0.009
R3482 net6.n1367 net6.n1366 0.009
R3483 net6.n1350 net6.n1349 0.009
R3484 net6.n1242 net6.n1230 0.009
R3485 net6.n1227 net6.n1226 0.009
R3486 net6.n1158 net6.n1157 0.009
R3487 net6.n1400 net6.n1395 0.009
R3488 net6.n1394 net6.n1393 0.009
R3489 net6.n1389 net6.n1384 0.009
R3490 net6.n1383 net6.n1382 0.009
R3491 net6.n1358 net6.n1353 0.009
R3492 net6.n1352 net6.n1351 0.009
R3493 net6.n1347 net6.n1342 0.009
R3494 net6.n1341 net6.n1340 0.009
R3495 net6.n1314 net6.n1264 0.009
R3496 net6.n1263 net6.n1262 0.009
R3497 net6.n1258 net6.n1253 0.009
R3498 net6.n1252 net6.n1251 0.009
R3499 net6.n1219 net6.n1214 0.009
R3500 net6.n1213 net6.n1212 0.009
R3501 net6.n1208 net6.n1207 0.009
R3502 net6.n1206 net6.n1205 0.009
R3503 net6.n1130 net6.n1128 0.009
R3504 net6.n1102 net6.n1101 0.009
R3505 net6.n876 net6.n875 0.009
R3506 net6.n806 net6.n805 0.009
R3507 net6.n837 net6.n836 0.009
R3508 net6.n1147 net6.n1146 0.009
R3509 net6.n1005 net6.n1004 0.009
R3510 net6.n988 net6.n987 0.009
R3511 net6.n880 net6.n868 0.009
R3512 net6.n865 net6.n864 0.009
R3513 net6.n796 net6.n795 0.009
R3514 net6.n1038 net6.n1033 0.009
R3515 net6.n1032 net6.n1031 0.009
R3516 net6.n1027 net6.n1022 0.009
R3517 net6.n1021 net6.n1020 0.009
R3518 net6.n996 net6.n991 0.009
R3519 net6.n990 net6.n989 0.009
R3520 net6.n985 net6.n980 0.009
R3521 net6.n979 net6.n978 0.009
R3522 net6.n952 net6.n902 0.009
R3523 net6.n901 net6.n900 0.009
R3524 net6.n896 net6.n891 0.009
R3525 net6.n890 net6.n889 0.009
R3526 net6.n857 net6.n852 0.009
R3527 net6.n851 net6.n850 0.009
R3528 net6.n846 net6.n845 0.009
R3529 net6.n844 net6.n843 0.009
R3530 net6.n768 net6.n766 0.009
R3531 net6.n740 net6.n739 0.009
R3532 net6.n514 net6.n513 0.009
R3533 net6.n444 net6.n443 0.009
R3534 net6.n475 net6.n474 0.009
R3535 net6.n785 net6.n784 0.009
R3536 net6.n643 net6.n642 0.009
R3537 net6.n626 net6.n625 0.009
R3538 net6.n518 net6.n506 0.009
R3539 net6.n503 net6.n502 0.009
R3540 net6.n434 net6.n433 0.009
R3541 net6.n676 net6.n671 0.009
R3542 net6.n670 net6.n669 0.009
R3543 net6.n665 net6.n660 0.009
R3544 net6.n659 net6.n658 0.009
R3545 net6.n634 net6.n629 0.009
R3546 net6.n628 net6.n627 0.009
R3547 net6.n623 net6.n618 0.009
R3548 net6.n617 net6.n616 0.009
R3549 net6.n590 net6.n540 0.009
R3550 net6.n539 net6.n538 0.009
R3551 net6.n534 net6.n529 0.009
R3552 net6.n528 net6.n527 0.009
R3553 net6.n495 net6.n490 0.009
R3554 net6.n489 net6.n488 0.009
R3555 net6.n484 net6.n483 0.009
R3556 net6.n482 net6.n481 0.009
R3557 net6.n406 net6.n404 0.009
R3558 net6.n378 net6.n377 0.009
R3559 net6.n152 net6.n151 0.009
R3560 net6.n82 net6.n81 0.009
R3561 net6.n113 net6.n112 0.009
R3562 net6.n423 net6.n422 0.009
R3563 net6.n281 net6.n280 0.009
R3564 net6.n264 net6.n263 0.009
R3565 net6.n156 net6.n144 0.009
R3566 net6.n141 net6.n140 0.009
R3567 net6.n72 net6.n71 0.009
R3568 net6.n314 net6.n309 0.009
R3569 net6.n308 net6.n307 0.009
R3570 net6.n303 net6.n298 0.009
R3571 net6.n297 net6.n296 0.009
R3572 net6.n272 net6.n267 0.009
R3573 net6.n266 net6.n265 0.009
R3574 net6.n261 net6.n256 0.009
R3575 net6.n255 net6.n254 0.009
R3576 net6.n228 net6.n178 0.009
R3577 net6.n177 net6.n176 0.009
R3578 net6.n172 net6.n167 0.009
R3579 net6.n166 net6.n165 0.009
R3580 net6.n133 net6.n128 0.009
R3581 net6.n127 net6.n126 0.009
R3582 net6.n122 net6.n121 0.009
R3583 net6.n120 net6.n119 0.009
R3584 net6.n11 net6.n10 0.007
R3585 net6.n5 net6.n4 0.007
R3586 net6.n15 net6.n14 0.007
R3587 net6.n3667 net6.n3666 0.007
R3588 net6.n3657 net6.n3656 0.007
R3589 net6.n3637 net6.n3636 0.007
R3590 net6.n3631 net6.n3630 0.007
R3591 net6.n3608 net6.n3607 0.007
R3592 net6.n3436 net6.n3435 0.007
R3593 net6.n3445 net6.n3444 0.007
R3594 net6.n3467 net6.n3466 0.007
R3595 net6.n3462 net6.n3461 0.007
R3596 net6.n3460 net6.n3459 0.007
R3597 net6.n3456 net6.n3455 0.007
R3598 net6.n3407 net6.n3406 0.007
R3599 net6.n3360 net6.n3358 0.007
R3600 net6.n3673 net6.n3672 0.007
R3601 net6.n3560 net6.n3559 0.007
R3602 net6.n3543 net6.n3538 0.007
R3603 net6.n3542 net6.n3541 0.007
R3604 net6.n3494 net6.n3493 0.007
R3605 net6.n3496 net6.n3495 0.007
R3606 net6.n3489 net6.n3488 0.007
R3607 net6.n3425 net6.n3422 0.007
R3608 net6.n3418 net6.n3417 0.007
R3609 net6.n3416 net6.n3415 0.007
R3610 net6.n3306 net6.n3305 0.007
R3611 net6.n3296 net6.n3295 0.007
R3612 net6.n3276 net6.n3275 0.007
R3613 net6.n3270 net6.n3269 0.007
R3614 net6.n3247 net6.n3246 0.007
R3615 net6.n3075 net6.n3074 0.007
R3616 net6.n3084 net6.n3083 0.007
R3617 net6.n3106 net6.n3105 0.007
R3618 net6.n3101 net6.n3100 0.007
R3619 net6.n3099 net6.n3098 0.007
R3620 net6.n3095 net6.n3094 0.007
R3621 net6.n3046 net6.n3045 0.007
R3622 net6.n2999 net6.n2997 0.007
R3623 net6.n3312 net6.n3311 0.007
R3624 net6.n3199 net6.n3198 0.007
R3625 net6.n3182 net6.n3177 0.007
R3626 net6.n3181 net6.n3180 0.007
R3627 net6.n3133 net6.n3132 0.007
R3628 net6.n3135 net6.n3134 0.007
R3629 net6.n3128 net6.n3127 0.007
R3630 net6.n3064 net6.n3061 0.007
R3631 net6.n3057 net6.n3056 0.007
R3632 net6.n3055 net6.n3054 0.007
R3633 net6.n2945 net6.n2944 0.007
R3634 net6.n2935 net6.n2934 0.007
R3635 net6.n2915 net6.n2914 0.007
R3636 net6.n2909 net6.n2908 0.007
R3637 net6.n2886 net6.n2885 0.007
R3638 net6.n2714 net6.n2713 0.007
R3639 net6.n2723 net6.n2722 0.007
R3640 net6.n2745 net6.n2744 0.007
R3641 net6.n2740 net6.n2739 0.007
R3642 net6.n2738 net6.n2737 0.007
R3643 net6.n2734 net6.n2733 0.007
R3644 net6.n2685 net6.n2684 0.007
R3645 net6.n2638 net6.n2636 0.007
R3646 net6.n2951 net6.n2950 0.007
R3647 net6.n2838 net6.n2837 0.007
R3648 net6.n2821 net6.n2816 0.007
R3649 net6.n2820 net6.n2819 0.007
R3650 net6.n2772 net6.n2771 0.007
R3651 net6.n2774 net6.n2773 0.007
R3652 net6.n2767 net6.n2766 0.007
R3653 net6.n2703 net6.n2700 0.007
R3654 net6.n2696 net6.n2695 0.007
R3655 net6.n2694 net6.n2693 0.007
R3656 net6.n2584 net6.n2583 0.007
R3657 net6.n2574 net6.n2573 0.007
R3658 net6.n2554 net6.n2553 0.007
R3659 net6.n2548 net6.n2547 0.007
R3660 net6.n2525 net6.n2524 0.007
R3661 net6.n2353 net6.n2352 0.007
R3662 net6.n2362 net6.n2361 0.007
R3663 net6.n2384 net6.n2383 0.007
R3664 net6.n2379 net6.n2378 0.007
R3665 net6.n2377 net6.n2376 0.007
R3666 net6.n2373 net6.n2372 0.007
R3667 net6.n2324 net6.n2323 0.007
R3668 net6.n2277 net6.n2275 0.007
R3669 net6.n2590 net6.n2589 0.007
R3670 net6.n2477 net6.n2476 0.007
R3671 net6.n2460 net6.n2455 0.007
R3672 net6.n2459 net6.n2458 0.007
R3673 net6.n2411 net6.n2410 0.007
R3674 net6.n2413 net6.n2412 0.007
R3675 net6.n2406 net6.n2405 0.007
R3676 net6.n2342 net6.n2339 0.007
R3677 net6.n2335 net6.n2334 0.007
R3678 net6.n2333 net6.n2332 0.007
R3679 net6.n2223 net6.n2222 0.007
R3680 net6.n2213 net6.n2212 0.007
R3681 net6.n2193 net6.n2192 0.007
R3682 net6.n2187 net6.n2186 0.007
R3683 net6.n2164 net6.n2163 0.007
R3684 net6.n1992 net6.n1991 0.007
R3685 net6.n2001 net6.n2000 0.007
R3686 net6.n2023 net6.n2022 0.007
R3687 net6.n2018 net6.n2017 0.007
R3688 net6.n2016 net6.n2015 0.007
R3689 net6.n2012 net6.n2011 0.007
R3690 net6.n1963 net6.n1962 0.007
R3691 net6.n1916 net6.n1914 0.007
R3692 net6.n2229 net6.n2228 0.007
R3693 net6.n2116 net6.n2115 0.007
R3694 net6.n2099 net6.n2094 0.007
R3695 net6.n2098 net6.n2097 0.007
R3696 net6.n2050 net6.n2049 0.007
R3697 net6.n2052 net6.n2051 0.007
R3698 net6.n2045 net6.n2044 0.007
R3699 net6.n1981 net6.n1978 0.007
R3700 net6.n1974 net6.n1973 0.007
R3701 net6.n1972 net6.n1971 0.007
R3702 net6.n1861 net6.n1860 0.007
R3703 net6.n1851 net6.n1850 0.007
R3704 net6.n1831 net6.n1830 0.007
R3705 net6.n1825 net6.n1824 0.007
R3706 net6.n1802 net6.n1801 0.007
R3707 net6.n1630 net6.n1629 0.007
R3708 net6.n1639 net6.n1638 0.007
R3709 net6.n1661 net6.n1660 0.007
R3710 net6.n1656 net6.n1655 0.007
R3711 net6.n1654 net6.n1653 0.007
R3712 net6.n1650 net6.n1649 0.007
R3713 net6.n1601 net6.n1600 0.007
R3714 net6.n1554 net6.n1552 0.007
R3715 net6.n1867 net6.n1866 0.007
R3716 net6.n1754 net6.n1753 0.007
R3717 net6.n1737 net6.n1732 0.007
R3718 net6.n1736 net6.n1735 0.007
R3719 net6.n1688 net6.n1687 0.007
R3720 net6.n1690 net6.n1689 0.007
R3721 net6.n1683 net6.n1682 0.007
R3722 net6.n1619 net6.n1616 0.007
R3723 net6.n1612 net6.n1611 0.007
R3724 net6.n1610 net6.n1609 0.007
R3725 net6.n1499 net6.n1498 0.007
R3726 net6.n1489 net6.n1488 0.007
R3727 net6.n1469 net6.n1468 0.007
R3728 net6.n1463 net6.n1462 0.007
R3729 net6.n1440 net6.n1439 0.007
R3730 net6.n1268 net6.n1267 0.007
R3731 net6.n1277 net6.n1276 0.007
R3732 net6.n1299 net6.n1298 0.007
R3733 net6.n1294 net6.n1293 0.007
R3734 net6.n1292 net6.n1291 0.007
R3735 net6.n1288 net6.n1287 0.007
R3736 net6.n1239 net6.n1238 0.007
R3737 net6.n1192 net6.n1190 0.007
R3738 net6.n1505 net6.n1504 0.007
R3739 net6.n1392 net6.n1391 0.007
R3740 net6.n1375 net6.n1370 0.007
R3741 net6.n1374 net6.n1373 0.007
R3742 net6.n1326 net6.n1325 0.007
R3743 net6.n1328 net6.n1327 0.007
R3744 net6.n1321 net6.n1320 0.007
R3745 net6.n1257 net6.n1254 0.007
R3746 net6.n1250 net6.n1249 0.007
R3747 net6.n1248 net6.n1247 0.007
R3748 net6.n1137 net6.n1136 0.007
R3749 net6.n1127 net6.n1126 0.007
R3750 net6.n1107 net6.n1106 0.007
R3751 net6.n1101 net6.n1100 0.007
R3752 net6.n1078 net6.n1077 0.007
R3753 net6.n906 net6.n905 0.007
R3754 net6.n915 net6.n914 0.007
R3755 net6.n937 net6.n936 0.007
R3756 net6.n932 net6.n931 0.007
R3757 net6.n930 net6.n929 0.007
R3758 net6.n926 net6.n925 0.007
R3759 net6.n877 net6.n876 0.007
R3760 net6.n830 net6.n828 0.007
R3761 net6.n1143 net6.n1142 0.007
R3762 net6.n1030 net6.n1029 0.007
R3763 net6.n1013 net6.n1008 0.007
R3764 net6.n1012 net6.n1011 0.007
R3765 net6.n964 net6.n963 0.007
R3766 net6.n966 net6.n965 0.007
R3767 net6.n959 net6.n958 0.007
R3768 net6.n895 net6.n892 0.007
R3769 net6.n888 net6.n887 0.007
R3770 net6.n886 net6.n885 0.007
R3771 net6.n775 net6.n774 0.007
R3772 net6.n765 net6.n764 0.007
R3773 net6.n745 net6.n744 0.007
R3774 net6.n739 net6.n738 0.007
R3775 net6.n716 net6.n715 0.007
R3776 net6.n544 net6.n543 0.007
R3777 net6.n553 net6.n552 0.007
R3778 net6.n575 net6.n574 0.007
R3779 net6.n570 net6.n569 0.007
R3780 net6.n568 net6.n567 0.007
R3781 net6.n564 net6.n563 0.007
R3782 net6.n515 net6.n514 0.007
R3783 net6.n468 net6.n466 0.007
R3784 net6.n781 net6.n780 0.007
R3785 net6.n668 net6.n667 0.007
R3786 net6.n651 net6.n646 0.007
R3787 net6.n650 net6.n649 0.007
R3788 net6.n602 net6.n601 0.007
R3789 net6.n604 net6.n603 0.007
R3790 net6.n597 net6.n596 0.007
R3791 net6.n533 net6.n530 0.007
R3792 net6.n526 net6.n525 0.007
R3793 net6.n524 net6.n523 0.007
R3794 net6.n413 net6.n412 0.007
R3795 net6.n403 net6.n402 0.007
R3796 net6.n383 net6.n382 0.007
R3797 net6.n377 net6.n376 0.007
R3798 net6.n354 net6.n353 0.007
R3799 net6.n182 net6.n181 0.007
R3800 net6.n191 net6.n190 0.007
R3801 net6.n213 net6.n212 0.007
R3802 net6.n208 net6.n207 0.007
R3803 net6.n206 net6.n205 0.007
R3804 net6.n202 net6.n201 0.007
R3805 net6.n153 net6.n152 0.007
R3806 net6.n106 net6.n104 0.007
R3807 net6.n419 net6.n418 0.007
R3808 net6.n306 net6.n305 0.007
R3809 net6.n289 net6.n284 0.007
R3810 net6.n288 net6.n287 0.007
R3811 net6.n240 net6.n239 0.007
R3812 net6.n242 net6.n241 0.007
R3813 net6.n235 net6.n234 0.007
R3814 net6.n171 net6.n168 0.007
R3815 net6.n164 net6.n163 0.007
R3816 net6.n162 net6.n161 0.007
R3817 net6.n3654 net6.n3653 0.005
R3818 net6.n3651 net6.n3649 0.005
R3819 net6.n3634 net6.n3633 0.005
R3820 net6.n3625 net6.n3624 0.005
R3821 net6.n3623 net6.n3622 0.005
R3822 net6.n3620 net6.n3619 0.005
R3823 net6.n3619 net6.n3616 0.005
R3824 net6.n3615 net6.n3614 0.005
R3825 net6.n3590 net6.n3589 0.005
R3826 net6.n3434 net6.n3433 0.005
R3827 net6.n3401 net6.n3400 0.005
R3828 net6.n3330 net6.n3329 0.005
R3829 net6.n3357 net6.n3356 0.005
R3830 net6.n3535 net6.n3529 0.005
R3831 net6.n3531 net6.n3530 0.005
R3832 net6.n3525 net6.n3522 0.005
R3833 net6.n3498 net6.n3497 0.005
R3834 net6.n3410 net6.n3409 0.005
R3835 net6.n3319 net6.n3318 0.005
R3836 net6.n3563 net6.n3562 0.005
R3837 net6.n3552 net6.n3551 0.005
R3838 net6.n3521 net6.n3520 0.005
R3839 net6.n3510 net6.n3509 0.005
R3840 net6.n3432 net6.n3431 0.005
R3841 net6.n3421 net6.n3420 0.005
R3842 net6.n3382 net6.n3381 0.005
R3843 net6.n3375 net6.n3374 0.005
R3844 net6.n3293 net6.n3292 0.005
R3845 net6.n3290 net6.n3288 0.005
R3846 net6.n3273 net6.n3272 0.005
R3847 net6.n3264 net6.n3263 0.005
R3848 net6.n3262 net6.n3261 0.005
R3849 net6.n3259 net6.n3258 0.005
R3850 net6.n3258 net6.n3255 0.005
R3851 net6.n3254 net6.n3253 0.005
R3852 net6.n3229 net6.n3228 0.005
R3853 net6.n3073 net6.n3072 0.005
R3854 net6.n3040 net6.n3039 0.005
R3855 net6.n2969 net6.n2968 0.005
R3856 net6.n2996 net6.n2995 0.005
R3857 net6.n3174 net6.n3168 0.005
R3858 net6.n3170 net6.n3169 0.005
R3859 net6.n3164 net6.n3161 0.005
R3860 net6.n3137 net6.n3136 0.005
R3861 net6.n3049 net6.n3048 0.005
R3862 net6.n2958 net6.n2957 0.005
R3863 net6.n3202 net6.n3201 0.005
R3864 net6.n3191 net6.n3190 0.005
R3865 net6.n3160 net6.n3159 0.005
R3866 net6.n3149 net6.n3148 0.005
R3867 net6.n3071 net6.n3070 0.005
R3868 net6.n3060 net6.n3059 0.005
R3869 net6.n3021 net6.n3020 0.005
R3870 net6.n3014 net6.n3013 0.005
R3871 net6.n2932 net6.n2931 0.005
R3872 net6.n2929 net6.n2927 0.005
R3873 net6.n2912 net6.n2911 0.005
R3874 net6.n2903 net6.n2902 0.005
R3875 net6.n2901 net6.n2900 0.005
R3876 net6.n2898 net6.n2897 0.005
R3877 net6.n2897 net6.n2894 0.005
R3878 net6.n2893 net6.n2892 0.005
R3879 net6.n2868 net6.n2867 0.005
R3880 net6.n2712 net6.n2711 0.005
R3881 net6.n2679 net6.n2678 0.005
R3882 net6.n2608 net6.n2607 0.005
R3883 net6.n2635 net6.n2634 0.005
R3884 net6.n2813 net6.n2807 0.005
R3885 net6.n2809 net6.n2808 0.005
R3886 net6.n2803 net6.n2800 0.005
R3887 net6.n2776 net6.n2775 0.005
R3888 net6.n2688 net6.n2687 0.005
R3889 net6.n2597 net6.n2596 0.005
R3890 net6.n2841 net6.n2840 0.005
R3891 net6.n2830 net6.n2829 0.005
R3892 net6.n2799 net6.n2798 0.005
R3893 net6.n2788 net6.n2787 0.005
R3894 net6.n2710 net6.n2709 0.005
R3895 net6.n2699 net6.n2698 0.005
R3896 net6.n2660 net6.n2659 0.005
R3897 net6.n2653 net6.n2652 0.005
R3898 net6.n2571 net6.n2570 0.005
R3899 net6.n2568 net6.n2566 0.005
R3900 net6.n2551 net6.n2550 0.005
R3901 net6.n2542 net6.n2541 0.005
R3902 net6.n2540 net6.n2539 0.005
R3903 net6.n2537 net6.n2536 0.005
R3904 net6.n2536 net6.n2533 0.005
R3905 net6.n2532 net6.n2531 0.005
R3906 net6.n2507 net6.n2506 0.005
R3907 net6.n2351 net6.n2350 0.005
R3908 net6.n2318 net6.n2317 0.005
R3909 net6.n2247 net6.n2246 0.005
R3910 net6.n2274 net6.n2273 0.005
R3911 net6.n2452 net6.n2446 0.005
R3912 net6.n2448 net6.n2447 0.005
R3913 net6.n2442 net6.n2439 0.005
R3914 net6.n2415 net6.n2414 0.005
R3915 net6.n2327 net6.n2326 0.005
R3916 net6.n2236 net6.n2235 0.005
R3917 net6.n2480 net6.n2479 0.005
R3918 net6.n2469 net6.n2468 0.005
R3919 net6.n2438 net6.n2437 0.005
R3920 net6.n2427 net6.n2426 0.005
R3921 net6.n2349 net6.n2348 0.005
R3922 net6.n2338 net6.n2337 0.005
R3923 net6.n2299 net6.n2298 0.005
R3924 net6.n2292 net6.n2291 0.005
R3925 net6.n2210 net6.n2209 0.005
R3926 net6.n2207 net6.n2205 0.005
R3927 net6.n2190 net6.n2189 0.005
R3928 net6.n2181 net6.n2180 0.005
R3929 net6.n2179 net6.n2178 0.005
R3930 net6.n2176 net6.n2175 0.005
R3931 net6.n2175 net6.n2172 0.005
R3932 net6.n2171 net6.n2170 0.005
R3933 net6.n2146 net6.n2145 0.005
R3934 net6.n1990 net6.n1989 0.005
R3935 net6.n1957 net6.n1956 0.005
R3936 net6.n1886 net6.n1885 0.005
R3937 net6.n1913 net6.n1912 0.005
R3938 net6.n2091 net6.n2085 0.005
R3939 net6.n2087 net6.n2086 0.005
R3940 net6.n2081 net6.n2078 0.005
R3941 net6.n2054 net6.n2053 0.005
R3942 net6.n1966 net6.n1965 0.005
R3943 net6.n1875 net6.n1874 0.005
R3944 net6.n2119 net6.n2118 0.005
R3945 net6.n2108 net6.n2107 0.005
R3946 net6.n2077 net6.n2076 0.005
R3947 net6.n2066 net6.n2065 0.005
R3948 net6.n1988 net6.n1987 0.005
R3949 net6.n1977 net6.n1976 0.005
R3950 net6.n1938 net6.n1937 0.005
R3951 net6.n1931 net6.n1930 0.005
R3952 net6.n1848 net6.n1847 0.005
R3953 net6.n1845 net6.n1843 0.005
R3954 net6.n1828 net6.n1827 0.005
R3955 net6.n1819 net6.n1818 0.005
R3956 net6.n1817 net6.n1816 0.005
R3957 net6.n1814 net6.n1813 0.005
R3958 net6.n1813 net6.n1810 0.005
R3959 net6.n1809 net6.n1808 0.005
R3960 net6.n1784 net6.n1783 0.005
R3961 net6.n1628 net6.n1627 0.005
R3962 net6.n1595 net6.n1594 0.005
R3963 net6.n1524 net6.n1523 0.005
R3964 net6.n1551 net6.n1550 0.005
R3965 net6.n1729 net6.n1723 0.005
R3966 net6.n1725 net6.n1724 0.005
R3967 net6.n1719 net6.n1716 0.005
R3968 net6.n1692 net6.n1691 0.005
R3969 net6.n1604 net6.n1603 0.005
R3970 net6.n1513 net6.n1512 0.005
R3971 net6.n1757 net6.n1756 0.005
R3972 net6.n1746 net6.n1745 0.005
R3973 net6.n1715 net6.n1714 0.005
R3974 net6.n1704 net6.n1703 0.005
R3975 net6.n1626 net6.n1625 0.005
R3976 net6.n1615 net6.n1614 0.005
R3977 net6.n1576 net6.n1575 0.005
R3978 net6.n1569 net6.n1568 0.005
R3979 net6.n1486 net6.n1485 0.005
R3980 net6.n1483 net6.n1481 0.005
R3981 net6.n1466 net6.n1465 0.005
R3982 net6.n1457 net6.n1456 0.005
R3983 net6.n1455 net6.n1454 0.005
R3984 net6.n1452 net6.n1451 0.005
R3985 net6.n1451 net6.n1448 0.005
R3986 net6.n1447 net6.n1446 0.005
R3987 net6.n1422 net6.n1421 0.005
R3988 net6.n1266 net6.n1265 0.005
R3989 net6.n1233 net6.n1232 0.005
R3990 net6.n1162 net6.n1161 0.005
R3991 net6.n1189 net6.n1188 0.005
R3992 net6.n1367 net6.n1361 0.005
R3993 net6.n1363 net6.n1362 0.005
R3994 net6.n1357 net6.n1354 0.005
R3995 net6.n1330 net6.n1329 0.005
R3996 net6.n1242 net6.n1241 0.005
R3997 net6.n1151 net6.n1150 0.005
R3998 net6.n1395 net6.n1394 0.005
R3999 net6.n1384 net6.n1383 0.005
R4000 net6.n1353 net6.n1352 0.005
R4001 net6.n1342 net6.n1341 0.005
R4002 net6.n1264 net6.n1263 0.005
R4003 net6.n1253 net6.n1252 0.005
R4004 net6.n1214 net6.n1213 0.005
R4005 net6.n1207 net6.n1206 0.005
R4006 net6.n1124 net6.n1123 0.005
R4007 net6.n1121 net6.n1119 0.005
R4008 net6.n1104 net6.n1103 0.005
R4009 net6.n1095 net6.n1094 0.005
R4010 net6.n1093 net6.n1092 0.005
R4011 net6.n1090 net6.n1089 0.005
R4012 net6.n1089 net6.n1086 0.005
R4013 net6.n1085 net6.n1084 0.005
R4014 net6.n1060 net6.n1059 0.005
R4015 net6.n904 net6.n903 0.005
R4016 net6.n871 net6.n870 0.005
R4017 net6.n800 net6.n799 0.005
R4018 net6.n827 net6.n826 0.005
R4019 net6.n1005 net6.n999 0.005
R4020 net6.n1001 net6.n1000 0.005
R4021 net6.n995 net6.n992 0.005
R4022 net6.n968 net6.n967 0.005
R4023 net6.n880 net6.n879 0.005
R4024 net6.n789 net6.n788 0.005
R4025 net6.n1033 net6.n1032 0.005
R4026 net6.n1022 net6.n1021 0.005
R4027 net6.n991 net6.n990 0.005
R4028 net6.n980 net6.n979 0.005
R4029 net6.n902 net6.n901 0.005
R4030 net6.n891 net6.n890 0.005
R4031 net6.n852 net6.n851 0.005
R4032 net6.n845 net6.n844 0.005
R4033 net6.n762 net6.n761 0.005
R4034 net6.n759 net6.n757 0.005
R4035 net6.n742 net6.n741 0.005
R4036 net6.n733 net6.n732 0.005
R4037 net6.n731 net6.n730 0.005
R4038 net6.n728 net6.n727 0.005
R4039 net6.n727 net6.n724 0.005
R4040 net6.n723 net6.n722 0.005
R4041 net6.n698 net6.n697 0.005
R4042 net6.n542 net6.n541 0.005
R4043 net6.n509 net6.n508 0.005
R4044 net6.n438 net6.n437 0.005
R4045 net6.n465 net6.n464 0.005
R4046 net6.n643 net6.n637 0.005
R4047 net6.n639 net6.n638 0.005
R4048 net6.n633 net6.n630 0.005
R4049 net6.n606 net6.n605 0.005
R4050 net6.n518 net6.n517 0.005
R4051 net6.n427 net6.n426 0.005
R4052 net6.n671 net6.n670 0.005
R4053 net6.n660 net6.n659 0.005
R4054 net6.n629 net6.n628 0.005
R4055 net6.n618 net6.n617 0.005
R4056 net6.n540 net6.n539 0.005
R4057 net6.n529 net6.n528 0.005
R4058 net6.n490 net6.n489 0.005
R4059 net6.n483 net6.n482 0.005
R4060 net6.n400 net6.n399 0.005
R4061 net6.n397 net6.n395 0.005
R4062 net6.n380 net6.n379 0.005
R4063 net6.n371 net6.n370 0.005
R4064 net6.n369 net6.n368 0.005
R4065 net6.n366 net6.n365 0.005
R4066 net6.n365 net6.n362 0.005
R4067 net6.n361 net6.n360 0.005
R4068 net6.n336 net6.n335 0.005
R4069 net6.n180 net6.n179 0.005
R4070 net6.n147 net6.n146 0.005
R4071 net6.n76 net6.n75 0.005
R4072 net6.n103 net6.n102 0.005
R4073 net6.n281 net6.n275 0.005
R4074 net6.n277 net6.n276 0.005
R4075 net6.n271 net6.n268 0.005
R4076 net6.n244 net6.n243 0.005
R4077 net6.n156 net6.n155 0.005
R4078 net6.n65 net6.n64 0.005
R4079 net6.n309 net6.n308 0.005
R4080 net6.n298 net6.n297 0.005
R4081 net6.n267 net6.n266 0.005
R4082 net6.n256 net6.n255 0.005
R4083 net6.n178 net6.n177 0.005
R4084 net6.n167 net6.n166 0.005
R4085 net6.n128 net6.n127 0.005
R4086 net6.n121 net6.n120 0.005
R4087 net6.n22 net6.n21 0.004
R4088 net6.n29 net6.n28 0.004
R4089 net6.n33 net6.n32 0.004
R4090 net6.n43 net6.n42 0.004
R4091 net6.n39 net6.n38 0.004
R4092 net6.n10 net6.n9 0.004
R4093 net6.n6 net6.n5 0.004
R4094 net6.n16 net6.n15 0.004
R4095 net6.n20 net6.n19 0.004
R4096 net6.n22 net6.n20 0.004
R4097 net6.n3665 net6.n3664 0.003
R4098 net6.n3478 net6.n3447 0.003
R4099 net6.n3475 net6.n3473 0.003
R4100 net6.n3459 net6.n3458 0.003
R4101 net6.n3334 net6.n3330 0.003
R4102 net6.n3348 net6.n3346 0.003
R4103 net6.n3354 net6.n3353 0.003
R4104 net6.n3365 net6.n3364 0.003
R4105 net6.n3678 net6.n3570 0.003
R4106 net6.n3545 net6.n3544 0.003
R4107 net6.n3536 net6.n3528 0.003
R4108 net6.n3501 net6.n3500 0.003
R4109 net6.n3491 net6.n3484 0.003
R4110 net6.n3412 net6.n3411 0.003
R4111 net6.n3396 net6.n3389 0.003
R4112 net6.n3304 net6.n3303 0.003
R4113 net6.n3117 net6.n3086 0.003
R4114 net6.n3114 net6.n3112 0.003
R4115 net6.n3098 net6.n3097 0.003
R4116 net6.n2973 net6.n2969 0.003
R4117 net6.n2987 net6.n2985 0.003
R4118 net6.n2993 net6.n2992 0.003
R4119 net6.n3004 net6.n3003 0.003
R4120 net6.n3317 net6.n3209 0.003
R4121 net6.n3184 net6.n3183 0.003
R4122 net6.n3175 net6.n3167 0.003
R4123 net6.n3140 net6.n3139 0.003
R4124 net6.n3130 net6.n3123 0.003
R4125 net6.n3051 net6.n3050 0.003
R4126 net6.n3035 net6.n3028 0.003
R4127 net6.n2943 net6.n2942 0.003
R4128 net6.n2756 net6.n2725 0.003
R4129 net6.n2753 net6.n2751 0.003
R4130 net6.n2737 net6.n2736 0.003
R4131 net6.n2612 net6.n2608 0.003
R4132 net6.n2626 net6.n2624 0.003
R4133 net6.n2632 net6.n2631 0.003
R4134 net6.n2643 net6.n2642 0.003
R4135 net6.n2956 net6.n2848 0.003
R4136 net6.n2823 net6.n2822 0.003
R4137 net6.n2814 net6.n2806 0.003
R4138 net6.n2779 net6.n2778 0.003
R4139 net6.n2769 net6.n2762 0.003
R4140 net6.n2690 net6.n2689 0.003
R4141 net6.n2674 net6.n2667 0.003
R4142 net6.n2582 net6.n2581 0.003
R4143 net6.n2395 net6.n2364 0.003
R4144 net6.n2392 net6.n2390 0.003
R4145 net6.n2376 net6.n2375 0.003
R4146 net6.n2251 net6.n2247 0.003
R4147 net6.n2265 net6.n2263 0.003
R4148 net6.n2271 net6.n2270 0.003
R4149 net6.n2282 net6.n2281 0.003
R4150 net6.n2595 net6.n2487 0.003
R4151 net6.n2462 net6.n2461 0.003
R4152 net6.n2453 net6.n2445 0.003
R4153 net6.n2418 net6.n2417 0.003
R4154 net6.n2408 net6.n2401 0.003
R4155 net6.n2329 net6.n2328 0.003
R4156 net6.n2313 net6.n2306 0.003
R4157 net6.n2221 net6.n2220 0.003
R4158 net6.n2034 net6.n2003 0.003
R4159 net6.n2031 net6.n2029 0.003
R4160 net6.n2015 net6.n2014 0.003
R4161 net6.n1890 net6.n1886 0.003
R4162 net6.n1904 net6.n1902 0.003
R4163 net6.n1910 net6.n1909 0.003
R4164 net6.n1921 net6.n1920 0.003
R4165 net6.n2234 net6.n2126 0.003
R4166 net6.n2101 net6.n2100 0.003
R4167 net6.n2092 net6.n2084 0.003
R4168 net6.n2057 net6.n2056 0.003
R4169 net6.n2047 net6.n2040 0.003
R4170 net6.n1968 net6.n1967 0.003
R4171 net6.n1952 net6.n1945 0.003
R4172 net6.n1859 net6.n1858 0.003
R4173 net6.n1672 net6.n1641 0.003
R4174 net6.n1669 net6.n1667 0.003
R4175 net6.n1653 net6.n1652 0.003
R4176 net6.n1528 net6.n1524 0.003
R4177 net6.n1542 net6.n1540 0.003
R4178 net6.n1548 net6.n1547 0.003
R4179 net6.n1559 net6.n1558 0.003
R4180 net6.n1872 net6.n1764 0.003
R4181 net6.n1739 net6.n1738 0.003
R4182 net6.n1730 net6.n1722 0.003
R4183 net6.n1695 net6.n1694 0.003
R4184 net6.n1685 net6.n1678 0.003
R4185 net6.n1606 net6.n1605 0.003
R4186 net6.n1590 net6.n1583 0.003
R4187 net6.n1497 net6.n1496 0.003
R4188 net6.n1310 net6.n1279 0.003
R4189 net6.n1307 net6.n1305 0.003
R4190 net6.n1291 net6.n1290 0.003
R4191 net6.n1166 net6.n1162 0.003
R4192 net6.n1180 net6.n1178 0.003
R4193 net6.n1186 net6.n1185 0.003
R4194 net6.n1197 net6.n1196 0.003
R4195 net6.n1510 net6.n1402 0.003
R4196 net6.n1377 net6.n1376 0.003
R4197 net6.n1368 net6.n1360 0.003
R4198 net6.n1333 net6.n1332 0.003
R4199 net6.n1323 net6.n1316 0.003
R4200 net6.n1244 net6.n1243 0.003
R4201 net6.n1228 net6.n1221 0.003
R4202 net6.n1135 net6.n1134 0.003
R4203 net6.n948 net6.n917 0.003
R4204 net6.n945 net6.n943 0.003
R4205 net6.n929 net6.n928 0.003
R4206 net6.n804 net6.n800 0.003
R4207 net6.n818 net6.n816 0.003
R4208 net6.n824 net6.n823 0.003
R4209 net6.n835 net6.n834 0.003
R4210 net6.n1148 net6.n1040 0.003
R4211 net6.n1015 net6.n1014 0.003
R4212 net6.n1006 net6.n998 0.003
R4213 net6.n971 net6.n970 0.003
R4214 net6.n961 net6.n954 0.003
R4215 net6.n882 net6.n881 0.003
R4216 net6.n866 net6.n859 0.003
R4217 net6.n773 net6.n772 0.003
R4218 net6.n586 net6.n555 0.003
R4219 net6.n583 net6.n581 0.003
R4220 net6.n567 net6.n566 0.003
R4221 net6.n442 net6.n438 0.003
R4222 net6.n456 net6.n454 0.003
R4223 net6.n462 net6.n461 0.003
R4224 net6.n473 net6.n472 0.003
R4225 net6.n786 net6.n678 0.003
R4226 net6.n653 net6.n652 0.003
R4227 net6.n644 net6.n636 0.003
R4228 net6.n609 net6.n608 0.003
R4229 net6.n599 net6.n592 0.003
R4230 net6.n520 net6.n519 0.003
R4231 net6.n504 net6.n497 0.003
R4232 net6.n411 net6.n410 0.003
R4233 net6.n224 net6.n193 0.003
R4234 net6.n221 net6.n219 0.003
R4235 net6.n205 net6.n204 0.003
R4236 net6.n80 net6.n76 0.003
R4237 net6.n94 net6.n92 0.003
R4238 net6.n100 net6.n99 0.003
R4239 net6.n111 net6.n110 0.003
R4240 net6.n424 net6.n316 0.003
R4241 net6.n291 net6.n290 0.003
R4242 net6.n282 net6.n274 0.003
R4243 net6.n247 net6.n246 0.003
R4244 net6.n237 net6.n230 0.003
R4245 net6.n158 net6.n157 0.003
R4246 net6.n142 net6.n135 0.003
R4247 net6.n59 net6.n13 0.002
R4248 net6.n3646 net6.n3645 0.001
R4249 net6.n3641 net6.n3639 0.001
R4250 net6.n3635 net6.n3634 0.001
R4251 net6.n3630 net6.n3629 0.001
R4252 net6.n3613 net6.n3610 0.001
R4253 net6.n3607 net6.n3606 0.001
R4254 net6.n3602 net6.n3599 0.001
R4255 net6.n3597 net6.n3596 0.001
R4256 net6.n3596 net6.n3593 0.001
R4257 net6.n3592 net6.n3591 0.001
R4258 net6.n3586 net6.n3585 0.001
R4259 net6.n3441 net6.n3437 0.001
R4260 net6.n3342 net6.n3339 0.001
R4261 net6.n3344 net6.n3343 0.001
R4262 net6.n3538 net6.n3537 0.001
R4263 net6.n3540 net6.n3539 0.001
R4264 net6.n3507 net6.n3506 0.001
R4265 net6.n3505 net6.n3504 0.001
R4266 net6.n3499 net6.n3494 0.001
R4267 net6.n3490 net6.n3489 0.001
R4268 net6.n3392 net6.n3391 0.001
R4269 net6.n3386 net6.n3385 0.001
R4270 net6.n3322 net6.n3321 0.001
R4271 net6.n3285 net6.n3284 0.001
R4272 net6.n3280 net6.n3278 0.001
R4273 net6.n3274 net6.n3273 0.001
R4274 net6.n3269 net6.n3268 0.001
R4275 net6.n3252 net6.n3249 0.001
R4276 net6.n3246 net6.n3245 0.001
R4277 net6.n3241 net6.n3238 0.001
R4278 net6.n3236 net6.n3235 0.001
R4279 net6.n3235 net6.n3232 0.001
R4280 net6.n3231 net6.n3230 0.001
R4281 net6.n3225 net6.n3224 0.001
R4282 net6.n3080 net6.n3076 0.001
R4283 net6.n2981 net6.n2978 0.001
R4284 net6.n2983 net6.n2982 0.001
R4285 net6.n3177 net6.n3176 0.001
R4286 net6.n3179 net6.n3178 0.001
R4287 net6.n3146 net6.n3145 0.001
R4288 net6.n3144 net6.n3143 0.001
R4289 net6.n3138 net6.n3133 0.001
R4290 net6.n3129 net6.n3128 0.001
R4291 net6.n3031 net6.n3030 0.001
R4292 net6.n3025 net6.n3024 0.001
R4293 net6.n2961 net6.n2960 0.001
R4294 net6.n2924 net6.n2923 0.001
R4295 net6.n2919 net6.n2917 0.001
R4296 net6.n2913 net6.n2912 0.001
R4297 net6.n2908 net6.n2907 0.001
R4298 net6.n2891 net6.n2888 0.001
R4299 net6.n2885 net6.n2884 0.001
R4300 net6.n2880 net6.n2877 0.001
R4301 net6.n2875 net6.n2874 0.001
R4302 net6.n2874 net6.n2871 0.001
R4303 net6.n2870 net6.n2869 0.001
R4304 net6.n2864 net6.n2863 0.001
R4305 net6.n2719 net6.n2715 0.001
R4306 net6.n2620 net6.n2617 0.001
R4307 net6.n2622 net6.n2621 0.001
R4308 net6.n2816 net6.n2815 0.001
R4309 net6.n2818 net6.n2817 0.001
R4310 net6.n2785 net6.n2784 0.001
R4311 net6.n2783 net6.n2782 0.001
R4312 net6.n2777 net6.n2772 0.001
R4313 net6.n2768 net6.n2767 0.001
R4314 net6.n2670 net6.n2669 0.001
R4315 net6.n2664 net6.n2663 0.001
R4316 net6.n2600 net6.n2599 0.001
R4317 net6.n2563 net6.n2562 0.001
R4318 net6.n2558 net6.n2556 0.001
R4319 net6.n2552 net6.n2551 0.001
R4320 net6.n2547 net6.n2546 0.001
R4321 net6.n2530 net6.n2527 0.001
R4322 net6.n2524 net6.n2523 0.001
R4323 net6.n2519 net6.n2516 0.001
R4324 net6.n2514 net6.n2513 0.001
R4325 net6.n2513 net6.n2510 0.001
R4326 net6.n2509 net6.n2508 0.001
R4327 net6.n2503 net6.n2502 0.001
R4328 net6.n2358 net6.n2354 0.001
R4329 net6.n2259 net6.n2256 0.001
R4330 net6.n2261 net6.n2260 0.001
R4331 net6.n2455 net6.n2454 0.001
R4332 net6.n2457 net6.n2456 0.001
R4333 net6.n2424 net6.n2423 0.001
R4334 net6.n2422 net6.n2421 0.001
R4335 net6.n2416 net6.n2411 0.001
R4336 net6.n2407 net6.n2406 0.001
R4337 net6.n2309 net6.n2308 0.001
R4338 net6.n2303 net6.n2302 0.001
R4339 net6.n2239 net6.n2238 0.001
R4340 net6.n2202 net6.n2201 0.001
R4341 net6.n2197 net6.n2195 0.001
R4342 net6.n2191 net6.n2190 0.001
R4343 net6.n2186 net6.n2185 0.001
R4344 net6.n2169 net6.n2166 0.001
R4345 net6.n2163 net6.n2162 0.001
R4346 net6.n2158 net6.n2155 0.001
R4347 net6.n2153 net6.n2152 0.001
R4348 net6.n2152 net6.n2149 0.001
R4349 net6.n2148 net6.n2147 0.001
R4350 net6.n2142 net6.n2141 0.001
R4351 net6.n1997 net6.n1993 0.001
R4352 net6.n1898 net6.n1895 0.001
R4353 net6.n1900 net6.n1899 0.001
R4354 net6.n2094 net6.n2093 0.001
R4355 net6.n2096 net6.n2095 0.001
R4356 net6.n2063 net6.n2062 0.001
R4357 net6.n2061 net6.n2060 0.001
R4358 net6.n2055 net6.n2050 0.001
R4359 net6.n2046 net6.n2045 0.001
R4360 net6.n1948 net6.n1947 0.001
R4361 net6.n1942 net6.n1941 0.001
R4362 net6.n1878 net6.n1877 0.001
R4363 net6.n1840 net6.n1839 0.001
R4364 net6.n1835 net6.n1833 0.001
R4365 net6.n1829 net6.n1828 0.001
R4366 net6.n1824 net6.n1823 0.001
R4367 net6.n1807 net6.n1804 0.001
R4368 net6.n1801 net6.n1800 0.001
R4369 net6.n1796 net6.n1793 0.001
R4370 net6.n1791 net6.n1790 0.001
R4371 net6.n1790 net6.n1787 0.001
R4372 net6.n1786 net6.n1785 0.001
R4373 net6.n1780 net6.n1779 0.001
R4374 net6.n1635 net6.n1631 0.001
R4375 net6.n1536 net6.n1533 0.001
R4376 net6.n1538 net6.n1537 0.001
R4377 net6.n1732 net6.n1731 0.001
R4378 net6.n1734 net6.n1733 0.001
R4379 net6.n1701 net6.n1700 0.001
R4380 net6.n1699 net6.n1698 0.001
R4381 net6.n1693 net6.n1688 0.001
R4382 net6.n1684 net6.n1683 0.001
R4383 net6.n1586 net6.n1585 0.001
R4384 net6.n1580 net6.n1579 0.001
R4385 net6.n1516 net6.n1515 0.001
R4386 net6.n1478 net6.n1477 0.001
R4387 net6.n1473 net6.n1471 0.001
R4388 net6.n1467 net6.n1466 0.001
R4389 net6.n1462 net6.n1461 0.001
R4390 net6.n1445 net6.n1442 0.001
R4391 net6.n1439 net6.n1438 0.001
R4392 net6.n1434 net6.n1431 0.001
R4393 net6.n1429 net6.n1428 0.001
R4394 net6.n1428 net6.n1425 0.001
R4395 net6.n1424 net6.n1423 0.001
R4396 net6.n1418 net6.n1417 0.001
R4397 net6.n1273 net6.n1269 0.001
R4398 net6.n1174 net6.n1171 0.001
R4399 net6.n1176 net6.n1175 0.001
R4400 net6.n1370 net6.n1369 0.001
R4401 net6.n1372 net6.n1371 0.001
R4402 net6.n1339 net6.n1338 0.001
R4403 net6.n1337 net6.n1336 0.001
R4404 net6.n1331 net6.n1326 0.001
R4405 net6.n1322 net6.n1321 0.001
R4406 net6.n1224 net6.n1223 0.001
R4407 net6.n1218 net6.n1217 0.001
R4408 net6.n1154 net6.n1153 0.001
R4409 net6.n1116 net6.n1115 0.001
R4410 net6.n1111 net6.n1109 0.001
R4411 net6.n1105 net6.n1104 0.001
R4412 net6.n1100 net6.n1099 0.001
R4413 net6.n1083 net6.n1080 0.001
R4414 net6.n1077 net6.n1076 0.001
R4415 net6.n1072 net6.n1069 0.001
R4416 net6.n1067 net6.n1066 0.001
R4417 net6.n1066 net6.n1063 0.001
R4418 net6.n1062 net6.n1061 0.001
R4419 net6.n1056 net6.n1055 0.001
R4420 net6.n911 net6.n907 0.001
R4421 net6.n812 net6.n809 0.001
R4422 net6.n814 net6.n813 0.001
R4423 net6.n1008 net6.n1007 0.001
R4424 net6.n1010 net6.n1009 0.001
R4425 net6.n977 net6.n976 0.001
R4426 net6.n975 net6.n974 0.001
R4427 net6.n969 net6.n964 0.001
R4428 net6.n960 net6.n959 0.001
R4429 net6.n862 net6.n861 0.001
R4430 net6.n856 net6.n855 0.001
R4431 net6.n792 net6.n791 0.001
R4432 net6.n754 net6.n753 0.001
R4433 net6.n749 net6.n747 0.001
R4434 net6.n743 net6.n742 0.001
R4435 net6.n738 net6.n737 0.001
R4436 net6.n721 net6.n718 0.001
R4437 net6.n715 net6.n714 0.001
R4438 net6.n710 net6.n707 0.001
R4439 net6.n705 net6.n704 0.001
R4440 net6.n704 net6.n701 0.001
R4441 net6.n700 net6.n699 0.001
R4442 net6.n694 net6.n693 0.001
R4443 net6.n549 net6.n545 0.001
R4444 net6.n450 net6.n447 0.001
R4445 net6.n452 net6.n451 0.001
R4446 net6.n646 net6.n645 0.001
R4447 net6.n648 net6.n647 0.001
R4448 net6.n615 net6.n614 0.001
R4449 net6.n613 net6.n612 0.001
R4450 net6.n607 net6.n602 0.001
R4451 net6.n598 net6.n597 0.001
R4452 net6.n500 net6.n499 0.001
R4453 net6.n494 net6.n493 0.001
R4454 net6.n430 net6.n429 0.001
R4455 net6.n392 net6.n391 0.001
R4456 net6.n387 net6.n385 0.001
R4457 net6.n381 net6.n380 0.001
R4458 net6.n376 net6.n375 0.001
R4459 net6.n359 net6.n356 0.001
R4460 net6.n353 net6.n352 0.001
R4461 net6.n348 net6.n345 0.001
R4462 net6.n343 net6.n342 0.001
R4463 net6.n342 net6.n339 0.001
R4464 net6.n338 net6.n337 0.001
R4465 net6.n332 net6.n331 0.001
R4466 net6.n187 net6.n183 0.001
R4467 net6.n88 net6.n85 0.001
R4468 net6.n90 net6.n89 0.001
R4469 net6.n284 net6.n283 0.001
R4470 net6.n286 net6.n285 0.001
R4471 net6.n253 net6.n252 0.001
R4472 net6.n251 net6.n250 0.001
R4473 net6.n245 net6.n240 0.001
R4474 net6.n236 net6.n235 0.001
R4475 net6.n138 net6.n137 0.001
R4476 net6.n132 net6.n131 0.001
R4477 net6.n68 net6.n67 0.001
R4478 net6.n62 net6.n61 0.001
R4479 net6.n63 net6.n62 0.001
R4480 net6.n13 net6.n12 0.001
R4481 net6.n60 net6.n59 0.001
R4482 net6.n12 net6.n3 0.001
R4483 net6.n61 net6.n60 0.001
R4484 VDD.n10018 VDD.t21 879.678
R4485 VDD.n10062 VDD.t27 774.86
R4486 VDD.n4634 VDD.n2769 390.923
R4487 VDD.n10572 VDD.t2 389.377
R4488 VDD.n10455 VDD.t43 380.543
R4489 VDD.n10109 VDD.t56 372.549
R4490 VDD.n11456 VDD.t28 368.288
R4491 VDD.n11461 VDD.t58 367.617
R4492 VDD.n4632 VDD.n4631 348.776
R4493 VDD.n10225 VDD.t54 343.942
R4494 VDD.n12228 VDD.t17 338.594
R4495 VDD.n11946 VDD.t34 338.283
R4496 VDD.n2029 VDD.n2026 335.489
R4497 VDD.n2030 VDD.n2022 335.203
R4498 VDD.n27 VDD.t0 304.27
R4499 VDD.n12258 VDD.t19 302.58
R4500 VDD.t54 VDD.t35 296.708
R4501 VDD.t56 VDD.t39 265.441
R4502 VDD.t28 VDD.t24 241.976
R4503 VDD.t24 VDD.t29 241.976
R4504 VDD.t29 VDD.t26 241.976
R4505 VDD.t26 VDD.t8 241.976
R4506 VDD.t8 VDD.t25 241.976
R4507 VDD.t9 VDD.t5 241.976
R4508 VDD.t7 VDD.t9 241.976
R4509 VDD.t10 VDD.t7 241.976
R4510 VDD.t6 VDD.t10 241.976
R4511 VDD.t34 VDD.t6 241.976
R4512 VDD.t58 VDD.t50 241.853
R4513 VDD.t50 VDD.t46 241.853
R4514 VDD.t46 VDD.t37 241.853
R4515 VDD.t37 VDD.t48 241.853
R4516 VDD.t48 VDD.t11 241.853
R4517 VDD.t15 VDD.t52 241.853
R4518 VDD.t41 VDD.t15 241.853
R4519 VDD.t30 VDD.t41 241.853
R4520 VDD.t13 VDD.t30 241.853
R4521 VDD.t32 VDD.t13 241.853
R4522 VDD.t17 VDD.t32 241.853
R4523 VDD.n3 VDD.t1 232.401
R4524 VDD.n12234 VDD.t20 232.401
R4525 VDD.n11861 VDD.t22 212.514
R4526 VDD.n11130 VDD.t23 202.483
R4527 VDD.n9 VDD.n8 188.161
R4528 VDD.n12240 VDD.n12239 188.161
R4529 VDD.n2830 VDD.n2829 175.251
R4530 VDD.n4478 VDD.n4477 175.251
R4531 VDD.n233 VDD.n232 175.251
R4532 VDD.n1931 VDD.n1930 175.251
R4533 VDD.n3126 VDD.n3123 172.727
R4534 VDD.n3364 VDD.n3361 172.727
R4535 VDD.n3601 VDD.n3598 172.727
R4536 VDD.n3839 VDD.n3836 172.727
R4537 VDD.n4076 VDD.n4073 172.727
R4538 VDD.n4314 VDD.n4311 172.727
R4539 VDD.n4629 VDD.n2772 172.727
R4540 VDD.n2175 VDD.n2172 172.727
R4541 VDD.n2406 VDD.n2403 172.727
R4542 VDD.n5010 VDD.n5009 172.727
R4543 VDD.n4779 VDD.n4778 172.727
R4544 VDD.n2022 VDD.n198 140.689
R4545 VDD.n4477 VDD.t4 131.474
R4546 VDD.n2829 VDD.t45 131.474
R4547 VDD.n232 VDD.t44 122.709
R4548 VDD.n1930 VDD.t3 122.709
R4549 VDD.n2783 VDD.n2782 102.972
R4550 VDD.n211 VDD.n210 102.972
R4551 VDD.n2026 VDD.n2025 102.972
R4552 VDD.n2022 VDD.n2021 97.033
R4553 VDD.n219 VDD.n218 92.5
R4554 VDD.n333 VDD.n332 92.5
R4555 VDD.n332 VDD.n331 92.5
R4556 VDD.n537 VDD.n536 92.5
R4557 VDD.n536 VDD.n535 92.5
R4558 VDD.n540 VDD.n539 92.5
R4559 VDD.n539 VDD.n538 92.5
R4560 VDD.n771 VDD.n770 92.5
R4561 VDD.n770 VDD.n769 92.5
R4562 VDD.n774 VDD.n773 92.5
R4563 VDD.n773 VDD.n772 92.5
R4564 VDD.n1004 VDD.n1003 92.5
R4565 VDD.n1003 VDD.n1002 92.5
R4566 VDD.n1007 VDD.n1006 92.5
R4567 VDD.n1006 VDD.n1005 92.5
R4568 VDD.n1238 VDD.n1237 92.5
R4569 VDD.n1237 VDD.n1236 92.5
R4570 VDD.n1241 VDD.n1240 92.5
R4571 VDD.n1240 VDD.n1239 92.5
R4572 VDD.n1471 VDD.n1470 92.5
R4573 VDD.n1470 VDD.n1469 92.5
R4574 VDD.n1474 VDD.n1473 92.5
R4575 VDD.n1473 VDD.n1472 92.5
R4576 VDD.n1705 VDD.n1704 92.5
R4577 VDD.n1704 VDD.n1703 92.5
R4578 VDD.n1708 VDD.n1707 92.5
R4579 VDD.n1707 VDD.n1706 92.5
R4580 VDD.n2791 VDD.n2790 92.5
R4581 VDD.n3116 VDD.n3115 92.5
R4582 VDD.n3354 VDD.n3353 92.5
R4583 VDD.n3591 VDD.n3590 92.5
R4584 VDD.n3829 VDD.n3828 92.5
R4585 VDD.n4066 VDD.n4065 92.5
R4586 VDD.n4304 VDD.n4303 92.5
R4587 VDD.n2774 VDD.n2773 92.5
R4588 VDD.n4767 VDD.n4766 92.5
R4589 VDD.n5230 VDD.n5229 92.5
R4590 VDD.n5229 VDD.n5228 92.5
R4591 VDD.n4998 VDD.n4997 92.5
R4592 VDD.n2163 VDD.n2162 92.5
R4593 VDD.n2394 VDD.n2393 92.5
R4594 VDD.n11786 VDD.n11785 92.5
R4595 VDD.n11498 VDD.n11497 92.5
R4596 VDD.n4424 VDD.n4422 89.685
R4597 VDD.n1820 VDD.n1817 86.363
R4598 VDD.n11330 VDD.n11329 61.333
R4599 VDD.n2999 VDD.n2998 56.468
R4600 VDD.n3236 VDD.n3235 56.468
R4601 VDD.n3711 VDD.n3710 56.468
R4602 VDD.n3949 VDD.n3948 56.468
R4603 VDD.n4186 VDD.n4185 56.468
R4604 VDD.n4424 VDD.n4423 56.468
R4605 VDD.n566 VDD.n565 56.468
R4606 VDD.n2805 VDD.n2804 53.146
R4607 VDD.n3109 VDD.n3108 53.146
R4608 VDD.n3126 VDD.n3125 53.146
R4609 VDD.n3153 VDD.n3152 53.146
R4610 VDD.n3347 VDD.n3346 53.146
R4611 VDD.n3364 VDD.n3363 53.146
R4612 VDD.n3584 VDD.n3583 53.146
R4613 VDD.n3601 VDD.n3600 53.146
R4614 VDD.n3822 VDD.n3821 53.146
R4615 VDD.n3839 VDD.n3838 53.146
R4616 VDD.n4059 VDD.n4058 53.146
R4617 VDD.n4076 VDD.n4075 53.146
R4618 VDD.n4267 VDD.n4266 53.146
R4619 VDD.n4297 VDD.n4296 53.146
R4620 VDD.n4314 VDD.n4313 53.146
R4621 VDD.n4620 VDD.n4619 53.146
R4622 VDD.n4630 VDD.n4629 53.146
R4623 VDD.n2154 VDD.n2153 53.146
R4624 VDD.n2175 VDD.n2174 53.146
R4625 VDD.n2385 VDD.n2384 53.146
R4626 VDD.n2406 VDD.n2405 53.146
R4627 VDD.n5219 VDD.n5218 53.146
R4628 VDD.n5285 VDD.n5284 53.146
R4629 VDD.n5010 VDD.n5008 53.146
R4630 VDD.n4989 VDD.n4988 53.146
R4631 VDD.n4779 VDD.n4777 53.146
R4632 VDD.n4758 VDD.n4757 53.146
R4633 VDD.n418 VDD.n417 53.146
R4634 VDD.n430 VDD.n429 53.146
R4635 VDD.n651 VDD.n650 53.146
R4636 VDD.n663 VDD.n662 53.146
R4637 VDD.n897 VDD.n896 53.146
R4638 VDD.n1118 VDD.n1117 53.146
R4639 VDD.n1130 VDD.n1129 53.146
R4640 VDD.n1352 VDD.n1351 53.146
R4641 VDD.n1364 VDD.n1363 53.146
R4642 VDD.n1585 VDD.n1584 53.146
R4643 VDD.n1597 VDD.n1596 53.146
R4644 VDD.n1819 VDD.n1818 53.146
R4645 VDD.n1831 VDD.n1830 53.146
R4646 VDD.n3000 VDD.n2996 51
R4647 VDD.n3237 VDD.n3234 51
R4648 VDD.n3475 VDD.n3471 51
R4649 VDD.n3712 VDD.n3709 51
R4650 VDD.n3950 VDD.n3946 51
R4651 VDD.n4187 VDD.n4184 51
R4652 VDD.n4425 VDD.n4421 51
R4653 VDD.n2986 VDD.n2985 49.825
R4654 VDD.n3010 VDD.n3009 49.825
R4655 VDD.n3224 VDD.n3223 49.825
R4656 VDD.n3247 VDD.n3246 49.825
R4657 VDD.n3461 VDD.n3460 49.825
R4658 VDD.n3485 VDD.n3484 49.825
R4659 VDD.n3699 VDD.n3698 49.825
R4660 VDD.n3722 VDD.n3721 49.825
R4661 VDD.n3936 VDD.n3935 49.825
R4662 VDD.n3960 VDD.n3959 49.825
R4663 VDD.n4174 VDD.n4173 49.825
R4664 VDD.n4197 VDD.n4196 49.825
R4665 VDD.n4411 VDD.n4410 49.825
R4666 VDD.n4435 VDD.n4434 49.825
R4667 VDD.n2041 VDD.n2040 49.825
R4668 VDD.n2055 VDD.n2054 49.825
R4669 VDD.n2272 VDD.n2271 49.825
R4670 VDD.n2286 VDD.n2285 49.825
R4671 VDD.n2511 VDD.n2510 49.825
R4672 VDD.n2581 VDD.n2580 49.825
R4673 VDD.n2736 VDD.n2735 49.825
R4674 VDD.n5114 VDD.n5113 49.825
R4675 VDD.n4890 VDD.n4889 49.825
R4676 VDD.n4876 VDD.n4875 49.825
R4677 VDD.n4659 VDD.n4658 49.825
R4678 VDD.n4645 VDD.n4644 49.825
R4679 VDD.n253 VDD.n252 49.825
R4680 VDD.n529 VDD.n528 49.825
R4681 VDD.n553 VDD.n552 49.825
R4682 VDD.n763 VDD.n762 49.825
R4683 VDD.n787 VDD.n786 49.825
R4684 VDD.n996 VDD.n995 49.825
R4685 VDD.n1020 VDD.n1019 49.825
R4686 VDD.n1230 VDD.n1229 49.825
R4687 VDD.n1254 VDD.n1253 49.825
R4688 VDD.n1463 VDD.n1462 49.825
R4689 VDD.n1487 VDD.n1486 49.825
R4690 VDD.n1667 VDD.n1666 49.825
R4691 VDD.n1697 VDD.n1696 49.825
R4692 VDD.n1721 VDD.n1720 49.825
R4693 VDD.n2015 VDD.n2014 49.825
R4694 VDD.n2785 VDD.n2781 48
R4695 VDD.n2806 VDD.n2802 48
R4696 VDD.n3110 VDD.n3106 48
R4697 VDD.n3127 VDD.n3122 48
R4698 VDD.n3348 VDD.n3344 48
R4699 VDD.n3365 VDD.n3360 48
R4700 VDD.n3585 VDD.n3581 48
R4701 VDD.n3602 VDD.n3597 48
R4702 VDD.n3823 VDD.n3819 48
R4703 VDD.n3840 VDD.n3835 48
R4704 VDD.n4060 VDD.n4056 48
R4705 VDD.n4077 VDD.n4072 48
R4706 VDD.n4298 VDD.n4294 48
R4707 VDD.n4315 VDD.n4310 48
R4708 VDD.n4621 VDD.n4617 48
R4709 VDD.n2837 VDD.n2836 46.503
R4710 VDD.n3095 VDD.n3094 46.503
R4711 VDD.n3140 VDD.n3139 46.503
R4712 VDD.n3333 VDD.n3332 46.503
R4713 VDD.n3378 VDD.n3377 46.503
R4714 VDD.n3570 VDD.n3569 46.503
R4715 VDD.n3615 VDD.n3614 46.503
R4716 VDD.n3808 VDD.n3807 46.503
R4717 VDD.n3853 VDD.n3852 46.503
R4718 VDD.n4045 VDD.n4044 46.503
R4719 VDD.n4090 VDD.n4089 46.503
R4720 VDD.n4283 VDD.n4282 46.503
R4721 VDD.n4328 VDD.n4327 46.503
R4722 VDD.n4557 VDD.n4556 46.503
R4723 VDD.n2140 VDD.n2139 46.503
R4724 VDD.n2189 VDD.n2188 46.503
R4725 VDD.n2371 VDD.n2370 46.503
R4726 VDD.n2420 VDD.n2419 46.503
R4727 VDD.n5199 VDD.n5198 46.503
R4728 VDD.n5266 VDD.n5265 46.503
R4729 VDD.n5024 VDD.n5023 46.503
R4730 VDD.n4975 VDD.n4974 46.503
R4731 VDD.n4793 VDD.n4792 46.503
R4732 VDD.n4744 VDD.n4743 46.503
R4733 VDD.n403 VDD.n402 46.503
R4734 VDD.n444 VDD.n443 46.503
R4735 VDD.n637 VDD.n636 46.503
R4736 VDD.n677 VDD.n676 46.503
R4737 VDD.n870 VDD.n869 46.503
R4738 VDD.n911 VDD.n910 46.503
R4739 VDD.n1104 VDD.n1103 46.503
R4740 VDD.n1144 VDD.n1143 46.503
R4741 VDD.n1337 VDD.n1336 46.503
R4742 VDD.n1378 VDD.n1377 46.503
R4743 VDD.n1571 VDD.n1570 46.503
R4744 VDD.n1611 VDD.n1610 46.503
R4745 VDD.n1804 VDD.n1803 46.503
R4746 VDD.n1845 VDD.n1844 46.503
R4747 VDD.n2984 VDD.n2983 45
R4748 VDD.n3008 VDD.n3007 45
R4749 VDD.n3222 VDD.n3221 45
R4750 VDD.n3245 VDD.n3244 45
R4751 VDD.n3459 VDD.n3458 45
R4752 VDD.n3483 VDD.n3482 45
R4753 VDD.n3697 VDD.n3696 45
R4754 VDD.n3720 VDD.n3719 45
R4755 VDD.n3934 VDD.n3933 45
R4756 VDD.n3958 VDD.n3957 45
R4757 VDD.n4172 VDD.n4171 45
R4758 VDD.n4195 VDD.n4194 45
R4759 VDD.n4409 VDD.n4408 45
R4760 VDD.n4433 VDD.n4432 45
R4761 VDD.n11697 VDD.n11696 44.982
R4762 VDD.n11599 VDD.n11598 44.982
R4763 VDD.n2972 VDD.n2971 43.181
R4764 VDD.n3024 VDD.n3023 43.181
R4765 VDD.n3210 VDD.n3209 43.181
R4766 VDD.n3261 VDD.n3260 43.181
R4767 VDD.n3447 VDD.n3446 43.181
R4768 VDD.n3499 VDD.n3498 43.181
R4769 VDD.n3685 VDD.n3684 43.181
R4770 VDD.n3736 VDD.n3735 43.181
R4771 VDD.n3922 VDD.n3921 43.181
R4772 VDD.n3974 VDD.n3973 43.181
R4773 VDD.n4160 VDD.n4159 43.181
R4774 VDD.n4211 VDD.n4210 43.181
R4775 VDD.n4397 VDD.n4396 43.181
R4776 VDD.n4449 VDD.n4448 43.181
R4777 VDD.n2028 VDD.n2027 43.181
R4778 VDD.n2069 VDD.n2068 43.181
R4779 VDD.n2258 VDD.n2257 43.181
R4780 VDD.n2300 VDD.n2299 43.181
R4781 VDD.n2491 VDD.n2490 43.181
R4782 VDD.n2557 VDD.n2556 43.181
R4783 VDD.n2718 VDD.n2717 43.181
R4784 VDD.n5094 VDD.n5093 43.181
R4785 VDD.n4904 VDD.n4903 43.181
R4786 VDD.n4862 VDD.n4861 43.181
R4787 VDD.n4673 VDD.n4672 43.181
R4788 VDD.n276 VDD.n275 43.181
R4789 VDD.n515 VDD.n514 43.181
R4790 VDD.n568 VDD.n567 43.181
R4791 VDD.n749 VDD.n748 43.181
R4792 VDD.n801 VDD.n800 43.181
R4793 VDD.n982 VDD.n981 43.181
R4794 VDD.n1035 VDD.n1034 43.181
R4795 VDD.n1216 VDD.n1215 43.181
R4796 VDD.n1268 VDD.n1267 43.181
R4797 VDD.n1449 VDD.n1448 43.181
R4798 VDD.n1502 VDD.n1501 43.181
R4799 VDD.n1683 VDD.n1682 43.181
R4800 VDD.n1735 VDD.n1734 43.181
R4801 VDD.n1942 VDD.n1941 43.181
R4802 VDD.n11456 VDD.n11455 42.661
R4803 VDD.n2838 VDD.n2834 42
R4804 VDD.n3096 VDD.n3092 42
R4805 VDD.n3141 VDD.n3137 42
R4806 VDD.n3334 VDD.n3330 42
R4807 VDD.n3379 VDD.n3375 42
R4808 VDD.n3571 VDD.n3567 42
R4809 VDD.n3616 VDD.n3612 42
R4810 VDD.n3809 VDD.n3805 42
R4811 VDD.n3854 VDD.n3850 42
R4812 VDD.n4046 VDD.n4042 42
R4813 VDD.n4091 VDD.n4087 42
R4814 VDD.n4284 VDD.n4280 42
R4815 VDD.n4329 VDD.n4325 42
R4816 VDD.n4558 VDD.n4554 42
R4817 VDD.n2863 VDD.n2862 39.86
R4818 VDD.n3081 VDD.n3080 39.86
R4819 VDD.n3155 VDD.n3154 39.86
R4820 VDD.n3319 VDD.n3317 39.86
R4821 VDD.n3392 VDD.n3391 39.86
R4822 VDD.n3556 VDD.n3555 39.86
R4823 VDD.n3630 VDD.n3629 39.86
R4824 VDD.n3794 VDD.n3793 39.86
R4825 VDD.n3867 VDD.n3866 39.86
R4826 VDD.n4031 VDD.n4030 39.86
R4827 VDD.n4105 VDD.n4104 39.86
R4828 VDD.n4269 VDD.n4268 39.86
R4829 VDD.n4342 VDD.n4341 39.86
R4830 VDD.n4529 VDD.n4528 39.86
R4831 VDD.n2126 VDD.n2125 39.86
R4832 VDD.n2203 VDD.n2202 39.86
R4833 VDD.n2357 VDD.n2356 39.86
R4834 VDD.n2434 VDD.n2433 39.86
R4835 VDD.n5178 VDD.n5177 39.86
R4836 VDD.n5245 VDD.n5244 39.86
R4837 VDD.n5038 VDD.n5037 39.86
R4838 VDD.n4961 VDD.n4960 39.86
R4839 VDD.n4807 VDD.n4806 39.86
R4840 VDD.n4730 VDD.n4729 39.86
R4841 VDD.n389 VDD.n388 39.86
R4842 VDD.n458 VDD.n457 39.86
R4843 VDD.n623 VDD.n622 39.86
R4844 VDD.n691 VDD.n690 39.86
R4845 VDD.n856 VDD.n855 39.86
R4846 VDD.n925 VDD.n924 39.86
R4847 VDD.n1090 VDD.n1089 39.86
R4848 VDD.n1158 VDD.n1157 39.86
R4849 VDD.n1323 VDD.n1322 39.86
R4850 VDD.n1392 VDD.n1391 39.86
R4851 VDD.n1557 VDD.n1556 39.86
R4852 VDD.n1625 VDD.n1624 39.86
R4853 VDD.n1790 VDD.n1789 39.86
R4854 VDD.n1863 VDD.n1862 39.86
R4855 VDD.n2970 VDD.n2969 39
R4856 VDD.n3022 VDD.n3021 39
R4857 VDD.n3208 VDD.n3207 39
R4858 VDD.n3259 VDD.n3258 39
R4859 VDD.n3445 VDD.n3444 39
R4860 VDD.n3497 VDD.n3496 39
R4861 VDD.n3683 VDD.n3682 39
R4862 VDD.n3734 VDD.n3733 39
R4863 VDD.n3920 VDD.n3919 39
R4864 VDD.n3972 VDD.n3971 39
R4865 VDD.n4158 VDD.n4157 39
R4866 VDD.n4209 VDD.n4208 39
R4867 VDD.n4395 VDD.n4394 39
R4868 VDD.n4447 VDD.n4446 39
R4869 VDD.n10688 VDD.n10687 38.453
R4870 VDD.n10567 VDD.n10566 37.672
R4871 VDD.n11945 VDD.n11943 37.055
R4872 VDD.n11945 VDD.n11944 37.055
R4873 VDD.n11126 VDD.n11124 37.055
R4874 VDD.n11129 VDD.n11127 37.055
R4875 VDD.n11126 VDD.n11125 37.055
R4876 VDD.n11129 VDD.n11128 37.055
R4877 VDD.n2958 VDD.n2957 36.538
R4878 VDD.n3038 VDD.n3037 36.538
R4879 VDD.n3196 VDD.n3195 36.538
R4880 VDD.n3275 VDD.n3274 36.538
R4881 VDD.n3433 VDD.n3432 36.538
R4882 VDD.n3513 VDD.n3512 36.538
R4883 VDD.n3671 VDD.n3670 36.538
R4884 VDD.n3750 VDD.n3749 36.538
R4885 VDD.n3908 VDD.n3907 36.538
R4886 VDD.n3988 VDD.n3987 36.538
R4887 VDD.n4146 VDD.n4145 36.538
R4888 VDD.n4225 VDD.n4224 36.538
R4889 VDD.n4383 VDD.n4382 36.538
R4890 VDD.n4468 VDD.n4467 36.538
R4891 VDD.n2083 VDD.n2082 36.538
R4892 VDD.n2244 VDD.n2243 36.538
R4893 VDD.n2314 VDD.n2313 36.538
R4894 VDD.n2475 VDD.n2474 36.538
R4895 VDD.n124 VDD.n123 36.538
R4896 VDD.n2664 VDD.n2663 36.538
R4897 VDD.n5079 VDD.n5078 36.538
R4898 VDD.n4918 VDD.n4917 36.538
R4899 VDD.n4848 VDD.n4847 36.538
R4900 VDD.n4687 VDD.n4686 36.538
R4901 VDD.n307 VDD.n306 36.538
R4902 VDD.n417 VDD.n416 36.538
R4903 VDD.n501 VDD.n500 36.538
R4904 VDD.n582 VDD.n581 36.538
R4905 VDD.n735 VDD.n733 36.538
R4906 VDD.n815 VDD.n814 36.538
R4907 VDD.n968 VDD.n967 36.538
R4908 VDD.n1049 VDD.n1048 36.538
R4909 VDD.n1202 VDD.n1201 36.538
R4910 VDD.n1282 VDD.n1281 36.538
R4911 VDD.n1435 VDD.n1434 36.538
R4912 VDD.n1516 VDD.n1515 36.538
R4913 VDD.n1669 VDD.n1668 36.538
R4914 VDD.n1749 VDD.n1748 36.538
R4915 VDD.n1920 VDD.n1919 36.538
R4916 VDD.n2864 VDD.n2860 36
R4917 VDD.n3082 VDD.n3078 36
R4918 VDD.n3156 VDD.n3151 36
R4919 VDD.n3320 VDD.n3315 36
R4920 VDD.n3393 VDD.n3389 36
R4921 VDD.n3557 VDD.n3553 36
R4922 VDD.n3631 VDD.n3626 36
R4923 VDD.n3795 VDD.n3790 36
R4924 VDD.n3868 VDD.n3864 36
R4925 VDD.n4032 VDD.n4028 36
R4926 VDD.n4106 VDD.n4101 36
R4927 VDD.n4270 VDD.n4265 36
R4928 VDD.n4343 VDD.n4339 36
R4929 VDD.n4530 VDD.n4526 36
R4930 VDD.n10175 VDD.n10174 33.333
R4931 VDD.n10080 VDD.n10079 33.333
R4932 VDD.n10048 VDD.n10047 33.333
R4933 VDD.n2893 VDD.n2892 33.216
R4934 VDD.n2998 VDD.n2997 33.216
R4935 VDD.n3067 VDD.n3066 33.216
R4936 VDD.n3169 VDD.n3168 33.216
R4937 VDD.n3304 VDD.n3303 33.216
R4938 VDD.n3406 VDD.n3405 33.216
R4939 VDD.n3542 VDD.n3541 33.216
R4940 VDD.n3644 VDD.n3643 33.216
R4941 VDD.n3779 VDD.n3778 33.216
R4942 VDD.n3881 VDD.n3880 33.216
R4943 VDD.n4017 VDD.n4016 33.216
R4944 VDD.n4119 VDD.n4118 33.216
R4945 VDD.n4254 VDD.n4253 33.216
R4946 VDD.n4356 VDD.n4355 33.216
R4947 VDD.n4509 VDD.n4508 33.216
R4948 VDD.n2112 VDD.n2111 33.216
R4949 VDD.n2217 VDD.n2216 33.216
R4950 VDD.n2343 VDD.n2342 33.216
R4951 VDD.n2448 VDD.n2447 33.216
R4952 VDD.n5160 VDD.n5159 33.216
R4953 VDD.n2641 VDD.n2640 33.216
R4954 VDD.n5052 VDD.n5051 33.216
R4955 VDD.n4947 VDD.n4946 33.216
R4956 VDD.n4821 VDD.n4820 33.216
R4957 VDD.n4716 VDD.n4715 33.216
R4958 VDD.n375 VDD.n374 33.216
R4959 VDD.n472 VDD.n471 33.216
R4960 VDD.n609 VDD.n608 33.216
R4961 VDD.n705 VDD.n704 33.216
R4962 VDD.n842 VDD.n841 33.216
R4963 VDD.n939 VDD.n938 33.216
R4964 VDD.n1076 VDD.n1075 33.216
R4965 VDD.n1172 VDD.n1171 33.216
R4966 VDD.n1309 VDD.n1308 33.216
R4967 VDD.n1406 VDD.n1405 33.216
R4968 VDD.n1543 VDD.n1542 33.216
R4969 VDD.n1639 VDD.n1638 33.216
R4970 VDD.n1776 VDD.n1775 33.216
R4971 VDD.n1881 VDD.n1880 33.216
R4972 VDD.n415 VDD.n414 33.103
R4973 VDD.n428 VDD.n427 33.103
R4974 VDD.n649 VDD.n648 33.103
R4975 VDD.n661 VDD.n660 33.103
R4976 VDD.n882 VDD.n881 33.103
R4977 VDD.n895 VDD.n894 33.103
R4978 VDD.n1116 VDD.n1115 33.103
R4979 VDD.n1128 VDD.n1127 33.103
R4980 VDD.n1349 VDD.n1348 33.103
R4981 VDD.n1362 VDD.n1361 33.103
R4982 VDD.n1583 VDD.n1582 33.103
R4983 VDD.n1595 VDD.n1594 33.103
R4984 VDD.n1816 VDD.n1815 33.103
R4985 VDD.n1829 VDD.n1828 33.103
R4986 VDD.n2956 VDD.n2955 33
R4987 VDD.n3036 VDD.n3035 33
R4988 VDD.n3194 VDD.n3193 33
R4989 VDD.n3273 VDD.n3272 33
R4990 VDD.n3431 VDD.n3430 33
R4991 VDD.n3511 VDD.n3510 33
R4992 VDD.n3669 VDD.n3668 33
R4993 VDD.n3748 VDD.n3747 33
R4994 VDD.n3906 VDD.n3905 33
R4995 VDD.n3986 VDD.n3985 33
R4996 VDD.n4144 VDD.n4143 33
R4997 VDD.n4223 VDD.n4222 33
R4998 VDD.n4381 VDD.n4380 33
R4999 VDD.n4466 VDD.n4465 33
R5000 VDD.n10293 VDD.n10292 32.727
R5001 VDD.n10640 VDD.n10639 32.727
R5002 VDD.n10521 VDD.n10520 32.727
R5003 VDD.n213 VDD.n209 31.034
R5004 VDD.n254 VDD.n250 31.034
R5005 VDD.n530 VDD.n526 31.034
R5006 VDD.n554 VDD.n550 31.034
R5007 VDD.n764 VDD.n760 31.034
R5008 VDD.n788 VDD.n784 31.034
R5009 VDD.n997 VDD.n993 31.034
R5010 VDD.n1021 VDD.n1017 31.034
R5011 VDD.n1231 VDD.n1227 31.034
R5012 VDD.n1255 VDD.n1251 31.034
R5013 VDD.n1464 VDD.n1460 31.034
R5014 VDD.n1488 VDD.n1484 31.034
R5015 VDD.n1698 VDD.n1694 31.034
R5016 VDD.n1722 VDD.n1718 31.034
R5017 VDD.n2016 VDD.n2012 31.034
R5018 VDD.n2894 VDD.n2890 30
R5019 VDD.n3068 VDD.n3064 30
R5020 VDD.n3170 VDD.n3166 30
R5021 VDD.n3305 VDD.n3301 30
R5022 VDD.n3407 VDD.n3403 30
R5023 VDD.n3543 VDD.n3539 30
R5024 VDD.n3645 VDD.n3641 30
R5025 VDD.n3780 VDD.n3776 30
R5026 VDD.n3882 VDD.n3878 30
R5027 VDD.n4018 VDD.n4014 30
R5028 VDD.n4120 VDD.n4116 30
R5029 VDD.n4255 VDD.n4251 30
R5030 VDD.n4357 VDD.n4353 30
R5031 VDD.n4510 VDD.n4506 30
R5032 VDD.n2911 VDD.n2910 29.895
R5033 VDD.n3052 VDD.n3051 29.895
R5034 VDD.n3182 VDD.n3181 29.895
R5035 VDD.n3289 VDD.n3288 29.895
R5036 VDD.n3419 VDD.n3418 29.895
R5037 VDD.n3474 VDD.n3473 29.895
R5038 VDD.n3527 VDD.n3526 29.895
R5039 VDD.n3657 VDD.n3656 29.895
R5040 VDD.n3764 VDD.n3763 29.895
R5041 VDD.n3894 VDD.n3893 29.895
R5042 VDD.n3949 VDD.n3947 29.895
R5043 VDD.n4002 VDD.n4001 29.895
R5044 VDD.n4132 VDD.n4131 29.895
R5045 VDD.n4239 VDD.n4238 29.895
R5046 VDD.n4369 VDD.n4368 29.895
R5047 VDD.n4488 VDD.n4487 29.895
R5048 VDD.n2097 VDD.n2096 29.895
R5049 VDD.n2230 VDD.n2229 29.895
R5050 VDD.n2328 VDD.n2327 29.895
R5051 VDD.n2461 VDD.n2460 29.895
R5052 VDD.n143 VDD.n142 29.895
R5053 VDD.n2683 VDD.n2682 29.895
R5054 VDD.n5065 VDD.n5064 29.895
R5055 VDD.n4932 VDD.n4931 29.895
R5056 VDD.n4834 VDD.n4833 29.895
R5057 VDD.n4701 VDD.n4700 29.895
R5058 VDD.n325 VDD.n324 29.895
R5059 VDD.n487 VDD.n486 29.895
R5060 VDD.n596 VDD.n595 29.895
R5061 VDD.n720 VDD.n719 29.895
R5062 VDD.n829 VDD.n828 29.895
R5063 VDD.n885 VDD.n884 29.895
R5064 VDD.n954 VDD.n953 29.895
R5065 VDD.n1063 VDD.n1062 29.895
R5066 VDD.n1187 VDD.n1186 29.895
R5067 VDD.n1296 VDD.n1295 29.895
R5068 VDD.n1421 VDD.n1420 29.895
R5069 VDD.n1530 VDD.n1529 29.895
R5070 VDD.n1654 VDD.n1653 29.895
R5071 VDD.n1763 VDD.n1762 29.895
R5072 VDD.n1901 VDD.n1900 29.895
R5073 VDD.n2155 VDD.n2151 29.538
R5074 VDD.n2176 VDD.n2171 29.538
R5075 VDD.n2386 VDD.n2382 29.538
R5076 VDD.n2407 VDD.n2402 29.538
R5077 VDD.n5220 VDD.n5216 29.538
R5078 VDD.n5286 VDD.n5282 29.538
R5079 VDD.n5011 VDD.n5006 29.538
R5080 VDD.n4990 VDD.n4986 29.538
R5081 VDD.n4780 VDD.n4775 29.538
R5082 VDD.n4759 VDD.n4755 29.538
R5083 VDD.n65 VDD.n64 29.09
R5084 VDD.n56 VDD.n55 29.09
R5085 VDD.n11421 VDD.n11420 29.09
R5086 VDD.n11223 VDD.n11222 29.09
R5087 VDD.n11932 VDD.n11931 29.09
R5088 VDD.n12296 VDD.n12295 29.09
R5089 VDD.n12287 VDD.n12286 29.09
R5090 VDD.n401 VDD.n400 28.965
R5091 VDD.n442 VDD.n441 28.965
R5092 VDD.n635 VDD.n634 28.965
R5093 VDD.n675 VDD.n674 28.965
R5094 VDD.n868 VDD.n867 28.965
R5095 VDD.n909 VDD.n908 28.965
R5096 VDD.n1102 VDD.n1101 28.965
R5097 VDD.n1142 VDD.n1141 28.965
R5098 VDD.n1335 VDD.n1334 28.965
R5099 VDD.n1376 VDD.n1375 28.965
R5100 VDD.n1569 VDD.n1568 28.965
R5101 VDD.n1609 VDD.n1608 28.965
R5102 VDD.n1802 VDD.n1801 28.965
R5103 VDD.n1843 VDD.n1842 28.965
R5104 VDD.n10187 VDD.n10186 28.888
R5105 VDD.n10061 VDD.n10060 28.888
R5106 VDD.n10024 VDD.n10023 28.888
R5107 VDD.n11455 VDD.n11454 28.51
R5108 VDD.n10268 VDD.n10267 28.363
R5109 VDD.n10615 VDD.n10614 28.363
R5110 VDD.n10533 VDD.n10532 28.363
R5111 VDD.n64 VDD.n63 27.808
R5112 VDD.n12295 VDD.n12294 27.808
R5113 VDD.n11946 VDD.n11945 27.723
R5114 VDD.n11130 VDD.n11126 27.723
R5115 VDD.n11130 VDD.n11129 27.723
R5116 VDD.n2039 VDD.n2038 27.692
R5117 VDD.n2053 VDD.n2052 27.692
R5118 VDD.n2270 VDD.n2269 27.692
R5119 VDD.n2284 VDD.n2283 27.692
R5120 VDD.n2509 VDD.n2508 27.692
R5121 VDD.n2579 VDD.n2578 27.692
R5122 VDD.n2734 VDD.n2733 27.692
R5123 VDD.n5112 VDD.n5111 27.692
R5124 VDD.n4888 VDD.n4887 27.692
R5125 VDD.n4874 VDD.n4873 27.692
R5126 VDD.n4657 VDD.n4656 27.692
R5127 VDD.n4643 VDD.n4642 27.692
R5128 VDD.n11331 VDD.n11328 27.272
R5129 VDD.n11698 VDD.n11695 27.272
R5130 VDD.n11600 VDD.n11597 27.272
R5131 VDD.n2909 VDD.n2908 27
R5132 VDD.n3050 VDD.n3049 27
R5133 VDD.n3180 VDD.n3179 27
R5134 VDD.n3287 VDD.n3286 27
R5135 VDD.n3417 VDD.n3416 27
R5136 VDD.n3525 VDD.n3524 27
R5137 VDD.n3655 VDD.n3654 27
R5138 VDD.n3762 VDD.n3761 27
R5139 VDD.n3892 VDD.n3891 27
R5140 VDD.n4000 VDD.n3999 27
R5141 VDD.n4130 VDD.n4129 27
R5142 VDD.n4237 VDD.n4236 27
R5143 VDD.n4367 VDD.n4366 27
R5144 VDD.n4486 VDD.n4485 27
R5145 VDD.n277 VDD.n273 26.896
R5146 VDD.n516 VDD.n512 26.896
R5147 VDD.n569 VDD.n564 26.896
R5148 VDD.n750 VDD.n746 26.896
R5149 VDD.n802 VDD.n798 26.896
R5150 VDD.n983 VDD.n979 26.896
R5151 VDD.n1036 VDD.n1031 26.896
R5152 VDD.n1217 VDD.n1213 26.896
R5153 VDD.n1269 VDD.n1265 26.896
R5154 VDD.n1450 VDD.n1446 26.896
R5155 VDD.n1503 VDD.n1498 26.896
R5156 VDD.n1684 VDD.n1680 26.896
R5157 VDD.n1736 VDD.n1732 26.896
R5158 VDD.n1943 VDD.n1939 26.896
R5159 VDD.n2912 VDD.n2911 26.573
R5160 VDD.n3053 VDD.n3052 26.573
R5161 VDD.n3183 VDD.n3182 26.573
R5162 VDD.n3290 VDD.n3289 26.573
R5163 VDD.n3420 VDD.n3419 26.573
R5164 VDD.n3473 VDD.n3472 26.573
R5165 VDD.n3528 VDD.n3527 26.573
R5166 VDD.n3658 VDD.n3657 26.573
R5167 VDD.n3765 VDD.n3764 26.573
R5168 VDD.n3895 VDD.n3894 26.573
R5169 VDD.n4003 VDD.n4002 26.573
R5170 VDD.n4133 VDD.n4132 26.573
R5171 VDD.n4240 VDD.n4239 26.573
R5172 VDD.n4370 VDD.n4369 26.573
R5173 VDD.n4489 VDD.n4488 26.573
R5174 VDD.n2098 VDD.n2097 26.573
R5175 VDD.n2231 VDD.n2230 26.573
R5176 VDD.n2329 VDD.n2328 26.573
R5177 VDD.n2462 VDD.n2461 26.573
R5178 VDD.n144 VDD.n143 26.573
R5179 VDD.n2684 VDD.n2683 26.573
R5180 VDD.n5066 VDD.n5065 26.573
R5181 VDD.n4933 VDD.n4932 26.573
R5182 VDD.n4835 VDD.n4834 26.573
R5183 VDD.n4702 VDD.n4701 26.573
R5184 VDD.n324 VDD.n323 26.573
R5185 VDD.n486 VDD.n485 26.573
R5186 VDD.n595 VDD.n594 26.573
R5187 VDD.n719 VDD.n718 26.573
R5188 VDD.n828 VDD.n827 26.573
R5189 VDD.n953 VDD.n952 26.573
R5190 VDD.n1062 VDD.n1061 26.573
R5191 VDD.n1186 VDD.n1185 26.573
R5192 VDD.n1295 VDD.n1294 26.573
R5193 VDD.n1353 VDD.n1350 26.573
R5194 VDD.n1420 VDD.n1419 26.573
R5195 VDD.n1529 VDD.n1528 26.573
R5196 VDD.n1653 VDD.n1652 26.573
R5197 VDD.n1762 VDD.n1761 26.573
R5198 VDD.n1900 VDD.n1899 26.573
R5199 VDD.n2141 VDD.n2137 25.846
R5200 VDD.n2190 VDD.n2186 25.846
R5201 VDD.n2372 VDD.n2368 25.846
R5202 VDD.n2421 VDD.n2417 25.846
R5203 VDD.n5200 VDD.n5196 25.846
R5204 VDD.n5267 VDD.n5263 25.846
R5205 VDD.n5025 VDD.n5021 25.846
R5206 VDD.n4976 VDD.n4972 25.846
R5207 VDD.n4794 VDD.n4790 25.846
R5208 VDD.n4745 VDD.n4741 25.846
R5209 VDD.n11433 VDD.n11432 25.454
R5210 VDD.n11235 VDD.n11234 25.454
R5211 VDD.n12205 VDD.n12204 25.454
R5212 VDD.n12171 VDD.n12170 25.454
R5213 VDD.n12001 VDD.n12000 25.454
R5214 VDD.n11967 VDD.n11966 25.454
R5215 VDD.n11161 VDD.n11160 25.454
R5216 VDD.n11110 VDD.n11109 25.454
R5217 VDD.n11919 VDD.n11918 25.454
R5218 VDD.n387 VDD.n386 24.827
R5219 VDD.n456 VDD.n455 24.827
R5220 VDD.n621 VDD.n620 24.827
R5221 VDD.n689 VDD.n688 24.827
R5222 VDD.n854 VDD.n853 24.827
R5223 VDD.n923 VDD.n922 24.827
R5224 VDD.n1088 VDD.n1087 24.827
R5225 VDD.n1156 VDD.n1155 24.827
R5226 VDD.n1321 VDD.n1320 24.827
R5227 VDD.n1390 VDD.n1389 24.827
R5228 VDD.n1555 VDD.n1554 24.827
R5229 VDD.n1623 VDD.n1622 24.827
R5230 VDD.n1788 VDD.n1787 24.827
R5231 VDD.n1861 VDD.n1860 24.827
R5232 VDD.n10199 VDD.n10198 24.444
R5233 VDD.n2913 VDD.n2909 24
R5234 VDD.n3054 VDD.n3050 24
R5235 VDD.n3184 VDD.n3180 24
R5236 VDD.n3291 VDD.n3287 24
R5237 VDD.n3421 VDD.n3417 24
R5238 VDD.n3529 VDD.n3525 24
R5239 VDD.n3659 VDD.n3655 24
R5240 VDD.n3766 VDD.n3762 24
R5241 VDD.n3896 VDD.n3892 24
R5242 VDD.n4004 VDD.n4000 24
R5243 VDD.n4134 VDD.n4130 24
R5244 VDD.n4241 VDD.n4237 24
R5245 VDD.n4371 VDD.n4367 24
R5246 VDD.n4490 VDD.n4486 24
R5247 VDD.n2024 VDD.n2023 24
R5248 VDD.n2067 VDD.n2066 24
R5249 VDD.n2256 VDD.n2255 24
R5250 VDD.n2298 VDD.n2297 24
R5251 VDD.n2489 VDD.n2488 24
R5252 VDD.n2555 VDD.n2554 24
R5253 VDD.n2716 VDD.n2715 24
R5254 VDD.n5092 VDD.n5091 24
R5255 VDD.n4902 VDD.n4901 24
R5256 VDD.n4860 VDD.n4859 24
R5257 VDD.n4671 VDD.n4670 24
R5258 VDD.n2771 VDD.n2770 24
R5259 VDD.n10318 VDD.n10317 24
R5260 VDD.n10665 VDD.n10664 24
R5261 VDD.n10545 VDD.n10544 24
R5262 VDD.n11343 VDD.n11342 23.636
R5263 VDD.n12111 VDD.n12109 23.636
R5264 VDD.n12066 VDD.n12064 23.636
R5265 VDD.n10927 VDD.n10925 23.636
R5266 VDD.n11050 VDD.n11048 23.636
R5267 VDD.n10836 VDD.n10834 23.636
R5268 VDD.n10754 VDD.n10752 23.636
R5269 VDD.n11707 VDD.n11706 23.636
R5270 VDD.n11615 VDD.n11614 23.636
R5271 VDD.n2892 VDD.n2891 23.251
R5272 VDD.n3066 VDD.n3065 23.251
R5273 VDD.n3168 VDD.n3167 23.251
R5274 VDD.n3303 VDD.n3302 23.251
R5275 VDD.n3405 VDD.n3404 23.251
R5276 VDD.n3541 VDD.n3540 23.251
R5277 VDD.n3643 VDD.n3642 23.251
R5278 VDD.n3778 VDD.n3777 23.251
R5279 VDD.n3880 VDD.n3879 23.251
R5280 VDD.n4016 VDD.n4015 23.251
R5281 VDD.n4118 VDD.n4117 23.251
R5282 VDD.n4253 VDD.n4252 23.251
R5283 VDD.n4355 VDD.n4354 23.251
R5284 VDD.n4508 VDD.n4507 23.251
R5285 VDD.n2111 VDD.n2110 23.251
R5286 VDD.n2216 VDD.n2215 23.251
R5287 VDD.n2342 VDD.n2341 23.251
R5288 VDD.n2447 VDD.n2446 23.251
R5289 VDD.n5159 VDD.n5158 23.251
R5290 VDD.n2640 VDD.n2639 23.251
R5291 VDD.n5051 VDD.n5050 23.251
R5292 VDD.n4946 VDD.n4945 23.251
R5293 VDD.n4820 VDD.n4819 23.251
R5294 VDD.n4715 VDD.n4714 23.251
R5295 VDD.n376 VDD.n375 23.251
R5296 VDD.n473 VDD.n472 23.251
R5297 VDD.n610 VDD.n609 23.251
R5298 VDD.n706 VDD.n705 23.251
R5299 VDD.n843 VDD.n842 23.251
R5300 VDD.n884 VDD.n883 23.251
R5301 VDD.n940 VDD.n939 23.251
R5302 VDD.n1077 VDD.n1076 23.251
R5303 VDD.n1173 VDD.n1172 23.251
R5304 VDD.n1310 VDD.n1309 23.251
R5305 VDD.n1407 VDD.n1406 23.251
R5306 VDD.n1544 VDD.n1543 23.251
R5307 VDD.n1640 VDD.n1639 23.251
R5308 VDD.n1777 VDD.n1776 23.251
R5309 VDD.n1882 VDD.n1881 23.251
R5310 VDD.n11308 VDD.n11307 22.771
R5311 VDD.n12097 VDD.n12096 22.771
R5312 VDD.n12077 VDD.n12076 22.771
R5313 VDD.n10940 VDD.n10939 22.771
R5314 VDD.n10815 VDD.n10814 22.771
R5315 VDD.n11032 VDD.n11031 22.771
R5316 VDD.n10740 VDD.n10739 22.771
R5317 VDD.n11799 VDD.n11798 22.771
R5318 VDD.n11511 VDD.n11510 22.771
R5319 VDD.n308 VDD.n304 22.758
R5320 VDD.n502 VDD.n498 22.758
R5321 VDD.n583 VDD.n579 22.758
R5322 VDD.n736 VDD.n731 22.758
R5323 VDD.n816 VDD.n812 22.758
R5324 VDD.n969 VDD.n965 22.758
R5325 VDD.n1050 VDD.n1046 22.758
R5326 VDD.n1203 VDD.n1198 22.758
R5327 VDD.n1283 VDD.n1279 22.758
R5328 VDD.n1436 VDD.n1432 22.758
R5329 VDD.n1517 VDD.n1513 22.758
R5330 VDD.n1670 VDD.n1665 22.758
R5331 VDD.n1750 VDD.n1746 22.758
R5332 VDD.n1921 VDD.n1917 22.758
R5333 VDD.n10110 VDD.n10108 22.222
R5334 VDD.n2127 VDD.n2123 22.153
R5335 VDD.n2204 VDD.n2200 22.153
R5336 VDD.n2358 VDD.n2354 22.153
R5337 VDD.n2435 VDD.n2431 22.153
R5338 VDD.n5179 VDD.n5175 22.153
R5339 VDD.n5246 VDD.n5242 22.153
R5340 VDD.n5039 VDD.n5035 22.153
R5341 VDD.n4962 VDD.n4958 22.153
R5342 VDD.n4808 VDD.n4804 22.153
R5343 VDD.n4731 VDD.n4727 22.153
R5344 VDD.n26 VDD.n25 21.818
R5345 VDD.n33 VDD.n32 21.818
R5346 VDD.n10234 VDD.n10233 21.818
R5347 VDD.n10581 VDD.n10580 21.818
R5348 VDD.n10456 VDD.n10454 21.818
R5349 VDD.n11445 VDD.n11444 21.818
R5350 VDD.n11247 VDD.n11246 21.818
R5351 VDD.n11191 VDD.n11190 21.818
R5352 VDD.n11758 VDD.n11757 21.818
R5353 VDD.n12257 VDD.n12256 21.818
R5354 VDD.n12264 VDD.n12263 21.818
R5355 VDD.n2890 VDD.n2889 21
R5356 VDD.n3064 VDD.n3063 21
R5357 VDD.n3166 VDD.n3165 21
R5358 VDD.n3301 VDD.n3300 21
R5359 VDD.n3403 VDD.n3402 21
R5360 VDD.n3539 VDD.n3538 21
R5361 VDD.n3641 VDD.n3640 21
R5362 VDD.n3776 VDD.n3775 21
R5363 VDD.n3878 VDD.n3877 21
R5364 VDD.n4014 VDD.n4013 21
R5365 VDD.n4116 VDD.n4115 21
R5366 VDD.n4251 VDD.n4250 21
R5367 VDD.n4353 VDD.n4352 21
R5368 VDD.n4506 VDD.n4505 21
R5369 VDD.n373 VDD.n372 20.689
R5370 VDD.n470 VDD.n469 20.689
R5371 VDD.n607 VDD.n606 20.689
R5372 VDD.n703 VDD.n702 20.689
R5373 VDD.n840 VDD.n839 20.689
R5374 VDD.n937 VDD.n936 20.689
R5375 VDD.n1074 VDD.n1073 20.689
R5376 VDD.n1170 VDD.n1169 20.689
R5377 VDD.n1307 VDD.n1306 20.689
R5378 VDD.n1404 VDD.n1403 20.689
R5379 VDD.n1541 VDD.n1540 20.689
R5380 VDD.n1637 VDD.n1636 20.689
R5381 VDD.n1774 VDD.n1773 20.689
R5382 VDD.n1879 VDD.n1878 20.689
R5383 VDD.n2081 VDD.n2080 20.307
R5384 VDD.n2242 VDD.n2241 20.307
R5385 VDD.n2312 VDD.n2311 20.307
R5386 VDD.n2473 VDD.n2472 20.307
R5387 VDD.n122 VDD.n121 20.307
R5388 VDD.n2662 VDD.n2661 20.307
R5389 VDD.n5077 VDD.n5076 20.307
R5390 VDD.n4916 VDD.n4915 20.307
R5391 VDD.n4846 VDD.n4845 20.307
R5392 VDD.n4685 VDD.n4684 20.307
R5393 VDD.n11296 VDD.n11295 20.065
R5394 VDD.n11815 VDD.n11814 20.065
R5395 VDD.n11523 VDD.n11522 20.065
R5396 VDD.n10211 VDD.n10210 20
R5397 VDD.n11355 VDD.n11354 20
R5398 VDD.n11684 VDD.n11683 20
R5399 VDD.n11632 VDD.n11631 20
R5400 VDD.n2959 VDD.n2958 19.93
R5401 VDD.n3039 VDD.n3038 19.93
R5402 VDD.n3197 VDD.n3196 19.93
R5403 VDD.n3276 VDD.n3275 19.93
R5404 VDD.n3434 VDD.n3433 19.93
R5405 VDD.n3514 VDD.n3513 19.93
R5406 VDD.n3672 VDD.n3671 19.93
R5407 VDD.n3751 VDD.n3750 19.93
R5408 VDD.n3909 VDD.n3908 19.93
R5409 VDD.n3989 VDD.n3988 19.93
R5410 VDD.n4147 VDD.n4146 19.93
R5411 VDD.n4226 VDD.n4225 19.93
R5412 VDD.n4384 VDD.n4383 19.93
R5413 VDD.n4469 VDD.n4468 19.93
R5414 VDD.n2084 VDD.n2083 19.93
R5415 VDD.n2245 VDD.n2244 19.93
R5416 VDD.n2315 VDD.n2314 19.93
R5417 VDD.n2476 VDD.n2475 19.93
R5418 VDD.n125 VDD.n124 19.93
R5419 VDD.n2665 VDD.n2664 19.93
R5420 VDD.n5080 VDD.n5079 19.93
R5421 VDD.n4919 VDD.n4918 19.93
R5422 VDD.n4849 VDD.n4848 19.93
R5423 VDD.n4688 VDD.n4687 19.93
R5424 VDD.n306 VDD.n305 19.93
R5425 VDD.n500 VDD.n499 19.93
R5426 VDD.n581 VDD.n580 19.93
R5427 VDD.n733 VDD.n732 19.93
R5428 VDD.n814 VDD.n813 19.93
R5429 VDD.n967 VDD.n966 19.93
R5430 VDD.n1048 VDD.n1047 19.93
R5431 VDD.n1281 VDD.n1280 19.93
R5432 VDD.n1434 VDD.n1433 19.93
R5433 VDD.n1515 VDD.n1514 19.93
R5434 VDD.n1668 VDD.n1667 19.93
R5435 VDD.n1748 VDD.n1747 19.93
R5436 VDD.n1919 VDD.n1918 19.93
R5437 VDD.n10243 VDD.n10242 19.636
R5438 VDD.n10590 VDD.n10589 19.636
R5439 VDD.n10557 VDD.n10556 19.636
R5440 VDD.n10116 VDD.n10115 18.987
R5441 VDD.n10226 VDD.n10224 18.677
R5442 VDD.n10573 VDD.n10571 18.677
R5443 VDD.n10462 VDD.n10461 18.677
R5444 VDD.n326 VDD.n322 18.62
R5445 VDD.n488 VDD.n484 18.62
R5446 VDD.n597 VDD.n593 18.62
R5447 VDD.n721 VDD.n717 18.62
R5448 VDD.n830 VDD.n826 18.62
R5449 VDD.n955 VDD.n951 18.62
R5450 VDD.n1064 VDD.n1060 18.62
R5451 VDD.n1188 VDD.n1184 18.62
R5452 VDD.n1297 VDD.n1293 18.62
R5453 VDD.n1422 VDD.n1418 18.62
R5454 VDD.n1531 VDD.n1527 18.62
R5455 VDD.n1655 VDD.n1651 18.62
R5456 VDD.n1764 VDD.n1760 18.62
R5457 VDD.n1902 VDD.n1898 18.62
R5458 VDD.n11648 VDD.n11647 18.51
R5459 VDD.n11475 VDD.n11474 18.51
R5460 VDD.n2113 VDD.n2109 18.461
R5461 VDD.n2218 VDD.n2214 18.461
R5462 VDD.n2344 VDD.n2340 18.461
R5463 VDD.n2449 VDD.n2445 18.461
R5464 VDD.n5161 VDD.n5157 18.461
R5465 VDD.n2642 VDD.n2638 18.461
R5466 VDD.n5053 VDD.n5049 18.461
R5467 VDD.n4948 VDD.n4944 18.461
R5468 VDD.n4822 VDD.n4818 18.461
R5469 VDD.n4717 VDD.n4713 18.461
R5470 VDD.n11259 VDD.n11258 18.181
R5471 VDD.n12146 VDD.n12145 18.181
R5472 VDD.n12026 VDD.n12025 18.181
R5473 VDD.n10886 VDD.n10885 18.181
R5474 VDD.n11003 VDD.n11002 18.181
R5475 VDD.n11092 VDD.n11091 18.181
R5476 VDD.n10712 VDD.n10711 18.181
R5477 VDD.n11771 VDD.n11770 18.181
R5478 VDD.n11482 VDD.n11481 18.181
R5479 VDD.n2960 VDD.n2956 18
R5480 VDD.n3040 VDD.n3036 18
R5481 VDD.n3198 VDD.n3194 18
R5482 VDD.n3277 VDD.n3273 18
R5483 VDD.n3435 VDD.n3431 18
R5484 VDD.n3515 VDD.n3511 18
R5485 VDD.n3673 VDD.n3669 18
R5486 VDD.n3752 VDD.n3748 18
R5487 VDD.n3910 VDD.n3906 18
R5488 VDD.n3990 VDD.n3986 18
R5489 VDD.n4148 VDD.n4144 18
R5490 VDD.n4227 VDD.n4223 18
R5491 VDD.n4385 VDD.n4381 18
R5492 VDD.n4470 VDD.n4466 18
R5493 VDD.n10129 VDD.n10127 17.777
R5494 VDD.n10333 VDD.n10331 17.454
R5495 VDD.n10680 VDD.n10678 17.454
R5496 VDD.n10475 VDD.n10473 17.454
R5497 VDD.n11284 VDD.n11283 17.266
R5498 VDD.n12122 VDD.n12121 17.266
R5499 VDD.n12052 VDD.n12051 17.266
R5500 VDD.n10915 VDD.n10914 17.266
R5501 VDD.n10850 VDD.n10849 17.266
R5502 VDD.n11065 VDD.n11064 17.266
R5503 VDD.n10775 VDD.n10774 17.266
R5504 VDD.n11831 VDD.n11830 17.266
R5505 VDD.n11545 VDD.n11544 17.266
R5506 VDD.n2095 VDD.n2094 16.615
R5507 VDD.n2228 VDD.n2227 16.615
R5508 VDD.n2326 VDD.n2325 16.615
R5509 VDD.n2459 VDD.n2458 16.615
R5510 VDD.n141 VDD.n140 16.615
R5511 VDD.n2681 VDD.n2680 16.615
R5512 VDD.n5063 VDD.n5062 16.615
R5513 VDD.n4930 VDD.n4929 16.615
R5514 VDD.n4832 VDD.n4831 16.615
R5515 VDD.n4699 VDD.n4698 16.615
R5516 VDD.n2862 VDD.n2861 16.608
R5517 VDD.n3080 VDD.n3079 16.608
R5518 VDD.n3154 VDD.n3153 16.608
R5519 VDD.n3317 VDD.n3316 16.608
R5520 VDD.n3391 VDD.n3390 16.608
R5521 VDD.n3555 VDD.n3554 16.608
R5522 VDD.n3866 VDD.n3865 16.608
R5523 VDD.n4030 VDD.n4029 16.608
R5524 VDD.n4104 VDD.n4103 16.608
R5525 VDD.n4268 VDD.n4267 16.608
R5526 VDD.n4341 VDD.n4340 16.608
R5527 VDD.n4528 VDD.n4527 16.608
R5528 VDD.n2125 VDD.n2124 16.608
R5529 VDD.n2202 VDD.n2201 16.608
R5530 VDD.n2356 VDD.n2355 16.608
R5531 VDD.n2433 VDD.n2432 16.608
R5532 VDD.n5177 VDD.n5176 16.608
R5533 VDD.n5244 VDD.n5243 16.608
R5534 VDD.n5037 VDD.n5036 16.608
R5535 VDD.n4960 VDD.n4959 16.608
R5536 VDD.n4806 VDD.n4805 16.608
R5537 VDD.n4729 VDD.n4728 16.608
R5538 VDD.n390 VDD.n389 16.608
R5539 VDD.n459 VDD.n458 16.608
R5540 VDD.n624 VDD.n623 16.608
R5541 VDD.n692 VDD.n691 16.608
R5542 VDD.n857 VDD.n856 16.608
R5543 VDD.n926 VDD.n925 16.608
R5544 VDD.n1091 VDD.n1090 16.608
R5545 VDD.n1159 VDD.n1158 16.608
R5546 VDD.n1324 VDD.n1323 16.608
R5547 VDD.n1393 VDD.n1392 16.608
R5548 VDD.n1558 VDD.n1557 16.608
R5549 VDD.n1626 VDD.n1625 16.608
R5550 VDD.n1791 VDD.n1790 16.608
R5551 VDD.n1864 VDD.n1863 16.608
R5552 VDD.n322 VDD.n321 16.551
R5553 VDD.n484 VDD.n483 16.551
R5554 VDD.n593 VDD.n592 16.551
R5555 VDD.n717 VDD.n716 16.551
R5556 VDD.n826 VDD.n825 16.551
R5557 VDD.n951 VDD.n950 16.551
R5558 VDD.n1060 VDD.n1059 16.551
R5559 VDD.n1184 VDD.n1183 16.551
R5560 VDD.n1293 VDD.n1292 16.551
R5561 VDD.n1418 VDD.n1417 16.551
R5562 VDD.n1527 VDD.n1526 16.551
R5563 VDD.n1651 VDD.n1650 16.551
R5564 VDD.n1760 VDD.n1759 16.551
R5565 VDD.n1898 VDD.n1897 16.551
R5566 VDD.n11367 VDD.n11366 16.363
R5567 VDD.n12136 VDD.n12134 16.363
R5568 VDD.n12041 VDD.n12039 16.363
R5569 VDD.n10904 VDD.n10902 16.363
R5570 VDD.n11082 VDD.n11080 16.363
R5571 VDD.n10869 VDD.n10867 16.363
R5572 VDD.n10696 VDD.n10694 16.363
R5573 VDD.n11672 VDD.n11671 16.363
R5574 VDD.n11586 VDD.n11585 16.363
R5575 VDD.n3 VDD.n2 15.764
R5576 VDD.n12234 VDD.n12233 15.764
R5577 VDD.n10115 VDD.n10114 15.555
R5578 VDD.n10212 VDD.n10211 15.508
R5579 VDD.n10164 VDD.n10163 15.29
R5580 VDD.n10163 VDD.n10162 15.29
R5581 VDD.n10093 VDD.n10092 15.29
R5582 VDD.n10092 VDD.n10091 15.29
R5583 VDD.n10036 VDD.n10035 15.29
R5584 VDD.n10035 VDD.n10034 15.29
R5585 VDD.n10224 VDD.n10223 15.272
R5586 VDD.n10571 VDD.n10570 15.272
R5587 VDD.n10461 VDD.n10460 15.272
R5588 VDD.n10244 VDD.n10243 15.249
R5589 VDD.n10591 VDD.n10590 15.249
R5590 VDD.n10558 VDD.n10557 15.249
R5591 VDD.n10280 VDD.n10279 15.034
R5592 VDD.n10281 VDD.n10280 15.034
R5593 VDD.n10627 VDD.n10626 15.034
R5594 VDD.n10628 VDD.n10627 15.034
R5595 VDD.n10510 VDD.n10509 15.034
R5596 VDD.n10509 VDD.n10508 15.034
R5597 VDD.n2860 VDD.n2859 15
R5598 VDD.n3078 VDD.n3077 15
R5599 VDD.n3151 VDD.n3150 15
R5600 VDD.n3315 VDD.n3314 15
R5601 VDD.n3389 VDD.n3388 15
R5602 VDD.n3553 VDD.n3552 15
R5603 VDD.n3626 VDD.n3625 15
R5604 VDD.n3790 VDD.n3789 15
R5605 VDD.n3864 VDD.n3863 15
R5606 VDD.n4028 VDD.n4027 15
R5607 VDD.n4101 VDD.n4100 15
R5608 VDD.n4265 VDD.n4264 15
R5609 VDD.n4339 VDD.n4338 15
R5610 VDD.n4526 VDD.n4525 15
R5611 VDD.n2099 VDD.n2095 14.769
R5612 VDD.n2232 VDD.n2228 14.769
R5613 VDD.n2330 VDD.n2326 14.769
R5614 VDD.n2463 VDD.n2459 14.769
R5615 VDD.n145 VDD.n141 14.769
R5616 VDD.n2685 VDD.n2681 14.769
R5617 VDD.n5067 VDD.n5063 14.769
R5618 VDD.n4934 VDD.n4930 14.769
R5619 VDD.n4836 VDD.n4832 14.769
R5620 VDD.n4703 VDD.n4699 14.769
R5621 VDD.n11271 VDD.n11270 14.545
R5622 VDD.n11847 VDD.n11846 14.545
R5623 VDD.n11466 VDD.n11465 14.545
R5624 VDD.n377 VDD.n373 14.482
R5625 VDD.n474 VDD.n470 14.482
R5626 VDD.n611 VDD.n607 14.482
R5627 VDD.n707 VDD.n703 14.482
R5628 VDD.n844 VDD.n840 14.482
R5629 VDD.n941 VDD.n937 14.482
R5630 VDD.n1078 VDD.n1074 14.482
R5631 VDD.n1174 VDD.n1170 14.482
R5632 VDD.n1311 VDD.n1307 14.482
R5633 VDD.n1408 VDD.n1404 14.482
R5634 VDD.n1545 VDD.n1541 14.482
R5635 VDD.n1641 VDD.n1637 14.482
R5636 VDD.n1778 VDD.n1774 14.482
R5637 VDD.n1883 VDD.n1879 14.482
R5638 VDD.n11272 VDD.n11271 14.37
R5639 VDD.n11848 VDD.n11847 14.37
R5640 VDD.n11467 VDD.n11466 14.37
R5641 VDD.n11414 VDD.n11413 13.485
R5642 VDD.n11216 VDD.n11215 13.485
R5643 VDD.n12193 VDD.n12192 13.485
R5644 VDD.n12183 VDD.n12182 13.485
R5645 VDD.n11989 VDD.n11988 13.485
R5646 VDD.n11979 VDD.n11978 13.485
R5647 VDD.n12184 VDD.n12183 13.485
R5648 VDD.n11980 VDD.n11979 13.485
R5649 VDD.n11988 VDD.n11987 13.485
R5650 VDD.n12192 VDD.n12191 13.485
R5651 VDD.n11175 VDD.n11174 13.485
R5652 VDD.n11145 VDD.n11144 13.485
R5653 VDD.n11146 VDD.n11145 13.485
R5654 VDD.n11174 VDD.n11173 13.485
R5655 VDD.n11905 VDD.n11904 13.485
R5656 VDD.n11904 VDD.n11903 13.485
R5657 VDD.n11413 VDD.n11412 13.485
R5658 VDD.n11215 VDD.n11214 13.485
R5659 VDD.n10152 VDD.n10151 13.398
R5660 VDD.n10151 VDD.n10150 13.398
R5661 VDD.n10069 VDD.n10068 13.398
R5662 VDD.n10070 VDD.n10069 13.398
R5663 VDD.n10016 VDD.n10015 13.398
R5664 VDD.n10017 VDD.n10016 13.398
R5665 VDD.n10141 VDD.n10140 13.333
R5666 VDD.n2973 VDD.n2972 13.286
R5667 VDD.n3025 VDD.n3024 13.286
R5668 VDD.n3211 VDD.n3210 13.286
R5669 VDD.n3262 VDD.n3261 13.286
R5670 VDD.n3448 VDD.n3447 13.286
R5671 VDD.n3500 VDD.n3499 13.286
R5672 VDD.n3686 VDD.n3685 13.286
R5673 VDD.n3737 VDD.n3736 13.286
R5674 VDD.n3923 VDD.n3922 13.286
R5675 VDD.n3975 VDD.n3974 13.286
R5676 VDD.n4161 VDD.n4160 13.286
R5677 VDD.n4212 VDD.n4211 13.286
R5678 VDD.n4398 VDD.n4397 13.286
R5679 VDD.n4450 VDD.n4449 13.286
R5680 VDD.n2029 VDD.n2028 13.286
R5681 VDD.n2070 VDD.n2069 13.286
R5682 VDD.n2259 VDD.n2258 13.286
R5683 VDD.n2301 VDD.n2300 13.286
R5684 VDD.n2492 VDD.n2491 13.286
R5685 VDD.n2558 VDD.n2557 13.286
R5686 VDD.n2719 VDD.n2718 13.286
R5687 VDD.n5095 VDD.n5094 13.286
R5688 VDD.n4905 VDD.n4904 13.286
R5689 VDD.n4863 VDD.n4862 13.286
R5690 VDD.n4674 VDD.n4673 13.286
R5691 VDD.n275 VDD.n274 13.286
R5692 VDD.n514 VDD.n513 13.286
R5693 VDD.n567 VDD.n566 13.286
R5694 VDD.n735 VDD.n734 13.286
R5695 VDD.n748 VDD.n747 13.286
R5696 VDD.n800 VDD.n799 13.286
R5697 VDD.n981 VDD.n980 13.286
R5698 VDD.n1215 VDD.n1214 13.286
R5699 VDD.n1267 VDD.n1266 13.286
R5700 VDD.n1448 VDD.n1447 13.286
R5701 VDD.n1501 VDD.n1500 13.286
R5702 VDD.n1682 VDD.n1681 13.286
R5703 VDD.n1734 VDD.n1733 13.286
R5704 VDD.n1941 VDD.n1940 13.286
R5705 VDD.n5506 VDD.n5505 13.176
R5706 VDD.n5867 VDD.n5866 13.176
R5707 VDD.n6229 VDD.n6228 13.176
R5708 VDD.n6591 VDD.n6590 13.176
R5709 VDD.n6953 VDD.n6952 13.176
R5710 VDD.n7315 VDD.n7314 13.176
R5711 VDD.n7677 VDD.n7676 13.176
R5712 VDD.n8039 VDD.n8038 13.176
R5713 VDD.n8401 VDD.n8400 13.176
R5714 VDD.n8763 VDD.n8762 13.176
R5715 VDD.n9125 VDD.n9124 13.176
R5716 VDD.n9487 VDD.n9486 13.176
R5717 VDD.n9849 VDD.n9848 13.176
R5718 VDD.n10306 VDD.n10305 13.172
R5719 VDD.n10305 VDD.n10304 13.172
R5720 VDD.n10653 VDD.n10652 13.172
R5721 VDD.n10652 VDD.n10651 13.172
R5722 VDD.n10498 VDD.n10497 13.172
R5723 VDD.n10497 VDD.n10496 13.172
R5724 VDD.n10258 VDD.n10256 13.09
R5725 VDD.n10605 VDD.n10603 13.09
R5726 VDD.n10487 VDD.n10486 13.09
R5727 VDD.n2109 VDD.n2108 12.923
R5728 VDD.n2214 VDD.n2213 12.923
R5729 VDD.n2340 VDD.n2339 12.923
R5730 VDD.n2445 VDD.n2444 12.923
R5731 VDD.n5157 VDD.n5156 12.923
R5732 VDD.n2638 VDD.n2637 12.923
R5733 VDD.n5049 VDD.n5048 12.923
R5734 VDD.n4944 VDD.n4943 12.923
R5735 VDD.n4818 VDD.n4817 12.923
R5736 VDD.n4713 VDD.n4712 12.923
R5737 VDD.n11379 VDD.n11378 12.727
R5738 VDD.n11657 VDD.n11656 12.727
R5739 VDD.n11869 VDD.n11868 12.727
R5740 VDD.n304 VDD.n303 12.413
R5741 VDD.n498 VDD.n497 12.413
R5742 VDD.n579 VDD.n578 12.413
R5743 VDD.n731 VDD.n730 12.413
R5744 VDD.n812 VDD.n811 12.413
R5745 VDD.n965 VDD.n964 12.413
R5746 VDD.n1046 VDD.n1045 12.413
R5747 VDD.n1198 VDD.n1197 12.413
R5748 VDD.n1279 VDD.n1278 12.413
R5749 VDD.n1432 VDD.n1431 12.413
R5750 VDD.n1513 VDD.n1512 12.413
R5751 VDD.n1665 VDD.n1664 12.413
R5752 VDD.n1746 VDD.n1745 12.413
R5753 VDD.n1917 VDD.n1916 12.413
R5754 VDD.n2974 VDD.n2970 12
R5755 VDD.n3026 VDD.n3022 12
R5756 VDD.n3212 VDD.n3208 12
R5757 VDD.n3263 VDD.n3259 12
R5758 VDD.n3449 VDD.n3445 12
R5759 VDD.n3501 VDD.n3497 12
R5760 VDD.n3687 VDD.n3683 12
R5761 VDD.n3738 VDD.n3734 12
R5762 VDD.n3924 VDD.n3920 12
R5763 VDD.n3976 VDD.n3972 12
R5764 VDD.n4162 VDD.n4158 12
R5765 VDD.n4213 VDD.n4209 12
R5766 VDD.n4399 VDD.n4395 12
R5767 VDD.n4451 VDD.n4447 12
R5768 VDD.n78 VDD.n77 11.908
R5769 VDD.n43 VDD.n42 11.908
R5770 VDD.n44 VDD.n43 11.908
R5771 VDD.n77 VDD.n76 11.908
R5772 VDD.n11402 VDD.n11401 11.908
R5773 VDD.n11203 VDD.n11202 11.908
R5774 VDD.n11891 VDD.n11890 11.908
R5775 VDD.n11890 VDD.n11889 11.908
R5776 VDD.n11401 VDD.n11400 11.908
R5777 VDD.n11202 VDD.n11201 11.908
R5778 VDD.n12309 VDD.n12308 11.908
R5779 VDD.n12274 VDD.n12273 11.908
R5780 VDD.n12275 VDD.n12274 11.908
R5781 VDD.n12308 VDD.n12307 11.908
R5782 VDD.n10200 VDD.n10199 11.88
R5783 VDD.n10319 VDD.n10318 11.677
R5784 VDD.n10666 VDD.n10665 11.677
R5785 VDD.n10546 VDD.n10545 11.677
R5786 VDD.n10140 VDD.n10139 11.465
R5787 VDD.n10139 VDD.n10138 11.465
R5788 VDD.n11260 VDD.n11259 11.373
R5789 VDD.n12147 VDD.n12146 11.373
R5790 VDD.n12027 VDD.n12026 11.373
R5791 VDD.n10887 VDD.n10886 11.373
R5792 VDD.n11093 VDD.n11092 11.373
R5793 VDD.n10713 VDD.n10712 11.373
R5794 VDD.n11004 VDD.n11003 11.373
R5795 VDD.n11772 VDD.n11771 11.373
R5796 VDD.n11483 VDD.n11482 11.373
R5797 VDD.n10255 VDD.n10254 11.27
R5798 VDD.n10256 VDD.n10255 11.27
R5799 VDD.n10602 VDD.n10601 11.27
R5800 VDD.n10603 VDD.n10602 11.27
R5801 VDD.n10486 VDD.n10485 11.27
R5802 VDD.n10485 VDD.n10484 11.27
R5803 VDD.n2085 VDD.n2081 11.076
R5804 VDD.n2246 VDD.n2242 11.076
R5805 VDD.n2316 VDD.n2312 11.076
R5806 VDD.n2477 VDD.n2473 11.076
R5807 VDD.n126 VDD.n122 11.076
R5808 VDD.n2666 VDD.n2662 11.076
R5809 VDD.n5081 VDD.n5077 11.076
R5810 VDD.n4920 VDD.n4916 11.076
R5811 VDD.n4850 VDD.n4846 11.076
R5812 VDD.n4689 VDD.n4685 11.076
R5813 VDD.n11283 VDD.n11282 10.909
R5814 VDD.n12121 VDD.n12120 10.909
R5815 VDD.n12051 VDD.n12050 10.909
R5816 VDD.n10914 VDD.n10913 10.909
R5817 VDD.n11064 VDD.n11063 10.909
R5818 VDD.n10849 VDD.n10848 10.909
R5819 VDD.n10774 VDD.n10773 10.909
R5820 VDD.n11830 VDD.n11829 10.909
R5821 VDD.n11544 VDD.n11543 10.909
R5822 VDD.n11959 VDD.n11951 10.868
R5823 VDD.n11194 VDD.n11187 10.867
R5824 VDD.n11647 VDD.n11646 10.37
R5825 VDD.n11474 VDD.n11473 10.37
R5826 VDD.n391 VDD.n387 10.344
R5827 VDD.n460 VDD.n456 10.344
R5828 VDD.n625 VDD.n621 10.344
R5829 VDD.n693 VDD.n689 10.344
R5830 VDD.n858 VDD.n854 10.344
R5831 VDD.n927 VDD.n923 10.344
R5832 VDD.n1092 VDD.n1088 10.344
R5833 VDD.n1160 VDD.n1156 10.344
R5834 VDD.n1325 VDD.n1321 10.344
R5835 VDD.n1394 VDD.n1390 10.344
R5836 VDD.n1559 VDD.n1555 10.344
R5837 VDD.n1627 VDD.n1623 10.344
R5838 VDD.n1792 VDD.n1788 10.344
R5839 VDD.n1865 VDD.n1861 10.344
R5840 VDD.n11390 VDD.n11389 10.302
R5841 VDD.n12218 VDD.n12217 10.302
R5842 VDD.n12158 VDD.n12157 10.302
R5843 VDD.n12014 VDD.n12013 10.302
R5844 VDD.n11955 VDD.n11954 10.302
R5845 VDD.n12159 VDD.n12158 10.302
R5846 VDD.n12013 VDD.n12012 10.302
R5847 VDD.n12217 VDD.n12216 10.302
R5848 VDD.n11956 VDD.n11955 10.302
R5849 VDD.n10877 VDD.n10876 10.302
R5850 VDD.n10989 VDD.n10988 10.302
R5851 VDD.n11122 VDD.n11121 10.302
R5852 VDD.n10704 VDD.n10703 10.302
R5853 VDD.n10703 VDD.n10702 10.302
R5854 VDD.n10878 VDD.n10877 10.302
R5855 VDD.n11123 VDD.n11122 10.302
R5856 VDD.n10988 VDD.n10987 10.302
R5857 VDD.n11860 VDD.n11859 10.302
R5858 VDD.n11859 VDD.n11858 10.302
R5859 VDD.n11389 VDD.n11388 10.302
R5860 VDD.n2836 VDD.n2835 9.965
R5861 VDD.n3094 VDD.n3093 9.965
R5862 VDD.n3139 VDD.n3138 9.965
R5863 VDD.n3319 VDD.n3318 9.965
R5864 VDD.n3332 VDD.n3331 9.965
R5865 VDD.n3377 VDD.n3376 9.965
R5866 VDD.n3569 VDD.n3568 9.965
R5867 VDD.n3614 VDD.n3613 9.965
R5868 VDD.n3629 VDD.n3628 9.965
R5869 VDD.n3793 VDD.n3792 9.965
R5870 VDD.n3807 VDD.n3806 9.965
R5871 VDD.n3852 VDD.n3851 9.965
R5872 VDD.n4044 VDD.n4043 9.965
R5873 VDD.n4089 VDD.n4088 9.965
R5874 VDD.n4105 VDD.n4102 9.965
R5875 VDD.n4282 VDD.n4281 9.965
R5876 VDD.n4327 VDD.n4326 9.965
R5877 VDD.n4556 VDD.n4555 9.965
R5878 VDD.n2139 VDD.n2138 9.965
R5879 VDD.n2188 VDD.n2187 9.965
R5880 VDD.n2370 VDD.n2369 9.965
R5881 VDD.n2419 VDD.n2418 9.965
R5882 VDD.n5198 VDD.n5197 9.965
R5883 VDD.n5265 VDD.n5264 9.965
R5884 VDD.n5023 VDD.n5022 9.965
R5885 VDD.n4974 VDD.n4973 9.965
R5886 VDD.n4792 VDD.n4791 9.965
R5887 VDD.n4743 VDD.n4742 9.965
R5888 VDD.n404 VDD.n403 9.965
R5889 VDD.n445 VDD.n444 9.965
R5890 VDD.n638 VDD.n637 9.965
R5891 VDD.n678 VDD.n677 9.965
R5892 VDD.n871 VDD.n870 9.965
R5893 VDD.n912 VDD.n911 9.965
R5894 VDD.n1034 VDD.n1033 9.965
R5895 VDD.n1105 VDD.n1104 9.965
R5896 VDD.n1145 VDD.n1144 9.965
R5897 VDD.n1200 VDD.n1199 9.965
R5898 VDD.n1201 VDD.n1200 9.965
R5899 VDD.n1338 VDD.n1337 9.965
R5900 VDD.n1379 VDD.n1378 9.965
R5901 VDD.n1572 VDD.n1571 9.965
R5902 VDD.n1612 VDD.n1611 9.965
R5903 VDD.n1805 VDD.n1804 9.965
R5904 VDD.n1846 VDD.n1845 9.965
R5905 VDD.n11460 VDD.n11459 9.72
R5906 VDD.n12227 VDD.n12226 9.72
R5907 VDD.n29 VDD.n28 9.716
R5908 VDD.n35 VDD.n34 9.716
R5909 VDD.n12260 VDD.n12259 9.716
R5910 VDD.n12266 VDD.n12265 9.716
R5911 VDD.n10127 VDD.n10126 9.488
R5912 VDD.n10126 VDD.n10125 9.488
R5913 VDD.n10331 VDD.n10330 9.324
R5914 VDD.n10330 VDD.n10329 9.324
R5915 VDD.n10678 VDD.n10677 9.324
R5916 VDD.n10677 VDD.n10676 9.324
R5917 VDD.n10473 VDD.n10472 9.324
R5918 VDD.n10472 VDD.n10471 9.324
R5919 VDD.n84 VDD.n83 9.3
R5920 VDD.n71 VDD.n70 9.3
R5921 VDD.n52 VDD.n51 9.3
R5922 VDD.n39 VDD.n38 9.3
R5923 VDD.n86 VDD.n85 9.3
R5924 VDD.n82 VDD.n81 9.3
R5925 VDD.n81 VDD.n80 9.3
R5926 VDD.n73 VDD.n72 9.3
R5927 VDD.n69 VDD.n68 9.3
R5928 VDD.n68 VDD.n67 9.3
R5929 VDD.n50 VDD.n49 9.3
R5930 VDD.n60 VDD.n59 9.3
R5931 VDD.n59 VDD.n58 9.3
R5932 VDD.n37 VDD.n36 9.3
R5933 VDD.n48 VDD.n47 9.3
R5934 VDD.n47 VDD.n46 9.3
R5935 VDD.n11 VDD.n10 9.3
R5936 VDD.n5 VDD.n4 9.3
R5937 VDD.n7 VDD.n6 9.3
R5938 VDD.n1933 VDD.n1932 9.3
R5939 VDD.n318 VDD.n316 9.3
R5940 VDD.n4681 VDD.n4680 9.3
R5941 VDD.n4709 VDD.n4708 9.3
R5942 VDD.n4737 VDD.n4736 9.3
R5943 VDD.n4765 VDD.n4764 9.3
R5944 VDD.n4796 VDD.n4795 9.3
R5945 VDD.n4795 VDD.n4794 9.3
R5946 VDD.n4794 VDD.n4793 9.3
R5947 VDD.n4824 VDD.n4823 9.3
R5948 VDD.n4823 VDD.n4822 9.3
R5949 VDD.n4822 VDD.n4821 9.3
R5950 VDD.n4852 VDD.n4851 9.3
R5951 VDD.n4851 VDD.n4850 9.3
R5952 VDD.n4850 VDD.n4849 9.3
R5953 VDD.n4880 VDD.n4879 9.3
R5954 VDD.n4879 VDD.n4878 9.3
R5955 VDD.n4878 VDD.n4877 9.3
R5956 VDD.n4898 VDD.n4897 9.3
R5957 VDD.n4926 VDD.n4925 9.3
R5958 VDD.n4954 VDD.n4953 9.3
R5959 VDD.n4982 VDD.n4981 9.3
R5960 VDD.n5013 VDD.n5012 9.3
R5961 VDD.n5012 VDD.n5011 9.3
R5962 VDD.n5011 VDD.n5010 9.3
R5963 VDD.n5041 VDD.n5040 9.3
R5964 VDD.n5040 VDD.n5039 9.3
R5965 VDD.n5039 VDD.n5038 9.3
R5966 VDD.n5069 VDD.n5068 9.3
R5967 VDD.n5068 VDD.n5067 9.3
R5968 VDD.n5067 VDD.n5066 9.3
R5969 VDD.n5083 VDD.n5082 9.3
R5970 VDD.n5082 VDD.n5081 9.3
R5971 VDD.n5081 VDD.n5080 9.3
R5972 VDD.n5071 VDD.n5070 9.3
R5973 VDD.n5073 VDD.n5072 9.3
R5974 VDD.n5059 VDD.n5058 9.3
R5975 VDD.n5057 VDD.n5056 9.3
R5976 VDD.n5055 VDD.n5054 9.3
R5977 VDD.n5054 VDD.n5053 9.3
R5978 VDD.n5053 VDD.n5052 9.3
R5979 VDD.n5043 VDD.n5042 9.3
R5980 VDD.n5045 VDD.n5044 9.3
R5981 VDD.n5031 VDD.n5030 9.3
R5982 VDD.n5029 VDD.n5028 9.3
R5983 VDD.n5027 VDD.n5026 9.3
R5984 VDD.n5026 VDD.n5025 9.3
R5985 VDD.n5025 VDD.n5024 9.3
R5986 VDD.n5015 VDD.n5014 9.3
R5987 VDD.n5017 VDD.n5016 9.3
R5988 VDD.n5002 VDD.n5001 9.3
R5989 VDD.n5000 VDD.n4999 9.3
R5990 VDD.n4996 VDD.n4995 9.3
R5991 VDD.n4992 VDD.n4991 9.3
R5992 VDD.n4991 VDD.n4990 9.3
R5993 VDD.n4990 VDD.n4989 9.3
R5994 VDD.n4994 VDD.n4993 9.3
R5995 VDD.n4980 VDD.n4979 9.3
R5996 VDD.n4978 VDD.n4977 9.3
R5997 VDD.n4977 VDD.n4976 9.3
R5998 VDD.n4976 VDD.n4975 9.3
R5999 VDD.n4968 VDD.n4967 9.3
R6000 VDD.n4964 VDD.n4963 9.3
R6001 VDD.n4963 VDD.n4962 9.3
R6002 VDD.n4962 VDD.n4961 9.3
R6003 VDD.n4966 VDD.n4965 9.3
R6004 VDD.n4952 VDD.n4951 9.3
R6005 VDD.n4950 VDD.n4949 9.3
R6006 VDD.n4949 VDD.n4948 9.3
R6007 VDD.n4948 VDD.n4947 9.3
R6008 VDD.n4940 VDD.n4939 9.3
R6009 VDD.n4936 VDD.n4935 9.3
R6010 VDD.n4935 VDD.n4934 9.3
R6011 VDD.n4934 VDD.n4933 9.3
R6012 VDD.n4938 VDD.n4937 9.3
R6013 VDD.n4924 VDD.n4923 9.3
R6014 VDD.n4922 VDD.n4921 9.3
R6015 VDD.n4921 VDD.n4920 9.3
R6016 VDD.n4920 VDD.n4919 9.3
R6017 VDD.n4912 VDD.n4911 9.3
R6018 VDD.n4908 VDD.n4907 9.3
R6019 VDD.n4907 VDD.n4906 9.3
R6020 VDD.n4906 VDD.n4905 9.3
R6021 VDD.n4910 VDD.n4909 9.3
R6022 VDD.n4896 VDD.n4895 9.3
R6023 VDD.n4894 VDD.n4893 9.3
R6024 VDD.n4893 VDD.n4892 9.3
R6025 VDD.n4892 VDD.n4891 9.3
R6026 VDD.n4870 VDD.n4869 9.3
R6027 VDD.n4868 VDD.n4867 9.3
R6028 VDD.n4866 VDD.n4865 9.3
R6029 VDD.n4865 VDD.n4864 9.3
R6030 VDD.n4864 VDD.n4863 9.3
R6031 VDD.n4854 VDD.n4853 9.3
R6032 VDD.n4856 VDD.n4855 9.3
R6033 VDD.n4842 VDD.n4841 9.3
R6034 VDD.n4840 VDD.n4839 9.3
R6035 VDD.n4838 VDD.n4837 9.3
R6036 VDD.n4837 VDD.n4836 9.3
R6037 VDD.n4836 VDD.n4835 9.3
R6038 VDD.n4826 VDD.n4825 9.3
R6039 VDD.n4828 VDD.n4827 9.3
R6040 VDD.n4814 VDD.n4813 9.3
R6041 VDD.n4812 VDD.n4811 9.3
R6042 VDD.n4810 VDD.n4809 9.3
R6043 VDD.n4809 VDD.n4808 9.3
R6044 VDD.n4808 VDD.n4807 9.3
R6045 VDD.n4798 VDD.n4797 9.3
R6046 VDD.n4800 VDD.n4799 9.3
R6047 VDD.n4786 VDD.n4785 9.3
R6048 VDD.n4784 VDD.n4783 9.3
R6049 VDD.n4782 VDD.n4781 9.3
R6050 VDD.n4781 VDD.n4780 9.3
R6051 VDD.n4780 VDD.n4779 9.3
R6052 VDD.n4769 VDD.n4768 9.3
R6053 VDD.n4771 VDD.n4770 9.3
R6054 VDD.n4763 VDD.n4762 9.3
R6055 VDD.n4761 VDD.n4760 9.3
R6056 VDD.n4760 VDD.n4759 9.3
R6057 VDD.n4759 VDD.n4758 9.3
R6058 VDD.n4751 VDD.n4750 9.3
R6059 VDD.n4747 VDD.n4746 9.3
R6060 VDD.n4746 VDD.n4745 9.3
R6061 VDD.n4745 VDD.n4744 9.3
R6062 VDD.n4749 VDD.n4748 9.3
R6063 VDD.n4735 VDD.n4734 9.3
R6064 VDD.n4733 VDD.n4732 9.3
R6065 VDD.n4732 VDD.n4731 9.3
R6066 VDD.n4731 VDD.n4730 9.3
R6067 VDD.n4723 VDD.n4722 9.3
R6068 VDD.n4719 VDD.n4718 9.3
R6069 VDD.n4718 VDD.n4717 9.3
R6070 VDD.n4717 VDD.n4716 9.3
R6071 VDD.n4721 VDD.n4720 9.3
R6072 VDD.n4707 VDD.n4706 9.3
R6073 VDD.n4705 VDD.n4704 9.3
R6074 VDD.n4704 VDD.n4703 9.3
R6075 VDD.n4703 VDD.n4702 9.3
R6076 VDD.n4695 VDD.n4694 9.3
R6077 VDD.n4691 VDD.n4690 9.3
R6078 VDD.n4690 VDD.n4689 9.3
R6079 VDD.n4689 VDD.n4688 9.3
R6080 VDD.n4693 VDD.n4692 9.3
R6081 VDD.n4679 VDD.n4678 9.3
R6082 VDD.n4677 VDD.n4676 9.3
R6083 VDD.n4676 VDD.n4675 9.3
R6084 VDD.n4675 VDD.n4674 9.3
R6085 VDD.n4667 VDD.n4666 9.3
R6086 VDD.n4663 VDD.n4662 9.3
R6087 VDD.n4662 VDD.n4661 9.3
R6088 VDD.n4661 VDD.n4660 9.3
R6089 VDD.n4665 VDD.n4664 9.3
R6090 VDD.n4649 VDD.n4648 9.3
R6091 VDD.n4648 VDD.n4647 9.3
R6092 VDD.n4647 VDD.n4646 9.3
R6093 VDD.n4637 VDD.n4636 9.3
R6094 VDD.n4639 VDD.n4638 9.3
R6095 VDD.n4635 VDD.n4634 9.3
R6096 VDD.n2035 VDD.n2034 9.3
R6097 VDD.n2061 VDD.n2060 9.3
R6098 VDD.n2075 VDD.n2074 9.3
R6099 VDD.n2089 VDD.n2088 9.3
R6100 VDD.n2103 VDD.n2102 9.3
R6101 VDD.n2117 VDD.n2116 9.3
R6102 VDD.n2131 VDD.n2130 9.3
R6103 VDD.n2145 VDD.n2144 9.3
R6104 VDD.n2159 VDD.n2158 9.3
R6105 VDD.n2167 VDD.n2166 9.3
R6106 VDD.n2182 VDD.n2181 9.3
R6107 VDD.n2196 VDD.n2195 9.3
R6108 VDD.n2210 VDD.n2209 9.3
R6109 VDD.n2224 VDD.n2223 9.3
R6110 VDD.n2238 VDD.n2237 9.3
R6111 VDD.n2252 VDD.n2251 9.3
R6112 VDD.n2266 VDD.n2265 9.3
R6113 VDD.n2292 VDD.n2291 9.3
R6114 VDD.n2306 VDD.n2305 9.3
R6115 VDD.n2320 VDD.n2319 9.3
R6116 VDD.n2334 VDD.n2333 9.3
R6117 VDD.n2348 VDD.n2347 9.3
R6118 VDD.n2362 VDD.n2361 9.3
R6119 VDD.n2376 VDD.n2375 9.3
R6120 VDD.n2390 VDD.n2389 9.3
R6121 VDD.n2398 VDD.n2397 9.3
R6122 VDD.n2413 VDD.n2412 9.3
R6123 VDD.n2427 VDD.n2426 9.3
R6124 VDD.n2441 VDD.n2440 9.3
R6125 VDD.n2455 VDD.n2454 9.3
R6126 VDD.n2469 VDD.n2468 9.3
R6127 VDD.n2465 VDD.n2464 9.3
R6128 VDD.n2464 VDD.n2463 9.3
R6129 VDD.n2463 VDD.n2462 9.3
R6130 VDD.n2453 VDD.n2452 9.3
R6131 VDD.n2437 VDD.n2436 9.3
R6132 VDD.n2436 VDD.n2435 9.3
R6133 VDD.n2435 VDD.n2434 9.3
R6134 VDD.n2425 VDD.n2424 9.3
R6135 VDD.n2409 VDD.n2408 9.3
R6136 VDD.n2408 VDD.n2407 9.3
R6137 VDD.n2407 VDD.n2406 9.3
R6138 VDD.n2396 VDD.n2395 9.3
R6139 VDD.n2378 VDD.n2377 9.3
R6140 VDD.n2350 VDD.n2349 9.3
R6141 VDD.n2322 VDD.n2321 9.3
R6142 VDD.n2294 VDD.n2293 9.3
R6143 VDD.n2262 VDD.n2261 9.3
R6144 VDD.n2261 VDD.n2260 9.3
R6145 VDD.n2260 VDD.n2259 9.3
R6146 VDD.n2250 VDD.n2249 9.3
R6147 VDD.n2234 VDD.n2233 9.3
R6148 VDD.n2233 VDD.n2232 9.3
R6149 VDD.n2232 VDD.n2231 9.3
R6150 VDD.n2222 VDD.n2221 9.3
R6151 VDD.n2206 VDD.n2205 9.3
R6152 VDD.n2205 VDD.n2204 9.3
R6153 VDD.n2204 VDD.n2203 9.3
R6154 VDD.n2194 VDD.n2193 9.3
R6155 VDD.n2178 VDD.n2177 9.3
R6156 VDD.n2177 VDD.n2176 9.3
R6157 VDD.n2176 VDD.n2175 9.3
R6158 VDD.n2165 VDD.n2164 9.3
R6159 VDD.n2147 VDD.n2146 9.3
R6160 VDD.n2119 VDD.n2118 9.3
R6161 VDD.n2091 VDD.n2090 9.3
R6162 VDD.n2063 VDD.n2062 9.3
R6163 VDD.n2031 VDD.n2030 9.3
R6164 VDD.n2030 VDD.n2029 9.3
R6165 VDD.n2033 VDD.n2032 9.3
R6166 VDD.n2045 VDD.n2044 9.3
R6167 VDD.n2044 VDD.n2043 9.3
R6168 VDD.n2043 VDD.n2042 9.3
R6169 VDD.n2059 VDD.n2058 9.3
R6170 VDD.n2058 VDD.n2057 9.3
R6171 VDD.n2057 VDD.n2056 9.3
R6172 VDD.n2073 VDD.n2072 9.3
R6173 VDD.n2072 VDD.n2071 9.3
R6174 VDD.n2071 VDD.n2070 9.3
R6175 VDD.n2077 VDD.n2076 9.3
R6176 VDD.n2087 VDD.n2086 9.3
R6177 VDD.n2086 VDD.n2085 9.3
R6178 VDD.n2085 VDD.n2084 9.3
R6179 VDD.n2101 VDD.n2100 9.3
R6180 VDD.n2100 VDD.n2099 9.3
R6181 VDD.n2099 VDD.n2098 9.3
R6182 VDD.n2105 VDD.n2104 9.3
R6183 VDD.n2115 VDD.n2114 9.3
R6184 VDD.n2114 VDD.n2113 9.3
R6185 VDD.n2113 VDD.n2112 9.3
R6186 VDD.n2129 VDD.n2128 9.3
R6187 VDD.n2128 VDD.n2127 9.3
R6188 VDD.n2127 VDD.n2126 9.3
R6189 VDD.n2133 VDD.n2132 9.3
R6190 VDD.n2143 VDD.n2142 9.3
R6191 VDD.n2142 VDD.n2141 9.3
R6192 VDD.n2141 VDD.n2140 9.3
R6193 VDD.n2157 VDD.n2156 9.3
R6194 VDD.n2156 VDD.n2155 9.3
R6195 VDD.n2155 VDD.n2154 9.3
R6196 VDD.n2161 VDD.n2160 9.3
R6197 VDD.n2180 VDD.n2179 9.3
R6198 VDD.n2192 VDD.n2191 9.3
R6199 VDD.n2191 VDD.n2190 9.3
R6200 VDD.n2190 VDD.n2189 9.3
R6201 VDD.n2208 VDD.n2207 9.3
R6202 VDD.n2220 VDD.n2219 9.3
R6203 VDD.n2219 VDD.n2218 9.3
R6204 VDD.n2218 VDD.n2217 9.3
R6205 VDD.n2236 VDD.n2235 9.3
R6206 VDD.n2248 VDD.n2247 9.3
R6207 VDD.n2247 VDD.n2246 9.3
R6208 VDD.n2246 VDD.n2245 9.3
R6209 VDD.n2264 VDD.n2263 9.3
R6210 VDD.n2276 VDD.n2275 9.3
R6211 VDD.n2275 VDD.n2274 9.3
R6212 VDD.n2274 VDD.n2273 9.3
R6213 VDD.n2290 VDD.n2289 9.3
R6214 VDD.n2289 VDD.n2288 9.3
R6215 VDD.n2288 VDD.n2287 9.3
R6216 VDD.n2304 VDD.n2303 9.3
R6217 VDD.n2303 VDD.n2302 9.3
R6218 VDD.n2302 VDD.n2301 9.3
R6219 VDD.n2308 VDD.n2307 9.3
R6220 VDD.n2318 VDD.n2317 9.3
R6221 VDD.n2317 VDD.n2316 9.3
R6222 VDD.n2316 VDD.n2315 9.3
R6223 VDD.n2332 VDD.n2331 9.3
R6224 VDD.n2331 VDD.n2330 9.3
R6225 VDD.n2330 VDD.n2329 9.3
R6226 VDD.n2336 VDD.n2335 9.3
R6227 VDD.n2346 VDD.n2345 9.3
R6228 VDD.n2345 VDD.n2344 9.3
R6229 VDD.n2344 VDD.n2343 9.3
R6230 VDD.n2360 VDD.n2359 9.3
R6231 VDD.n2359 VDD.n2358 9.3
R6232 VDD.n2358 VDD.n2357 9.3
R6233 VDD.n2364 VDD.n2363 9.3
R6234 VDD.n2374 VDD.n2373 9.3
R6235 VDD.n2373 VDD.n2372 9.3
R6236 VDD.n2372 VDD.n2371 9.3
R6237 VDD.n2388 VDD.n2387 9.3
R6238 VDD.n2387 VDD.n2386 9.3
R6239 VDD.n2386 VDD.n2385 9.3
R6240 VDD.n2392 VDD.n2391 9.3
R6241 VDD.n2411 VDD.n2410 9.3
R6242 VDD.n2423 VDD.n2422 9.3
R6243 VDD.n2422 VDD.n2421 9.3
R6244 VDD.n2421 VDD.n2420 9.3
R6245 VDD.n2439 VDD.n2438 9.3
R6246 VDD.n2451 VDD.n2450 9.3
R6247 VDD.n2450 VDD.n2449 9.3
R6248 VDD.n2449 VDD.n2448 9.3
R6249 VDD.n2467 VDD.n2466 9.3
R6250 VDD.n2479 VDD.n2478 9.3
R6251 VDD.n2478 VDD.n2477 9.3
R6252 VDD.n2477 VDD.n2476 9.3
R6253 VDD.n5097 VDD.n5096 9.3
R6254 VDD.n5096 VDD.n5095 9.3
R6255 VDD.n2686 VDD.n2685 9.3
R6256 VDD.n2685 VDD.n2684 9.3
R6257 VDD.n2643 VDD.n2642 9.3
R6258 VDD.n2642 VDD.n2641 9.3
R6259 VDD.n5247 VDD.n5246 9.3
R6260 VDD.n5246 VDD.n5245 9.3
R6261 VDD.n5268 VDD.n5267 9.3
R6262 VDD.n5267 VDD.n5266 9.3
R6263 VDD.n5287 VDD.n5286 9.3
R6264 VDD.n5286 VDD.n5285 9.3
R6265 VDD.n5221 VDD.n5220 9.3
R6266 VDD.n5220 VDD.n5219 9.3
R6267 VDD.n5201 VDD.n5200 9.3
R6268 VDD.n5200 VDD.n5199 9.3
R6269 VDD.n5180 VDD.n5179 9.3
R6270 VDD.n5179 VDD.n5178 9.3
R6271 VDD.n5162 VDD.n5161 9.3
R6272 VDD.n5161 VDD.n5160 9.3
R6273 VDD.n146 VDD.n145 9.3
R6274 VDD.n145 VDD.n144 9.3
R6275 VDD.n127 VDD.n126 9.3
R6276 VDD.n126 VDD.n125 9.3
R6277 VDD.n2560 VDD.n2559 9.3
R6278 VDD.n2559 VDD.n2558 9.3
R6279 VDD.n2584 VDD.n2583 9.3
R6280 VDD.n2583 VDD.n2582 9.3
R6281 VDD.n2514 VDD.n2513 9.3
R6282 VDD.n2513 VDD.n2512 9.3
R6283 VDD.n2667 VDD.n2666 9.3
R6284 VDD.n2666 VDD.n2665 9.3
R6285 VDD.n2721 VDD.n2720 9.3
R6286 VDD.n2720 VDD.n2719 9.3
R6287 VDD.n2739 VDD.n2738 9.3
R6288 VDD.n2738 VDD.n2737 9.3
R6289 VDD.n5117 VDD.n5116 9.3
R6290 VDD.n5116 VDD.n5115 9.3
R6291 VDD.n2494 VDD.n2493 9.3
R6292 VDD.n2493 VDD.n2492 9.3
R6293 VDD.n5482 VDD.n5481 9.3
R6294 VDD.n5363 VDD.n5362 9.3
R6295 VDD.n5365 VDD.n5364 9.3
R6296 VDD.n5374 VDD.n5373 9.3
R6297 VDD.n5356 VDD.n5355 9.3
R6298 VDD.n5358 VDD.n5357 9.3
R6299 VDD.n5469 VDD.n5468 9.3
R6300 VDD.n5511 VDD.n5510 9.3
R6301 VDD.n5495 VDD.n5494 9.3
R6302 VDD.n5484 VDD.n5483 9.3
R6303 VDD.n5471 VDD.n5470 9.3
R6304 VDD.n5525 VDD.n5524 9.3
R6305 VDD.n5527 VDD.n5526 9.3
R6306 VDD.n5655 VDD.n5654 9.3
R6307 VDD.n5643 VDD.n5642 9.3
R6308 VDD.n5641 VDD.n5640 9.3
R6309 VDD.n5843 VDD.n5842 9.3
R6310 VDD.n5724 VDD.n5723 9.3
R6311 VDD.n5726 VDD.n5725 9.3
R6312 VDD.n5735 VDD.n5734 9.3
R6313 VDD.n5717 VDD.n5716 9.3
R6314 VDD.n5719 VDD.n5718 9.3
R6315 VDD.n5830 VDD.n5829 9.3
R6316 VDD.n5872 VDD.n5871 9.3
R6317 VDD.n5856 VDD.n5855 9.3
R6318 VDD.n5845 VDD.n5844 9.3
R6319 VDD.n5832 VDD.n5831 9.3
R6320 VDD.n5886 VDD.n5885 9.3
R6321 VDD.n5888 VDD.n5887 9.3
R6322 VDD.n6016 VDD.n6015 9.3
R6323 VDD.n6004 VDD.n6003 9.3
R6324 VDD.n6002 VDD.n6001 9.3
R6325 VDD.n6205 VDD.n6204 9.3
R6326 VDD.n6086 VDD.n6085 9.3
R6327 VDD.n6088 VDD.n6087 9.3
R6328 VDD.n6097 VDD.n6096 9.3
R6329 VDD.n6079 VDD.n6078 9.3
R6330 VDD.n6081 VDD.n6080 9.3
R6331 VDD.n6192 VDD.n6191 9.3
R6332 VDD.n6234 VDD.n6233 9.3
R6333 VDD.n6218 VDD.n6217 9.3
R6334 VDD.n6207 VDD.n6206 9.3
R6335 VDD.n6194 VDD.n6193 9.3
R6336 VDD.n6248 VDD.n6247 9.3
R6337 VDD.n6250 VDD.n6249 9.3
R6338 VDD.n6378 VDD.n6377 9.3
R6339 VDD.n6366 VDD.n6365 9.3
R6340 VDD.n6364 VDD.n6363 9.3
R6341 VDD.n6567 VDD.n6566 9.3
R6342 VDD.n6448 VDD.n6447 9.3
R6343 VDD.n6450 VDD.n6449 9.3
R6344 VDD.n6459 VDD.n6458 9.3
R6345 VDD.n6441 VDD.n6440 9.3
R6346 VDD.n6443 VDD.n6442 9.3
R6347 VDD.n6554 VDD.n6553 9.3
R6348 VDD.n6596 VDD.n6595 9.3
R6349 VDD.n6580 VDD.n6579 9.3
R6350 VDD.n6569 VDD.n6568 9.3
R6351 VDD.n6556 VDD.n6555 9.3
R6352 VDD.n6610 VDD.n6609 9.3
R6353 VDD.n6612 VDD.n6611 9.3
R6354 VDD.n6740 VDD.n6739 9.3
R6355 VDD.n6728 VDD.n6727 9.3
R6356 VDD.n6726 VDD.n6725 9.3
R6357 VDD.n6929 VDD.n6928 9.3
R6358 VDD.n6810 VDD.n6809 9.3
R6359 VDD.n6812 VDD.n6811 9.3
R6360 VDD.n6821 VDD.n6820 9.3
R6361 VDD.n6803 VDD.n6802 9.3
R6362 VDD.n6805 VDD.n6804 9.3
R6363 VDD.n6916 VDD.n6915 9.3
R6364 VDD.n6958 VDD.n6957 9.3
R6365 VDD.n6942 VDD.n6941 9.3
R6366 VDD.n6931 VDD.n6930 9.3
R6367 VDD.n6918 VDD.n6917 9.3
R6368 VDD.n6972 VDD.n6971 9.3
R6369 VDD.n6974 VDD.n6973 9.3
R6370 VDD.n7102 VDD.n7101 9.3
R6371 VDD.n7090 VDD.n7089 9.3
R6372 VDD.n7088 VDD.n7087 9.3
R6373 VDD.n7291 VDD.n7290 9.3
R6374 VDD.n7172 VDD.n7171 9.3
R6375 VDD.n7174 VDD.n7173 9.3
R6376 VDD.n7183 VDD.n7182 9.3
R6377 VDD.n7165 VDD.n7164 9.3
R6378 VDD.n7167 VDD.n7166 9.3
R6379 VDD.n7278 VDD.n7277 9.3
R6380 VDD.n7320 VDD.n7319 9.3
R6381 VDD.n7304 VDD.n7303 9.3
R6382 VDD.n7293 VDD.n7292 9.3
R6383 VDD.n7280 VDD.n7279 9.3
R6384 VDD.n7334 VDD.n7333 9.3
R6385 VDD.n7336 VDD.n7335 9.3
R6386 VDD.n7464 VDD.n7463 9.3
R6387 VDD.n7452 VDD.n7451 9.3
R6388 VDD.n7450 VDD.n7449 9.3
R6389 VDD.n7653 VDD.n7652 9.3
R6390 VDD.n7534 VDD.n7533 9.3
R6391 VDD.n7536 VDD.n7535 9.3
R6392 VDD.n7545 VDD.n7544 9.3
R6393 VDD.n7527 VDD.n7526 9.3
R6394 VDD.n7529 VDD.n7528 9.3
R6395 VDD.n7640 VDD.n7639 9.3
R6396 VDD.n7682 VDD.n7681 9.3
R6397 VDD.n7666 VDD.n7665 9.3
R6398 VDD.n7655 VDD.n7654 9.3
R6399 VDD.n7642 VDD.n7641 9.3
R6400 VDD.n7696 VDD.n7695 9.3
R6401 VDD.n7698 VDD.n7697 9.3
R6402 VDD.n7826 VDD.n7825 9.3
R6403 VDD.n7814 VDD.n7813 9.3
R6404 VDD.n7812 VDD.n7811 9.3
R6405 VDD.n8015 VDD.n8014 9.3
R6406 VDD.n7896 VDD.n7895 9.3
R6407 VDD.n7898 VDD.n7897 9.3
R6408 VDD.n7907 VDD.n7906 9.3
R6409 VDD.n7889 VDD.n7888 9.3
R6410 VDD.n7891 VDD.n7890 9.3
R6411 VDD.n8002 VDD.n8001 9.3
R6412 VDD.n8044 VDD.n8043 9.3
R6413 VDD.n8028 VDD.n8027 9.3
R6414 VDD.n8017 VDD.n8016 9.3
R6415 VDD.n8004 VDD.n8003 9.3
R6416 VDD.n8058 VDD.n8057 9.3
R6417 VDD.n8060 VDD.n8059 9.3
R6418 VDD.n8188 VDD.n8187 9.3
R6419 VDD.n8176 VDD.n8175 9.3
R6420 VDD.n8174 VDD.n8173 9.3
R6421 VDD.n8377 VDD.n8376 9.3
R6422 VDD.n8258 VDD.n8257 9.3
R6423 VDD.n8260 VDD.n8259 9.3
R6424 VDD.n8269 VDD.n8268 9.3
R6425 VDD.n8251 VDD.n8250 9.3
R6426 VDD.n8253 VDD.n8252 9.3
R6427 VDD.n8364 VDD.n8363 9.3
R6428 VDD.n8406 VDD.n8405 9.3
R6429 VDD.n8390 VDD.n8389 9.3
R6430 VDD.n8379 VDD.n8378 9.3
R6431 VDD.n8366 VDD.n8365 9.3
R6432 VDD.n8420 VDD.n8419 9.3
R6433 VDD.n8422 VDD.n8421 9.3
R6434 VDD.n8550 VDD.n8549 9.3
R6435 VDD.n8538 VDD.n8537 9.3
R6436 VDD.n8536 VDD.n8535 9.3
R6437 VDD.n8739 VDD.n8738 9.3
R6438 VDD.n8620 VDD.n8619 9.3
R6439 VDD.n8622 VDD.n8621 9.3
R6440 VDD.n8631 VDD.n8630 9.3
R6441 VDD.n8613 VDD.n8612 9.3
R6442 VDD.n8615 VDD.n8614 9.3
R6443 VDD.n8726 VDD.n8725 9.3
R6444 VDD.n8768 VDD.n8767 9.3
R6445 VDD.n8752 VDD.n8751 9.3
R6446 VDD.n8741 VDD.n8740 9.3
R6447 VDD.n8728 VDD.n8727 9.3
R6448 VDD.n8782 VDD.n8781 9.3
R6449 VDD.n8784 VDD.n8783 9.3
R6450 VDD.n8912 VDD.n8911 9.3
R6451 VDD.n8900 VDD.n8899 9.3
R6452 VDD.n8898 VDD.n8897 9.3
R6453 VDD.n9101 VDD.n9100 9.3
R6454 VDD.n8982 VDD.n8981 9.3
R6455 VDD.n8984 VDD.n8983 9.3
R6456 VDD.n8993 VDD.n8992 9.3
R6457 VDD.n8975 VDD.n8974 9.3
R6458 VDD.n8977 VDD.n8976 9.3
R6459 VDD.n9088 VDD.n9087 9.3
R6460 VDD.n9130 VDD.n9129 9.3
R6461 VDD.n9114 VDD.n9113 9.3
R6462 VDD.n9103 VDD.n9102 9.3
R6463 VDD.n9090 VDD.n9089 9.3
R6464 VDD.n9144 VDD.n9143 9.3
R6465 VDD.n9146 VDD.n9145 9.3
R6466 VDD.n9274 VDD.n9273 9.3
R6467 VDD.n9262 VDD.n9261 9.3
R6468 VDD.n9260 VDD.n9259 9.3
R6469 VDD.n9463 VDD.n9462 9.3
R6470 VDD.n9344 VDD.n9343 9.3
R6471 VDD.n9346 VDD.n9345 9.3
R6472 VDD.n9355 VDD.n9354 9.3
R6473 VDD.n9337 VDD.n9336 9.3
R6474 VDD.n9339 VDD.n9338 9.3
R6475 VDD.n9450 VDD.n9449 9.3
R6476 VDD.n9492 VDD.n9491 9.3
R6477 VDD.n9476 VDD.n9475 9.3
R6478 VDD.n9465 VDD.n9464 9.3
R6479 VDD.n9452 VDD.n9451 9.3
R6480 VDD.n9506 VDD.n9505 9.3
R6481 VDD.n9508 VDD.n9507 9.3
R6482 VDD.n9636 VDD.n9635 9.3
R6483 VDD.n9624 VDD.n9623 9.3
R6484 VDD.n9622 VDD.n9621 9.3
R6485 VDD.n9825 VDD.n9824 9.3
R6486 VDD.n9706 VDD.n9705 9.3
R6487 VDD.n9708 VDD.n9707 9.3
R6488 VDD.n9717 VDD.n9716 9.3
R6489 VDD.n9699 VDD.n9698 9.3
R6490 VDD.n9701 VDD.n9700 9.3
R6491 VDD.n9812 VDD.n9811 9.3
R6492 VDD.n9854 VDD.n9853 9.3
R6493 VDD.n9838 VDD.n9837 9.3
R6494 VDD.n9827 VDD.n9826 9.3
R6495 VDD.n9814 VDD.n9813 9.3
R6496 VDD.n9868 VDD.n9867 9.3
R6497 VDD.n9870 VDD.n9869 9.3
R6498 VDD.n9998 VDD.n9997 9.3
R6499 VDD.n9986 VDD.n9985 9.3
R6500 VDD.n9984 VDD.n9983 9.3
R6501 VDD.n10337 VDD.n10336 9.3
R6502 VDD.n10324 VDD.n10323 9.3
R6503 VDD.n10312 VDD.n10311 9.3
R6504 VDD.n10299 VDD.n10298 9.3
R6505 VDD.n10276 VDD.n10275 9.3
R6506 VDD.n10264 VDD.n10263 9.3
R6507 VDD.n10251 VDD.n10250 9.3
R6508 VDD.n10239 VDD.n10238 9.3
R6509 VDD.n10237 VDD.n10236 9.3
R6510 VDD.n10249 VDD.n10248 9.3
R6511 VDD.n10262 VDD.n10261 9.3
R6512 VDD.n10274 VDD.n10273 9.3
R6513 VDD.n10339 VDD.n10338 9.3
R6514 VDD.n10326 VDD.n10325 9.3
R6515 VDD.n10314 VDD.n10313 9.3
R6516 VDD.n10301 VDD.n10300 9.3
R6517 VDD.n10235 VDD.n10234 9.3
R6518 VDD.n10228 VDD.n10227 9.3
R6519 VDD.n10335 VDD.n10334 9.3
R6520 VDD.n10334 VDD.n10333 9.3
R6521 VDD.n10322 VDD.n10321 9.3
R6522 VDD.n10321 VDD.n10320 9.3
R6523 VDD.n10310 VDD.n10309 9.3
R6524 VDD.n10309 VDD.n10308 9.3
R6525 VDD.n10297 VDD.n10296 9.3
R6526 VDD.n10296 VDD.n10295 9.3
R6527 VDD.n10285 VDD.n10284 9.3
R6528 VDD.n10284 VDD.n10283 9.3
R6529 VDD.n10272 VDD.n10271 9.3
R6530 VDD.n10271 VDD.n10270 9.3
R6531 VDD.n10260 VDD.n10259 9.3
R6532 VDD.n10259 VDD.n10258 9.3
R6533 VDD.n10247 VDD.n10246 9.3
R6534 VDD.n10246 VDD.n10245 9.3
R6535 VDD.n10111 VDD.n10110 9.3
R6536 VDD.n10110 VDD.n10109 9.3
R6537 VDD.n10217 VDD.n10216 9.3
R6538 VDD.n10205 VDD.n10204 9.3
R6539 VDD.n10193 VDD.n10192 9.3
R6540 VDD.n10181 VDD.n10180 9.3
R6541 VDD.n10159 VDD.n10158 9.3
R6542 VDD.n10147 VDD.n10146 9.3
R6543 VDD.n10135 VDD.n10134 9.3
R6544 VDD.n10122 VDD.n10121 9.3
R6545 VDD.n10118 VDD.n10117 9.3
R6546 VDD.n10120 VDD.n10119 9.3
R6547 VDD.n10133 VDD.n10132 9.3
R6548 VDD.n10145 VDD.n10144 9.3
R6549 VDD.n10157 VDD.n10156 9.3
R6550 VDD.n10219 VDD.n10218 9.3
R6551 VDD.n10215 VDD.n10214 9.3
R6552 VDD.n10214 VDD.n10213 9.3
R6553 VDD.n10207 VDD.n10206 9.3
R6554 VDD.n10203 VDD.n10202 9.3
R6555 VDD.n10202 VDD.n10201 9.3
R6556 VDD.n10195 VDD.n10194 9.3
R6557 VDD.n10191 VDD.n10190 9.3
R6558 VDD.n10190 VDD.n10189 9.3
R6559 VDD.n10183 VDD.n10182 9.3
R6560 VDD.n10179 VDD.n10178 9.3
R6561 VDD.n10178 VDD.n10177 9.3
R6562 VDD.n10167 VDD.n10166 9.3
R6563 VDD.n10166 VDD.n10165 9.3
R6564 VDD.n10155 VDD.n10154 9.3
R6565 VDD.n10154 VDD.n10153 9.3
R6566 VDD.n10143 VDD.n10142 9.3
R6567 VDD.n10142 VDD.n10141 9.3
R6568 VDD.n10131 VDD.n10130 9.3
R6569 VDD.n10130 VDD.n10129 9.3
R6570 VDD.n10099 VDD.n10098 9.3
R6571 VDD.n10076 VDD.n10075 9.3
R6572 VDD.n10074 VDD.n10073 9.3
R6573 VDD.n10101 VDD.n10100 9.3
R6574 VDD.n10072 VDD.n10071 9.3
R6575 VDD.n10065 VDD.n10064 9.3
R6576 VDD.n10097 VDD.n10096 9.3
R6577 VDD.n10096 VDD.n10095 9.3
R6578 VDD.n10084 VDD.n10083 9.3
R6579 VDD.n10083 VDD.n10082 9.3
R6580 VDD.n10020 VDD.n10019 9.3
R6581 VDD.n10019 VDD.n10018 9.3
R6582 VDD.n10054 VDD.n10053 9.3
R6583 VDD.n10031 VDD.n10030 9.3
R6584 VDD.n10027 VDD.n10026 9.3
R6585 VDD.n10029 VDD.n10028 9.3
R6586 VDD.n10056 VDD.n10055 9.3
R6587 VDD.n10052 VDD.n10051 9.3
R6588 VDD.n10051 VDD.n10050 9.3
R6589 VDD.n10040 VDD.n10039 9.3
R6590 VDD.n10039 VDD.n10038 9.3
R6591 VDD.n10684 VDD.n10683 9.3
R6592 VDD.n10671 VDD.n10670 9.3
R6593 VDD.n10659 VDD.n10658 9.3
R6594 VDD.n10646 VDD.n10645 9.3
R6595 VDD.n10623 VDD.n10622 9.3
R6596 VDD.n10611 VDD.n10610 9.3
R6597 VDD.n10598 VDD.n10597 9.3
R6598 VDD.n10586 VDD.n10585 9.3
R6599 VDD.n10584 VDD.n10583 9.3
R6600 VDD.n10596 VDD.n10595 9.3
R6601 VDD.n10609 VDD.n10608 9.3
R6602 VDD.n10621 VDD.n10620 9.3
R6603 VDD.n10686 VDD.n10685 9.3
R6604 VDD.n10673 VDD.n10672 9.3
R6605 VDD.n10661 VDD.n10660 9.3
R6606 VDD.n10648 VDD.n10647 9.3
R6607 VDD.n10582 VDD.n10581 9.3
R6608 VDD.n10575 VDD.n10574 9.3
R6609 VDD.n10682 VDD.n10681 9.3
R6610 VDD.n10681 VDD.n10680 9.3
R6611 VDD.n10669 VDD.n10668 9.3
R6612 VDD.n10668 VDD.n10667 9.3
R6613 VDD.n10657 VDD.n10656 9.3
R6614 VDD.n10656 VDD.n10655 9.3
R6615 VDD.n10644 VDD.n10643 9.3
R6616 VDD.n10643 VDD.n10642 9.3
R6617 VDD.n10632 VDD.n10631 9.3
R6618 VDD.n10631 VDD.n10630 9.3
R6619 VDD.n10619 VDD.n10618 9.3
R6620 VDD.n10618 VDD.n10617 9.3
R6621 VDD.n10607 VDD.n10606 9.3
R6622 VDD.n10606 VDD.n10605 9.3
R6623 VDD.n10594 VDD.n10593 9.3
R6624 VDD.n10593 VDD.n10592 9.3
R6625 VDD.n10457 VDD.n10456 9.3
R6626 VDD.n10456 VDD.n10455 9.3
R6627 VDD.n10563 VDD.n10562 9.3
R6628 VDD.n10551 VDD.n10550 9.3
R6629 VDD.n10539 VDD.n10538 9.3
R6630 VDD.n10527 VDD.n10526 9.3
R6631 VDD.n10505 VDD.n10504 9.3
R6632 VDD.n10493 VDD.n10492 9.3
R6633 VDD.n10481 VDD.n10480 9.3
R6634 VDD.n10468 VDD.n10467 9.3
R6635 VDD.n10464 VDD.n10463 9.3
R6636 VDD.n10466 VDD.n10465 9.3
R6637 VDD.n10479 VDD.n10478 9.3
R6638 VDD.n10491 VDD.n10490 9.3
R6639 VDD.n10503 VDD.n10502 9.3
R6640 VDD.n10565 VDD.n10564 9.3
R6641 VDD.n10561 VDD.n10560 9.3
R6642 VDD.n10560 VDD.n10559 9.3
R6643 VDD.n10553 VDD.n10552 9.3
R6644 VDD.n10549 VDD.n10548 9.3
R6645 VDD.n10548 VDD.n10547 9.3
R6646 VDD.n10541 VDD.n10540 9.3
R6647 VDD.n10537 VDD.n10536 9.3
R6648 VDD.n10536 VDD.n10535 9.3
R6649 VDD.n10529 VDD.n10528 9.3
R6650 VDD.n10525 VDD.n10524 9.3
R6651 VDD.n10524 VDD.n10523 9.3
R6652 VDD.n10513 VDD.n10512 9.3
R6653 VDD.n10512 VDD.n10511 9.3
R6654 VDD.n10501 VDD.n10500 9.3
R6655 VDD.n10500 VDD.n10499 9.3
R6656 VDD.n10489 VDD.n10488 9.3
R6657 VDD.n10488 VDD.n10487 9.3
R6658 VDD.n10477 VDD.n10476 9.3
R6659 VDD.n10476 VDD.n10475 9.3
R6660 VDD.n10720 VDD.n10719 9.3
R6661 VDD.n10718 VDD.n10717 9.3
R6662 VDD.n10894 VDD.n10893 9.3
R6663 VDD.n10892 VDD.n10891 9.3
R6664 VDD.n10697 VDD.n10696 9.3
R6665 VDD.n10716 VDD.n10715 9.3
R6666 VDD.n10715 VDD.n10714 9.3
R6667 VDD.n10755 VDD.n10754 9.3
R6668 VDD.n10817 VDD.n10816 9.3
R6669 VDD.n10852 VDD.n10851 9.3
R6670 VDD.n11095 VDD.n11094 9.3
R6671 VDD.n11113 VDD.n11112 9.3
R6672 VDD.n10928 VDD.n10927 9.3
R6673 VDD.n10942 VDD.n10941 9.3
R6674 VDD.n10905 VDD.n10904 9.3
R6675 VDD.n10881 VDD.n10880 9.3
R6676 VDD.n10890 VDD.n10889 9.3
R6677 VDD.n10889 VDD.n10888 9.3
R6678 VDD.n11034 VDD.n11033 9.3
R6679 VDD.n11051 VDD.n11050 9.3
R6680 VDD.n10917 VDD.n10916 9.3
R6681 VDD.n11067 VDD.n11066 9.3
R6682 VDD.n11083 VDD.n11082 9.3
R6683 VDD.n11006 VDD.n11005 9.3
R6684 VDD.n10992 VDD.n10991 9.3
R6685 VDD.n11164 VDD.n11163 9.3
R6686 VDD.n11178 VDD.n11177 9.3
R6687 VDD.n11149 VDD.n11148 9.3
R6688 VDD.n11133 VDD.n11132 9.3
R6689 VDD.n10870 VDD.n10869 9.3
R6690 VDD.n10837 VDD.n10836 9.3
R6691 VDD.n10742 VDD.n10741 9.3
R6692 VDD.n10777 VDD.n10776 9.3
R6693 VDD.n10707 VDD.n10706 9.3
R6694 VDD.n11661 VDD.n11660 9.3
R6695 VDD.n11488 VDD.n11487 9.3
R6696 VDD.n11663 VDD.n11662 9.3
R6697 VDD.n11659 VDD.n11658 9.3
R6698 VDD.n11658 VDD.n11657 9.3
R6699 VDD.n11673 VDD.n11672 9.3
R6700 VDD.n11708 VDD.n11707 9.3
R6701 VDD.n11699 VDD.n11698 9.3
R6702 VDD.n11801 VDD.n11800 9.3
R6703 VDD.n11817 VDD.n11816 9.3
R6704 VDD.n11833 VDD.n11832 9.3
R6705 VDD.n11685 VDD.n11684 9.3
R6706 VDD.n11850 VDD.n11849 9.3
R6707 VDD.n11774 VDD.n11773 9.3
R6708 VDD.n11761 VDD.n11760 9.3
R6709 VDD.n11922 VDD.n11921 9.3
R6710 VDD.n11935 VDD.n11934 9.3
R6711 VDD.n11907 VDD.n11906 9.3
R6712 VDD.n11893 VDD.n11892 9.3
R6713 VDD.n11870 VDD.n11869 9.3
R6714 VDD.n11587 VDD.n11586 9.3
R6715 VDD.n11633 VDD.n11632 9.3
R6716 VDD.n11616 VDD.n11615 9.3
R6717 VDD.n11601 VDD.n11600 9.3
R6718 VDD.n11513 VDD.n11512 9.3
R6719 VDD.n11525 VDD.n11524 9.3
R6720 VDD.n11863 VDD.n11862 9.3
R6721 VDD.n11862 VDD.n11861 9.3
R6722 VDD.n11547 VDD.n11546 9.3
R6723 VDD.n11469 VDD.n11468 9.3
R6724 VDD.n11490 VDD.n11489 9.3
R6725 VDD.n11486 VDD.n11485 9.3
R6726 VDD.n11485 VDD.n11484 9.3
R6727 VDD.n11477 VDD.n11476 9.3
R6728 VDD.n11650 VDD.n11649 9.3
R6729 VDD.n12223 VDD.n12222 9.3
R6730 VDD.n12211 VDD.n12210 9.3
R6731 VDD.n12199 VDD.n12198 9.3
R6732 VDD.n12179 VDD.n12178 9.3
R6733 VDD.n12167 VDD.n12166 9.3
R6734 VDD.n12154 VDD.n12153 9.3
R6735 VDD.n12142 VDD.n12141 9.3
R6736 VDD.n12129 VDD.n12128 9.3
R6737 VDD.n12117 VDD.n12116 9.3
R6738 VDD.n12104 VDD.n12103 9.3
R6739 VDD.n12092 VDD.n12091 9.3
R6740 VDD.n12082 VDD.n12081 9.3
R6741 VDD.n12070 VDD.n12069 9.3
R6742 VDD.n12057 VDD.n12056 9.3
R6743 VDD.n12045 VDD.n12044 9.3
R6744 VDD.n12032 VDD.n12031 9.3
R6745 VDD.n12020 VDD.n12019 9.3
R6746 VDD.n12007 VDD.n12006 9.3
R6747 VDD.n11995 VDD.n11994 9.3
R6748 VDD.n11975 VDD.n11974 9.3
R6749 VDD.n11963 VDD.n11962 9.3
R6750 VDD.n11961 VDD.n11960 9.3
R6751 VDD.n11973 VDD.n11972 9.3
R6752 VDD.n12090 VDD.n12089 9.3
R6753 VDD.n12102 VDD.n12101 9.3
R6754 VDD.n12115 VDD.n12114 9.3
R6755 VDD.n12127 VDD.n12126 9.3
R6756 VDD.n12140 VDD.n12139 9.3
R6757 VDD.n12152 VDD.n12151 9.3
R6758 VDD.n12165 VDD.n12164 9.3
R6759 VDD.n12177 VDD.n12176 9.3
R6760 VDD.n12225 VDD.n12224 9.3
R6761 VDD.n12221 VDD.n12220 9.3
R6762 VDD.n12220 VDD.n12219 9.3
R6763 VDD.n12213 VDD.n12212 9.3
R6764 VDD.n12209 VDD.n12208 9.3
R6765 VDD.n12208 VDD.n12207 9.3
R6766 VDD.n12201 VDD.n12200 9.3
R6767 VDD.n12197 VDD.n12196 9.3
R6768 VDD.n12196 VDD.n12195 9.3
R6769 VDD.n12188 VDD.n12187 9.3
R6770 VDD.n12187 VDD.n12186 9.3
R6771 VDD.n12175 VDD.n12174 9.3
R6772 VDD.n12174 VDD.n12173 9.3
R6773 VDD.n12163 VDD.n12162 9.3
R6774 VDD.n12162 VDD.n12161 9.3
R6775 VDD.n12150 VDD.n12149 9.3
R6776 VDD.n12149 VDD.n12148 9.3
R6777 VDD.n12138 VDD.n12137 9.3
R6778 VDD.n12137 VDD.n12136 9.3
R6779 VDD.n12125 VDD.n12124 9.3
R6780 VDD.n12124 VDD.n12123 9.3
R6781 VDD.n12113 VDD.n12112 9.3
R6782 VDD.n12112 VDD.n12111 9.3
R6783 VDD.n12100 VDD.n12099 9.3
R6784 VDD.n12099 VDD.n12098 9.3
R6785 VDD.n12084 VDD.n12083 9.3
R6786 VDD.n12080 VDD.n12079 9.3
R6787 VDD.n12079 VDD.n12078 9.3
R6788 VDD.n12072 VDD.n12071 9.3
R6789 VDD.n12068 VDD.n12067 9.3
R6790 VDD.n12067 VDD.n12066 9.3
R6791 VDD.n12059 VDD.n12058 9.3
R6792 VDD.n12055 VDD.n12054 9.3
R6793 VDD.n12054 VDD.n12053 9.3
R6794 VDD.n12047 VDD.n12046 9.3
R6795 VDD.n12043 VDD.n12042 9.3
R6796 VDD.n12042 VDD.n12041 9.3
R6797 VDD.n12034 VDD.n12033 9.3
R6798 VDD.n12030 VDD.n12029 9.3
R6799 VDD.n12029 VDD.n12028 9.3
R6800 VDD.n12022 VDD.n12021 9.3
R6801 VDD.n12018 VDD.n12017 9.3
R6802 VDD.n12017 VDD.n12016 9.3
R6803 VDD.n12009 VDD.n12008 9.3
R6804 VDD.n12005 VDD.n12004 9.3
R6805 VDD.n12004 VDD.n12003 9.3
R6806 VDD.n11997 VDD.n11996 9.3
R6807 VDD.n11993 VDD.n11992 9.3
R6808 VDD.n11992 VDD.n11991 9.3
R6809 VDD.n11984 VDD.n11983 9.3
R6810 VDD.n11983 VDD.n11982 9.3
R6811 VDD.n11971 VDD.n11970 9.3
R6812 VDD.n11970 VDD.n11969 9.3
R6813 VDD.n11958 VDD.n11957 9.3
R6814 VDD.n11198 VDD.n11197 9.3
R6815 VDD.n11211 VDD.n11210 9.3
R6816 VDD.n11229 VDD.n11228 9.3
R6817 VDD.n11241 VDD.n11240 9.3
R6818 VDD.n11253 VDD.n11252 9.3
R6819 VDD.n11265 VDD.n11264 9.3
R6820 VDD.n11277 VDD.n11276 9.3
R6821 VDD.n11289 VDD.n11288 9.3
R6822 VDD.n11301 VDD.n11300 9.3
R6823 VDD.n11313 VDD.n11312 9.3
R6824 VDD.n11323 VDD.n11322 9.3
R6825 VDD.n11337 VDD.n11336 9.3
R6826 VDD.n11349 VDD.n11348 9.3
R6827 VDD.n11361 VDD.n11360 9.3
R6828 VDD.n11373 VDD.n11372 9.3
R6829 VDD.n11385 VDD.n11384 9.3
R6830 VDD.n11397 VDD.n11396 9.3
R6831 VDD.n11409 VDD.n11408 9.3
R6832 VDD.n11427 VDD.n11426 9.3
R6833 VDD.n11439 VDD.n11438 9.3
R6834 VDD.n11451 VDD.n11450 9.3
R6835 VDD.n11196 VDD.n11195 9.3
R6836 VDD.n11209 VDD.n11208 9.3
R6837 VDD.n11321 VDD.n11320 9.3
R6838 VDD.n11335 VDD.n11334 9.3
R6839 VDD.n11347 VDD.n11346 9.3
R6840 VDD.n11359 VDD.n11358 9.3
R6841 VDD.n11371 VDD.n11370 9.3
R6842 VDD.n11383 VDD.n11382 9.3
R6843 VDD.n11395 VDD.n11394 9.3
R6844 VDD.n11407 VDD.n11406 9.3
R6845 VDD.n11453 VDD.n11452 9.3
R6846 VDD.n11449 VDD.n11448 9.3
R6847 VDD.n11448 VDD.n11447 9.3
R6848 VDD.n11441 VDD.n11440 9.3
R6849 VDD.n11437 VDD.n11436 9.3
R6850 VDD.n11436 VDD.n11435 9.3
R6851 VDD.n11429 VDD.n11428 9.3
R6852 VDD.n11425 VDD.n11424 9.3
R6853 VDD.n11424 VDD.n11423 9.3
R6854 VDD.n11417 VDD.n11416 9.3
R6855 VDD.n11416 VDD.n11415 9.3
R6856 VDD.n11405 VDD.n11404 9.3
R6857 VDD.n11404 VDD.n11403 9.3
R6858 VDD.n11393 VDD.n11392 9.3
R6859 VDD.n11392 VDD.n11391 9.3
R6860 VDD.n11381 VDD.n11380 9.3
R6861 VDD.n11380 VDD.n11379 9.3
R6862 VDD.n11369 VDD.n11368 9.3
R6863 VDD.n11368 VDD.n11367 9.3
R6864 VDD.n11357 VDD.n11356 9.3
R6865 VDD.n11356 VDD.n11355 9.3
R6866 VDD.n11345 VDD.n11344 9.3
R6867 VDD.n11344 VDD.n11343 9.3
R6868 VDD.n11333 VDD.n11332 9.3
R6869 VDD.n11332 VDD.n11331 9.3
R6870 VDD.n11315 VDD.n11314 9.3
R6871 VDD.n11311 VDD.n11310 9.3
R6872 VDD.n11310 VDD.n11309 9.3
R6873 VDD.n11303 VDD.n11302 9.3
R6874 VDD.n11299 VDD.n11298 9.3
R6875 VDD.n11298 VDD.n11297 9.3
R6876 VDD.n11291 VDD.n11290 9.3
R6877 VDD.n11287 VDD.n11286 9.3
R6878 VDD.n11286 VDD.n11285 9.3
R6879 VDD.n11279 VDD.n11278 9.3
R6880 VDD.n11275 VDD.n11274 9.3
R6881 VDD.n11274 VDD.n11273 9.3
R6882 VDD.n11267 VDD.n11266 9.3
R6883 VDD.n11263 VDD.n11262 9.3
R6884 VDD.n11262 VDD.n11261 9.3
R6885 VDD.n11255 VDD.n11254 9.3
R6886 VDD.n11251 VDD.n11250 9.3
R6887 VDD.n11250 VDD.n11249 9.3
R6888 VDD.n11243 VDD.n11242 9.3
R6889 VDD.n11239 VDD.n11238 9.3
R6890 VDD.n11238 VDD.n11237 9.3
R6891 VDD.n11231 VDD.n11230 9.3
R6892 VDD.n11227 VDD.n11226 9.3
R6893 VDD.n11226 VDD.n11225 9.3
R6894 VDD.n11219 VDD.n11218 9.3
R6895 VDD.n11218 VDD.n11217 9.3
R6896 VDD.n11207 VDD.n11206 9.3
R6897 VDD.n11206 VDD.n11205 9.3
R6898 VDD.n11193 VDD.n11192 9.3
R6899 VDD.n12242 VDD.n12241 9.3
R6900 VDD.n12236 VDD.n12235 9.3
R6901 VDD.n12238 VDD.n12237 9.3
R6902 VDD.n12315 VDD.n12314 9.3
R6903 VDD.n12302 VDD.n12301 9.3
R6904 VDD.n12283 VDD.n12282 9.3
R6905 VDD.n12270 VDD.n12269 9.3
R6906 VDD.n12313 VDD.n12312 9.3
R6907 VDD.n12312 VDD.n12311 9.3
R6908 VDD.n12304 VDD.n12303 9.3
R6909 VDD.n12300 VDD.n12299 9.3
R6910 VDD.n12299 VDD.n12298 9.3
R6911 VDD.n12281 VDD.n12280 9.3
R6912 VDD.n12291 VDD.n12290 9.3
R6913 VDD.n12290 VDD.n12289 9.3
R6914 VDD.n12268 VDD.n12267 9.3
R6915 VDD.n12279 VDD.n12278 9.3
R6916 VDD.n12278 VDD.n12277 9.3
R6917 VDD.n12317 VDD.n12316 9.3
R6918 VDD.n2785 VDD.n2784 9.249
R6919 VDD.n10404 VDD.t36 9.245
R6920 VDD.n2123 VDD.n2122 9.23
R6921 VDD.n2200 VDD.n2199 9.23
R6922 VDD.n2354 VDD.n2353 9.23
R6923 VDD.n2431 VDD.n2430 9.23
R6924 VDD.n5175 VDD.n5174 9.23
R6925 VDD.n5242 VDD.n5241 9.23
R6926 VDD.n5035 VDD.n5034 9.23
R6927 VDD.n4958 VDD.n4957 9.23
R6928 VDD.n4804 VDD.n4803 9.23
R6929 VDD.n4727 VDD.n4726 9.23
R6930 VDD.n10348 VDD.t57 9.217
R6931 VDD.n10430 VDD.t55 9.206
R6932 VDD.n10377 VDD.t40 9.206
R6933 VDD.n11391 VDD.n11390 9.09
R6934 VDD.n11192 VDD.n11191 9.09
R6935 VDD.n12219 VDD.n12218 9.09
R6936 VDD.n12161 VDD.n12159 9.09
R6937 VDD.n12016 VDD.n12014 9.09
R6938 VDD.n11957 VDD.n11956 9.09
R6939 VDD.n10880 VDD.n10878 9.09
R6940 VDD.n10991 VDD.n10989 9.09
R6941 VDD.n11132 VDD.n11123 9.09
R6942 VDD.n10706 VDD.n10704 9.09
R6943 VDD.n11862 VDD.n11860 9.09
R6944 VDD.n2799 VDD.n2798 9.013
R6945 VDD.n2953 VDD.n2952 9.013
R6946 VDD.n4460 VDD.n4459 9.013
R6947 VDD.n4566 VDD.n4565 9.013
R6948 VDD.n1963 VDD.n1962 9.013
R6949 VDD.n1856 VDD.n1855 9.013
R6950 VDD.n221 VDD.n220 9.013
R6951 VDD.n370 VDD.n369 9.013
R6952 VDD.n2834 VDD.n2833 9
R6953 VDD.n3092 VDD.n3091 9
R6954 VDD.n3137 VDD.n3136 9
R6955 VDD.n3330 VDD.n3329 9
R6956 VDD.n3375 VDD.n3374 9
R6957 VDD.n3567 VDD.n3566 9
R6958 VDD.n3612 VDD.n3611 9
R6959 VDD.n3805 VDD.n3804 9
R6960 VDD.n3850 VDD.n3849 9
R6961 VDD.n4042 VDD.n4041 9
R6962 VDD.n4087 VDD.n4086 9
R6963 VDD.n4280 VDD.n4279 9
R6964 VDD.n4325 VDD.n4324 9
R6965 VDD.n4554 VDD.n4553 9
R6966 VDD.n10153 VDD.n10152 8.888
R6967 VDD.n10071 VDD.n10070 8.888
R6968 VDD.n10019 VDD.n10017 8.888
R6969 VDD.n214 VDD.n213 8.855
R6970 VDD.n255 VDD.n254 8.855
R6971 VDD.n254 VDD.n253 8.855
R6972 VDD.n278 VDD.n277 8.855
R6973 VDD.n277 VDD.n276 8.855
R6974 VDD.n309 VDD.n308 8.855
R6975 VDD.n308 VDD.n307 8.855
R6976 VDD.n327 VDD.n326 8.855
R6977 VDD.n326 VDD.n325 8.855
R6978 VDD.n378 VDD.n377 8.855
R6979 VDD.n377 VDD.n376 8.855
R6980 VDD.n392 VDD.n391 8.855
R6981 VDD.n391 VDD.n390 8.855
R6982 VDD.n406 VDD.n405 8.855
R6983 VDD.n405 VDD.n404 8.855
R6984 VDD.n421 VDD.n420 8.855
R6985 VDD.n420 VDD.n419 8.855
R6986 VDD.n433 VDD.n432 8.855
R6987 VDD.n432 VDD.n431 8.855
R6988 VDD.n447 VDD.n446 8.855
R6989 VDD.n446 VDD.n445 8.855
R6990 VDD.n461 VDD.n460 8.855
R6991 VDD.n460 VDD.n459 8.855
R6992 VDD.n475 VDD.n474 8.855
R6993 VDD.n474 VDD.n473 8.855
R6994 VDD.n489 VDD.n488 8.855
R6995 VDD.n488 VDD.n487 8.855
R6996 VDD.n503 VDD.n502 8.855
R6997 VDD.n502 VDD.n501 8.855
R6998 VDD.n517 VDD.n516 8.855
R6999 VDD.n516 VDD.n515 8.855
R7000 VDD.n531 VDD.n530 8.855
R7001 VDD.n530 VDD.n529 8.855
R7002 VDD.n555 VDD.n554 8.855
R7003 VDD.n554 VDD.n553 8.855
R7004 VDD.n570 VDD.n569 8.855
R7005 VDD.n569 VDD.n568 8.855
R7006 VDD.n584 VDD.n583 8.855
R7007 VDD.n583 VDD.n582 8.855
R7008 VDD.n598 VDD.n597 8.855
R7009 VDD.n597 VDD.n596 8.855
R7010 VDD.n612 VDD.n611 8.855
R7011 VDD.n611 VDD.n610 8.855
R7012 VDD.n626 VDD.n625 8.855
R7013 VDD.n625 VDD.n624 8.855
R7014 VDD.n640 VDD.n639 8.855
R7015 VDD.n639 VDD.n638 8.855
R7016 VDD.n654 VDD.n653 8.855
R7017 VDD.n653 VDD.n652 8.855
R7018 VDD.n666 VDD.n665 8.855
R7019 VDD.n665 VDD.n664 8.855
R7020 VDD.n680 VDD.n679 8.855
R7021 VDD.n679 VDD.n678 8.855
R7022 VDD.n694 VDD.n693 8.855
R7023 VDD.n693 VDD.n692 8.855
R7024 VDD.n708 VDD.n707 8.855
R7025 VDD.n707 VDD.n706 8.855
R7026 VDD.n722 VDD.n721 8.855
R7027 VDD.n721 VDD.n720 8.855
R7028 VDD.n737 VDD.n736 8.855
R7029 VDD.n736 VDD.n735 8.855
R7030 VDD.n751 VDD.n750 8.855
R7031 VDD.n750 VDD.n749 8.855
R7032 VDD.n765 VDD.n764 8.855
R7033 VDD.n764 VDD.n763 8.855
R7034 VDD.n789 VDD.n788 8.855
R7035 VDD.n788 VDD.n787 8.855
R7036 VDD.n803 VDD.n802 8.855
R7037 VDD.n802 VDD.n801 8.855
R7038 VDD.n817 VDD.n816 8.855
R7039 VDD.n816 VDD.n815 8.855
R7040 VDD.n831 VDD.n830 8.855
R7041 VDD.n830 VDD.n829 8.855
R7042 VDD.n845 VDD.n844 8.855
R7043 VDD.n844 VDD.n843 8.855
R7044 VDD.n859 VDD.n858 8.855
R7045 VDD.n858 VDD.n857 8.855
R7046 VDD.n873 VDD.n872 8.855
R7047 VDD.n872 VDD.n871 8.855
R7048 VDD.n888 VDD.n887 8.855
R7049 VDD.n887 VDD.n886 8.855
R7050 VDD.n900 VDD.n899 8.855
R7051 VDD.n899 VDD.n898 8.855
R7052 VDD.n914 VDD.n913 8.855
R7053 VDD.n913 VDD.n912 8.855
R7054 VDD.n928 VDD.n927 8.855
R7055 VDD.n927 VDD.n926 8.855
R7056 VDD.n942 VDD.n941 8.855
R7057 VDD.n941 VDD.n940 8.855
R7058 VDD.n956 VDD.n955 8.855
R7059 VDD.n955 VDD.n954 8.855
R7060 VDD.n970 VDD.n969 8.855
R7061 VDD.n969 VDD.n968 8.855
R7062 VDD.n984 VDD.n983 8.855
R7063 VDD.n983 VDD.n982 8.855
R7064 VDD.n998 VDD.n997 8.855
R7065 VDD.n997 VDD.n996 8.855
R7066 VDD.n1022 VDD.n1021 8.855
R7067 VDD.n1021 VDD.n1020 8.855
R7068 VDD.n1037 VDD.n1036 8.855
R7069 VDD.n1036 VDD.n1035 8.855
R7070 VDD.n1051 VDD.n1050 8.855
R7071 VDD.n1050 VDD.n1049 8.855
R7072 VDD.n1065 VDD.n1064 8.855
R7073 VDD.n1064 VDD.n1063 8.855
R7074 VDD.n1079 VDD.n1078 8.855
R7075 VDD.n1078 VDD.n1077 8.855
R7076 VDD.n1093 VDD.n1092 8.855
R7077 VDD.n1092 VDD.n1091 8.855
R7078 VDD.n1107 VDD.n1106 8.855
R7079 VDD.n1106 VDD.n1105 8.855
R7080 VDD.n1121 VDD.n1120 8.855
R7081 VDD.n1120 VDD.n1119 8.855
R7082 VDD.n1133 VDD.n1132 8.855
R7083 VDD.n1132 VDD.n1131 8.855
R7084 VDD.n1147 VDD.n1146 8.855
R7085 VDD.n1146 VDD.n1145 8.855
R7086 VDD.n1161 VDD.n1160 8.855
R7087 VDD.n1160 VDD.n1159 8.855
R7088 VDD.n1175 VDD.n1174 8.855
R7089 VDD.n1174 VDD.n1173 8.855
R7090 VDD.n1189 VDD.n1188 8.855
R7091 VDD.n1188 VDD.n1187 8.855
R7092 VDD.n1204 VDD.n1203 8.855
R7093 VDD.n1203 VDD.n1202 8.855
R7094 VDD.n1218 VDD.n1217 8.855
R7095 VDD.n1217 VDD.n1216 8.855
R7096 VDD.n1232 VDD.n1231 8.855
R7097 VDD.n1231 VDD.n1230 8.855
R7098 VDD.n1256 VDD.n1255 8.855
R7099 VDD.n1255 VDD.n1254 8.855
R7100 VDD.n1270 VDD.n1269 8.855
R7101 VDD.n1269 VDD.n1268 8.855
R7102 VDD.n1284 VDD.n1283 8.855
R7103 VDD.n1283 VDD.n1282 8.855
R7104 VDD.n1298 VDD.n1297 8.855
R7105 VDD.n1297 VDD.n1296 8.855
R7106 VDD.n1312 VDD.n1311 8.855
R7107 VDD.n1311 VDD.n1310 8.855
R7108 VDD.n1326 VDD.n1325 8.855
R7109 VDD.n1325 VDD.n1324 8.855
R7110 VDD.n1340 VDD.n1339 8.855
R7111 VDD.n1339 VDD.n1338 8.855
R7112 VDD.n1355 VDD.n1354 8.855
R7113 VDD.n1354 VDD.n1353 8.855
R7114 VDD.n1367 VDD.n1366 8.855
R7115 VDD.n1366 VDD.n1365 8.855
R7116 VDD.n1381 VDD.n1380 8.855
R7117 VDD.n1380 VDD.n1379 8.855
R7118 VDD.n1395 VDD.n1394 8.855
R7119 VDD.n1394 VDD.n1393 8.855
R7120 VDD.n1409 VDD.n1408 8.855
R7121 VDD.n1408 VDD.n1407 8.855
R7122 VDD.n1423 VDD.n1422 8.855
R7123 VDD.n1422 VDD.n1421 8.855
R7124 VDD.n1437 VDD.n1436 8.855
R7125 VDD.n1436 VDD.n1435 8.855
R7126 VDD.n1451 VDD.n1450 8.855
R7127 VDD.n1450 VDD.n1449 8.855
R7128 VDD.n1465 VDD.n1464 8.855
R7129 VDD.n1464 VDD.n1463 8.855
R7130 VDD.n1489 VDD.n1488 8.855
R7131 VDD.n1488 VDD.n1487 8.855
R7132 VDD.n1504 VDD.n1503 8.855
R7133 VDD.n1503 VDD.n1502 8.855
R7134 VDD.n1518 VDD.n1517 8.855
R7135 VDD.n1517 VDD.n1516 8.855
R7136 VDD.n1532 VDD.n1531 8.855
R7137 VDD.n1531 VDD.n1530 8.855
R7138 VDD.n1546 VDD.n1545 8.855
R7139 VDD.n1545 VDD.n1544 8.855
R7140 VDD.n1560 VDD.n1559 8.855
R7141 VDD.n1559 VDD.n1558 8.855
R7142 VDD.n1574 VDD.n1573 8.855
R7143 VDD.n1573 VDD.n1572 8.855
R7144 VDD.n1588 VDD.n1587 8.855
R7145 VDD.n1587 VDD.n1586 8.855
R7146 VDD.n1600 VDD.n1599 8.855
R7147 VDD.n1599 VDD.n1598 8.855
R7148 VDD.n1614 VDD.n1613 8.855
R7149 VDD.n1613 VDD.n1612 8.855
R7150 VDD.n1628 VDD.n1627 8.855
R7151 VDD.n1627 VDD.n1626 8.855
R7152 VDD.n1642 VDD.n1641 8.855
R7153 VDD.n1641 VDD.n1640 8.855
R7154 VDD.n1656 VDD.n1655 8.855
R7155 VDD.n1655 VDD.n1654 8.855
R7156 VDD.n1671 VDD.n1670 8.855
R7157 VDD.n1670 VDD.n1669 8.855
R7158 VDD.n1685 VDD.n1684 8.855
R7159 VDD.n1684 VDD.n1683 8.855
R7160 VDD.n1699 VDD.n1698 8.855
R7161 VDD.n1698 VDD.n1697 8.855
R7162 VDD.n1723 VDD.n1722 8.855
R7163 VDD.n1722 VDD.n1721 8.855
R7164 VDD.n1737 VDD.n1736 8.855
R7165 VDD.n1736 VDD.n1735 8.855
R7166 VDD.n1751 VDD.n1750 8.855
R7167 VDD.n1750 VDD.n1749 8.855
R7168 VDD.n1765 VDD.n1764 8.855
R7169 VDD.n1764 VDD.n1763 8.855
R7170 VDD.n1779 VDD.n1778 8.855
R7171 VDD.n1778 VDD.n1777 8.855
R7172 VDD.n1793 VDD.n1792 8.855
R7173 VDD.n1792 VDD.n1791 8.855
R7174 VDD.n1807 VDD.n1806 8.855
R7175 VDD.n1806 VDD.n1805 8.855
R7176 VDD.n1822 VDD.n1821 8.855
R7177 VDD.n1821 VDD.n1820 8.855
R7178 VDD.n1834 VDD.n1833 8.855
R7179 VDD.n1833 VDD.n1832 8.855
R7180 VDD.n1848 VDD.n1847 8.855
R7181 VDD.n1847 VDD.n1846 8.855
R7182 VDD.n1884 VDD.n1883 8.855
R7183 VDD.n1883 VDD.n1882 8.855
R7184 VDD.n1903 VDD.n1902 8.855
R7185 VDD.n1902 VDD.n1901 8.855
R7186 VDD.n1922 VDD.n1921 8.855
R7187 VDD.n1921 VDD.n1920 8.855
R7188 VDD.n1866 VDD.n1865 8.855
R7189 VDD.n1865 VDD.n1864 8.855
R7190 VDD.n1944 VDD.n1943 8.855
R7191 VDD.n1943 VDD.n1942 8.855
R7192 VDD.n2017 VDD.n2016 8.855
R7193 VDD.n2016 VDD.n2015 8.855
R7194 VDD.n4628 VDD.n4627 8.855
R7195 VDD.n4629 VDD.n4628 8.855
R7196 VDD.n2975 VDD.n2974 8.855
R7197 VDD.n2974 VDD.n2973 8.855
R7198 VDD.n2989 VDD.n2988 8.855
R7199 VDD.n2988 VDD.n2987 8.855
R7200 VDD.n3128 VDD.n3127 8.855
R7201 VDD.n3127 VDD.n3126 8.855
R7202 VDD.n3142 VDD.n3141 8.855
R7203 VDD.n3141 VDD.n3140 8.855
R7204 VDD.n3157 VDD.n3156 8.855
R7205 VDD.n3156 VDD.n3155 8.855
R7206 VDD.n3171 VDD.n3170 8.855
R7207 VDD.n3170 VDD.n3169 8.855
R7208 VDD.n3185 VDD.n3184 8.855
R7209 VDD.n3184 VDD.n3183 8.855
R7210 VDD.n3199 VDD.n3198 8.855
R7211 VDD.n3198 VDD.n3197 8.855
R7212 VDD.n3213 VDD.n3212 8.855
R7213 VDD.n3212 VDD.n3211 8.855
R7214 VDD.n3227 VDD.n3226 8.855
R7215 VDD.n3226 VDD.n3225 8.855
R7216 VDD.n3366 VDD.n3365 8.855
R7217 VDD.n3365 VDD.n3364 8.855
R7218 VDD.n3380 VDD.n3379 8.855
R7219 VDD.n3379 VDD.n3378 8.855
R7220 VDD.n3394 VDD.n3393 8.855
R7221 VDD.n3393 VDD.n3392 8.855
R7222 VDD.n3408 VDD.n3407 8.855
R7223 VDD.n3407 VDD.n3406 8.855
R7224 VDD.n3422 VDD.n3421 8.855
R7225 VDD.n3421 VDD.n3420 8.855
R7226 VDD.n3436 VDD.n3435 8.855
R7227 VDD.n3435 VDD.n3434 8.855
R7228 VDD.n3450 VDD.n3449 8.855
R7229 VDD.n3449 VDD.n3448 8.855
R7230 VDD.n3464 VDD.n3463 8.855
R7231 VDD.n3463 VDD.n3462 8.855
R7232 VDD.n3603 VDD.n3602 8.855
R7233 VDD.n3602 VDD.n3601 8.855
R7234 VDD.n3617 VDD.n3616 8.855
R7235 VDD.n3616 VDD.n3615 8.855
R7236 VDD.n3632 VDD.n3631 8.855
R7237 VDD.n3631 VDD.n3630 8.855
R7238 VDD.n3646 VDD.n3645 8.855
R7239 VDD.n3645 VDD.n3644 8.855
R7240 VDD.n3660 VDD.n3659 8.855
R7241 VDD.n3659 VDD.n3658 8.855
R7242 VDD.n3674 VDD.n3673 8.855
R7243 VDD.n3673 VDD.n3672 8.855
R7244 VDD.n3688 VDD.n3687 8.855
R7245 VDD.n3687 VDD.n3686 8.855
R7246 VDD.n3702 VDD.n3701 8.855
R7247 VDD.n3701 VDD.n3700 8.855
R7248 VDD.n3841 VDD.n3840 8.855
R7249 VDD.n3840 VDD.n3839 8.855
R7250 VDD.n3855 VDD.n3854 8.855
R7251 VDD.n3854 VDD.n3853 8.855
R7252 VDD.n3869 VDD.n3868 8.855
R7253 VDD.n3868 VDD.n3867 8.855
R7254 VDD.n3883 VDD.n3882 8.855
R7255 VDD.n3882 VDD.n3881 8.855
R7256 VDD.n3897 VDD.n3896 8.855
R7257 VDD.n3896 VDD.n3895 8.855
R7258 VDD.n3911 VDD.n3910 8.855
R7259 VDD.n3910 VDD.n3909 8.855
R7260 VDD.n3925 VDD.n3924 8.855
R7261 VDD.n3924 VDD.n3923 8.855
R7262 VDD.n3939 VDD.n3938 8.855
R7263 VDD.n3938 VDD.n3937 8.855
R7264 VDD.n4078 VDD.n4077 8.855
R7265 VDD.n4077 VDD.n4076 8.855
R7266 VDD.n4092 VDD.n4091 8.855
R7267 VDD.n4091 VDD.n4090 8.855
R7268 VDD.n4107 VDD.n4106 8.855
R7269 VDD.n4106 VDD.n4105 8.855
R7270 VDD.n4121 VDD.n4120 8.855
R7271 VDD.n4120 VDD.n4119 8.855
R7272 VDD.n4135 VDD.n4134 8.855
R7273 VDD.n4134 VDD.n4133 8.855
R7274 VDD.n4149 VDD.n4148 8.855
R7275 VDD.n4148 VDD.n4147 8.855
R7276 VDD.n4163 VDD.n4162 8.855
R7277 VDD.n4162 VDD.n4161 8.855
R7278 VDD.n4177 VDD.n4176 8.855
R7279 VDD.n4176 VDD.n4175 8.855
R7280 VDD.n4316 VDD.n4315 8.855
R7281 VDD.n4315 VDD.n4314 8.855
R7282 VDD.n4330 VDD.n4329 8.855
R7283 VDD.n4329 VDD.n4328 8.855
R7284 VDD.n4344 VDD.n4343 8.855
R7285 VDD.n4343 VDD.n4342 8.855
R7286 VDD.n4358 VDD.n4357 8.855
R7287 VDD.n4357 VDD.n4356 8.855
R7288 VDD.n4372 VDD.n4371 8.855
R7289 VDD.n4371 VDD.n4370 8.855
R7290 VDD.n4386 VDD.n4385 8.855
R7291 VDD.n4385 VDD.n4384 8.855
R7292 VDD.n4400 VDD.n4399 8.855
R7293 VDD.n4399 VDD.n4398 8.855
R7294 VDD.n4414 VDD.n4413 8.855
R7295 VDD.n4413 VDD.n4412 8.855
R7296 VDD.n4559 VDD.n4558 8.855
R7297 VDD.n4558 VDD.n4557 8.855
R7298 VDD.n4511 VDD.n4510 8.855
R7299 VDD.n4510 VDD.n4509 8.855
R7300 VDD.n2961 VDD.n2960 8.855
R7301 VDD.n2960 VDD.n2959 8.855
R7302 VDD.n2895 VDD.n2894 8.855
R7303 VDD.n2894 VDD.n2893 8.855
R7304 VDD.n2839 VDD.n2838 8.855
R7305 VDD.n2838 VDD.n2837 8.855
R7306 VDD.n2786 VDD.n2785 8.855
R7307 VDD.n2807 VDD.n2806 8.855
R7308 VDD.n2806 VDD.n2805 8.855
R7309 VDD.n2865 VDD.n2864 8.855
R7310 VDD.n2864 VDD.n2863 8.855
R7311 VDD.n2914 VDD.n2913 8.855
R7312 VDD.n2913 VDD.n2912 8.855
R7313 VDD.n3013 VDD.n3012 8.855
R7314 VDD.n3012 VDD.n3011 8.855
R7315 VDD.n3027 VDD.n3026 8.855
R7316 VDD.n3026 VDD.n3025 8.855
R7317 VDD.n3041 VDD.n3040 8.855
R7318 VDD.n3040 VDD.n3039 8.855
R7319 VDD.n3055 VDD.n3054 8.855
R7320 VDD.n3054 VDD.n3053 8.855
R7321 VDD.n3069 VDD.n3068 8.855
R7322 VDD.n3068 VDD.n3067 8.855
R7323 VDD.n3083 VDD.n3082 8.855
R7324 VDD.n3082 VDD.n3081 8.855
R7325 VDD.n3097 VDD.n3096 8.855
R7326 VDD.n3096 VDD.n3095 8.855
R7327 VDD.n3111 VDD.n3110 8.855
R7328 VDD.n3110 VDD.n3109 8.855
R7329 VDD.n3250 VDD.n3249 8.855
R7330 VDD.n3249 VDD.n3248 8.855
R7331 VDD.n3264 VDD.n3263 8.855
R7332 VDD.n3263 VDD.n3262 8.855
R7333 VDD.n3278 VDD.n3277 8.855
R7334 VDD.n3277 VDD.n3276 8.855
R7335 VDD.n3292 VDD.n3291 8.855
R7336 VDD.n3291 VDD.n3290 8.855
R7337 VDD.n3306 VDD.n3305 8.855
R7338 VDD.n3305 VDD.n3304 8.855
R7339 VDD.n3321 VDD.n3320 8.855
R7340 VDD.n3320 VDD.n3319 8.855
R7341 VDD.n3335 VDD.n3334 8.855
R7342 VDD.n3334 VDD.n3333 8.855
R7343 VDD.n3349 VDD.n3348 8.855
R7344 VDD.n3348 VDD.n3347 8.855
R7345 VDD.n3488 VDD.n3487 8.855
R7346 VDD.n3487 VDD.n3486 8.855
R7347 VDD.n3502 VDD.n3501 8.855
R7348 VDD.n3501 VDD.n3500 8.855
R7349 VDD.n3516 VDD.n3515 8.855
R7350 VDD.n3515 VDD.n3514 8.855
R7351 VDD.n3530 VDD.n3529 8.855
R7352 VDD.n3529 VDD.n3528 8.855
R7353 VDD.n3544 VDD.n3543 8.855
R7354 VDD.n3543 VDD.n3542 8.855
R7355 VDD.n3558 VDD.n3557 8.855
R7356 VDD.n3557 VDD.n3556 8.855
R7357 VDD.n3572 VDD.n3571 8.855
R7358 VDD.n3571 VDD.n3570 8.855
R7359 VDD.n3586 VDD.n3585 8.855
R7360 VDD.n3585 VDD.n3584 8.855
R7361 VDD.n3725 VDD.n3724 8.855
R7362 VDD.n3724 VDD.n3723 8.855
R7363 VDD.n3739 VDD.n3738 8.855
R7364 VDD.n3738 VDD.n3737 8.855
R7365 VDD.n3753 VDD.n3752 8.855
R7366 VDD.n3752 VDD.n3751 8.855
R7367 VDD.n3767 VDD.n3766 8.855
R7368 VDD.n3766 VDD.n3765 8.855
R7369 VDD.n3781 VDD.n3780 8.855
R7370 VDD.n3780 VDD.n3779 8.855
R7371 VDD.n3796 VDD.n3795 8.855
R7372 VDD.n3795 VDD.n3794 8.855
R7373 VDD.n3810 VDD.n3809 8.855
R7374 VDD.n3809 VDD.n3808 8.855
R7375 VDD.n3824 VDD.n3823 8.855
R7376 VDD.n3823 VDD.n3822 8.855
R7377 VDD.n3963 VDD.n3962 8.855
R7378 VDD.n3962 VDD.n3961 8.855
R7379 VDD.n3977 VDD.n3976 8.855
R7380 VDD.n3976 VDD.n3975 8.855
R7381 VDD.n3991 VDD.n3990 8.855
R7382 VDD.n3990 VDD.n3989 8.855
R7383 VDD.n4005 VDD.n4004 8.855
R7384 VDD.n4004 VDD.n4003 8.855
R7385 VDD.n4019 VDD.n4018 8.855
R7386 VDD.n4018 VDD.n4017 8.855
R7387 VDD.n4033 VDD.n4032 8.855
R7388 VDD.n4032 VDD.n4031 8.855
R7389 VDD.n4047 VDD.n4046 8.855
R7390 VDD.n4046 VDD.n4045 8.855
R7391 VDD.n4061 VDD.n4060 8.855
R7392 VDD.n4060 VDD.n4059 8.855
R7393 VDD.n4200 VDD.n4199 8.855
R7394 VDD.n4199 VDD.n4198 8.855
R7395 VDD.n4214 VDD.n4213 8.855
R7396 VDD.n4213 VDD.n4212 8.855
R7397 VDD.n4228 VDD.n4227 8.855
R7398 VDD.n4227 VDD.n4226 8.855
R7399 VDD.n4242 VDD.n4241 8.855
R7400 VDD.n4241 VDD.n4240 8.855
R7401 VDD.n4256 VDD.n4255 8.855
R7402 VDD.n4255 VDD.n4254 8.855
R7403 VDD.n4271 VDD.n4270 8.855
R7404 VDD.n4270 VDD.n4269 8.855
R7405 VDD.n4285 VDD.n4284 8.855
R7406 VDD.n4284 VDD.n4283 8.855
R7407 VDD.n4299 VDD.n4298 8.855
R7408 VDD.n4298 VDD.n4297 8.855
R7409 VDD.n4438 VDD.n4437 8.855
R7410 VDD.n4437 VDD.n4436 8.855
R7411 VDD.n4452 VDD.n4451 8.855
R7412 VDD.n4451 VDD.n4450 8.855
R7413 VDD.n4471 VDD.n4470 8.855
R7414 VDD.n4470 VDD.n4469 8.855
R7415 VDD.n4491 VDD.n4490 8.855
R7416 VDD.n4490 VDD.n4489 8.855
R7417 VDD.n4531 VDD.n4530 8.855
R7418 VDD.n4530 VDD.n4529 8.855
R7419 VDD.n4622 VDD.n4621 8.855
R7420 VDD.n4621 VDD.n4620 8.855
R7421 VDD.n4883 VDD.n4882 8.855
R7422 VDD.n4882 VDD.n4881 8.855
R7423 VDD.n4652 VDD.n4651 8.855
R7424 VDD.n4651 VDD.n4650 8.855
R7425 VDD.n2048 VDD.n2047 8.855
R7426 VDD.n2047 VDD.n2046 8.855
R7427 VDD.n2279 VDD.n2278 8.855
R7428 VDD.n2278 VDD.n2277 8.855
R7429 VDD.n2523 VDD.n2522 8.855
R7430 VDD.n2522 VDD.n2521 8.855
R7431 VDD.n2762 VDD.n2761 8.855
R7432 VDD.n2761 VDD.n2760 8.855
R7433 VDD.n10288 VDD.n10287 8.855
R7434 VDD.n10170 VDD.n10169 8.855
R7435 VDD.n10087 VDD.n10086 8.855
R7436 VDD.n10043 VDD.n10042 8.855
R7437 VDD.n10635 VDD.n10634 8.855
R7438 VDD.n10516 VDD.n10515 8.855
R7439 VDD.n10308 VDD.n10306 8.727
R7440 VDD.n10655 VDD.n10653 8.727
R7441 VDD.n10499 VDD.n10498 8.727
R7442 VDD.n11378 VDD.n11377 8.665
R7443 VDD.n11656 VDD.n11655 8.665
R7444 VDD.n11868 VDD.n11867 8.665
R7445 VDD.n11655 VDD.n11654 8.665
R7446 VDD.n11867 VDD.n11866 8.665
R7447 VDD.n11377 VDD.n11376 8.665
R7448 VDD.n2164 VDD.n2163 8.615
R7449 VDD.n2395 VDD.n2394 8.615
R7450 VDD.n4999 VDD.n4998 8.615
R7451 VDD.n4768 VDD.n4767 8.615
R7452 VDD.n10883 VDD.n10882 8.55
R7453 VDD.n10709 VDD.n10708 8.55
R7454 VDD.n11652 VDD.n11651 8.55
R7455 VDD.n11479 VDD.n11478 8.55
R7456 VDD.n4633 VDD.n4632 8.531
R7457 VDD.n10063 VDD.n10062 8.468
R7458 VDD.n28 VDD.n27 8.46
R7459 VDD.n12259 VDD.n12258 8.46
R7460 VDD.n5382 VDD.n5381 8.454
R7461 VDD.n5743 VDD.n5742 8.454
R7462 VDD.n6105 VDD.n6104 8.454
R7463 VDD.n6467 VDD.n6466 8.454
R7464 VDD.n6829 VDD.n6828 8.454
R7465 VDD.n7191 VDD.n7190 8.454
R7466 VDD.n7553 VDD.n7552 8.454
R7467 VDD.n7915 VDD.n7914 8.454
R7468 VDD.n8277 VDD.n8276 8.454
R7469 VDD.n8639 VDD.n8638 8.454
R7470 VDD.n9001 VDD.n9000 8.454
R7471 VDD.n9363 VDD.n9362 8.454
R7472 VDD.n9725 VDD.n9724 8.454
R7473 VDD.n5666 VDD.n5665 8.453
R7474 VDD.n6027 VDD.n6026 8.453
R7475 VDD.n6389 VDD.n6388 8.453
R7476 VDD.n6751 VDD.n6750 8.453
R7477 VDD.n7113 VDD.n7112 8.453
R7478 VDD.n7475 VDD.n7474 8.453
R7479 VDD.n7837 VDD.n7836 8.453
R7480 VDD.n8199 VDD.n8198 8.453
R7481 VDD.n8561 VDD.n8560 8.453
R7482 VDD.n8923 VDD.n8922 8.453
R7483 VDD.n9285 VDD.n9284 8.453
R7484 VDD.n9647 VDD.n9646 8.453
R7485 VDD.n10009 VDD.n10008 8.453
R7486 VDD.n3001 VDD.n3000 8.45
R7487 VDD.n3000 VDD.n2999 8.45
R7488 VDD.n3238 VDD.n3237 8.45
R7489 VDD.n3237 VDD.n3236 8.45
R7490 VDD.n3476 VDD.n3475 8.45
R7491 VDD.n3475 VDD.n3474 8.45
R7492 VDD.n3713 VDD.n3712 8.45
R7493 VDD.n3712 VDD.n3711 8.45
R7494 VDD.n3951 VDD.n3950 8.45
R7495 VDD.n3950 VDD.n3949 8.45
R7496 VDD.n4188 VDD.n4187 8.45
R7497 VDD.n4187 VDD.n4186 8.45
R7498 VDD.n4426 VDD.n4425 8.45
R7499 VDD.n4425 VDD.n4424 8.45
R7500 VDD.n11457 VDD.n11456 8.45
R7501 VDD.n273 VDD.n272 8.275
R7502 VDD.n512 VDD.n511 8.275
R7503 VDD.n564 VDD.n563 8.275
R7504 VDD.n746 VDD.n745 8.275
R7505 VDD.n798 VDD.n797 8.275
R7506 VDD.n979 VDD.n978 8.275
R7507 VDD.n1031 VDD.n1030 8.275
R7508 VDD.n1213 VDD.n1212 8.275
R7509 VDD.n1265 VDD.n1264 8.275
R7510 VDD.n1446 VDD.n1445 8.275
R7511 VDD.n1498 VDD.n1497 8.275
R7512 VDD.n1680 VDD.n1679 8.275
R7513 VDD.n1732 VDD.n1731 8.275
R7514 VDD.n1939 VDD.n1938 8.275
R7515 VDD.n34 VDD.n33 8.269
R7516 VDD.n28 VDD.n26 8.269
R7517 VDD.n11446 VDD.n11445 8.269
R7518 VDD.n11248 VDD.n11247 8.269
R7519 VDD.n11759 VDD.n11758 8.269
R7520 VDD.n12265 VDD.n12264 8.269
R7521 VDD.n12259 VDD.n12257 8.269
R7522 VDD.n11949 VDD.n11948 8.258
R7523 VDD.n11458 VDD.n11457 8.258
R7524 VDD.n11462 VDD.n11461 8.17
R7525 VDD.n12229 VDD.n12228 8.126
R7526 VDD.n10188 VDD.n10187 8.093
R7527 VDD.n10063 VDD.n10061 8.093
R7528 VDD.n10025 VDD.n10024 8.093
R7529 VDD.n10226 VDD.n10225 7.961
R7530 VDD.n10573 VDD.n10572 7.961
R7531 VDD.n10269 VDD.n10268 7.953
R7532 VDD.n10616 VDD.n10615 7.953
R7533 VDD.n10534 VDD.n10533 7.953
R7534 VDD.n4626 VDD.n2774 7.886
R7535 VDD.n10107 VDD.n10106 7.464
R7536 VDD.n10108 VDD.n10107 7.464
R7537 VDD.n2030 VDD.n2024 7.384
R7538 VDD.n2071 VDD.n2067 7.384
R7539 VDD.n2260 VDD.n2256 7.384
R7540 VDD.n2302 VDD.n2298 7.384
R7541 VDD.n2493 VDD.n2489 7.384
R7542 VDD.n2559 VDD.n2555 7.384
R7543 VDD.n2720 VDD.n2716 7.384
R7544 VDD.n5096 VDD.n5092 7.384
R7545 VDD.n4906 VDD.n4902 7.384
R7546 VDD.n4864 VDD.n4860 7.384
R7547 VDD.n4675 VDD.n4671 7.384
R7548 VDD.n10232 VDD.n10231 7.334
R7549 VDD.n10233 VDD.n10232 7.334
R7550 VDD.n10579 VDD.n10578 7.334
R7551 VDD.n10580 VDD.n10579 7.334
R7552 VDD.n10453 VDD.n10452 7.334
R7553 VDD.n10454 VDD.n10453 7.334
R7554 VDD.n10103 VDD.n10057 7.279
R7555 VDD.n11295 VDD.n11294 7.272
R7556 VDD.n11814 VDD.n11813 7.272
R7557 VDD.n11522 VDD.n11521 7.272
R7558 VDD.n213 VDD.n212 7.136
R7559 VDD.n11366 VDD.n11365 6.998
R7560 VDD.n12133 VDD.n12132 6.998
R7561 VDD.n12039 VDD.n12038 6.998
R7562 VDD.n12134 VDD.n12133 6.998
R7563 VDD.n12038 VDD.n12037 6.998
R7564 VDD.n10901 VDD.n10900 6.998
R7565 VDD.n11080 VDD.n11079 6.998
R7566 VDD.n10866 VDD.n10865 6.998
R7567 VDD.n10694 VDD.n10693 6.998
R7568 VDD.n10693 VDD.n10692 6.998
R7569 VDD.n10902 VDD.n10901 6.998
R7570 VDD.n10867 VDD.n10866 6.998
R7571 VDD.n11079 VDD.n11078 6.998
R7572 VDD.n11671 VDD.n11670 6.998
R7573 VDD.n11585 VDD.n11584 6.998
R7574 VDD.n11670 VDD.n11669 6.998
R7575 VDD.n11584 VDD.n11583 6.998
R7576 VDD.n11365 VDD.n11364 6.998
R7577 VDD.n10810 VDD.n10809 6.981
R7578 VDD.n11625 VDD.n11624 6.981
R7579 VDD.n4633 VDD.n2771 6.774
R7580 VDD.n11187 VDD.n11186 6.687
R7581 VDD.n11948 VDD.n11947 6.687
R7582 VDD.n11951 VDD.n11950 6.687
R7583 VDD.n3117 VDD.n3116 6.686
R7584 VDD.n3355 VDD.n3354 6.686
R7585 VDD.n3592 VDD.n3591 6.686
R7586 VDD.n3830 VDD.n3829 6.686
R7587 VDD.n4067 VDD.n4066 6.686
R7588 VDD.n4305 VDD.n4304 6.686
R7589 VDD.n2987 VDD.n2986 6.643
R7590 VDD.n3011 VDD.n3010 6.643
R7591 VDD.n3225 VDD.n3224 6.643
R7592 VDD.n3248 VDD.n3247 6.643
R7593 VDD.n3462 VDD.n3461 6.643
R7594 VDD.n3486 VDD.n3485 6.643
R7595 VDD.n3628 VDD.n3627 6.643
R7596 VDD.n3700 VDD.n3699 6.643
R7597 VDD.n3723 VDD.n3722 6.643
R7598 VDD.n3792 VDD.n3791 6.643
R7599 VDD.n3937 VDD.n3936 6.643
R7600 VDD.n3961 VDD.n3960 6.643
R7601 VDD.n4175 VDD.n4174 6.643
R7602 VDD.n4198 VDD.n4197 6.643
R7603 VDD.n4412 VDD.n4411 6.643
R7604 VDD.n4436 VDD.n4435 6.643
R7605 VDD.n2042 VDD.n2041 6.643
R7606 VDD.n2056 VDD.n2055 6.643
R7607 VDD.n2273 VDD.n2272 6.643
R7608 VDD.n2287 VDD.n2286 6.643
R7609 VDD.n2512 VDD.n2511 6.643
R7610 VDD.n2582 VDD.n2581 6.643
R7611 VDD.n2737 VDD.n2736 6.643
R7612 VDD.n5115 VDD.n5114 6.643
R7613 VDD.n4891 VDD.n4890 6.643
R7614 VDD.n4877 VDD.n4876 6.643
R7615 VDD.n4660 VDD.n4659 6.643
R7616 VDD.n4646 VDD.n4645 6.643
R7617 VDD.n252 VDD.n251 6.643
R7618 VDD.n528 VDD.n527 6.643
R7619 VDD.n552 VDD.n551 6.643
R7620 VDD.n762 VDD.n761 6.643
R7621 VDD.n786 VDD.n785 6.643
R7622 VDD.n995 VDD.n994 6.643
R7623 VDD.n1019 VDD.n1018 6.643
R7624 VDD.n1229 VDD.n1228 6.643
R7625 VDD.n1253 VDD.n1252 6.643
R7626 VDD.n1462 VDD.n1461 6.643
R7627 VDD.n1486 VDD.n1485 6.643
R7628 VDD.n1502 VDD.n1499 6.643
R7629 VDD.n1696 VDD.n1695 6.643
R7630 VDD.n1720 VDD.n1719 6.643
R7631 VDD.n2014 VDD.n2013 6.643
R7632 VDD.n12087 VDD.n12085 6.593
R7633 VDD.n12087 VDD.n12086 6.593
R7634 VDD.n11020 VDD.n11018 6.593
R7635 VDD.n11020 VDD.n11019 6.593
R7636 VDD.n10728 VDD.n10726 6.593
R7637 VDD.n10728 VDD.n10727 6.593
R7638 VDD.n11787 VDD.n11784 6.593
R7639 VDD.n11787 VDD.n11786 6.593
R7640 VDD.n11499 VDD.n11496 6.593
R7641 VDD.n11499 VDD.n11498 6.593
R7642 VDD.n11318 VDD.n11316 6.593
R7643 VDD.n11318 VDD.n11317 6.593
R7644 VDD.n10341 VDD.n10220 6.452
R7645 VDD.n2831 VDD.n2830 6.413
R7646 VDD.n4479 VDD.n4478 6.413
R7647 VDD.n234 VDD.n233 6.413
R7648 VDD.n10767 VDD.n10765 6.4
R7649 VDD.n11537 VDD.n11535 6.4
R7650 VDD.n10103 VDD.n10102 6.389
R7651 VDD.n405 VDD.n401 6.206
R7652 VDD.n446 VDD.n442 6.206
R7653 VDD.n639 VDD.n635 6.206
R7654 VDD.n679 VDD.n675 6.206
R7655 VDD.n872 VDD.n868 6.206
R7656 VDD.n913 VDD.n909 6.206
R7657 VDD.n1106 VDD.n1102 6.206
R7658 VDD.n1146 VDD.n1142 6.206
R7659 VDD.n1339 VDD.n1335 6.206
R7660 VDD.n1380 VDD.n1376 6.206
R7661 VDD.n1573 VDD.n1569 6.206
R7662 VDD.n1613 VDD.n1609 6.206
R7663 VDD.n1806 VDD.n1802 6.206
R7664 VDD.n1847 VDD.n1843 6.206
R7665 VDD.n10921 VDD.n10920 6.206
R7666 VDD.n11720 VDD.n11719 6.206
R7667 VDD.n2793 VDD.n2791 6.068
R7668 VDD.n2988 VDD.n2984 6
R7669 VDD.n3012 VDD.n3008 6
R7670 VDD.n3226 VDD.n3222 6
R7671 VDD.n3249 VDD.n3245 6
R7672 VDD.n3463 VDD.n3459 6
R7673 VDD.n3487 VDD.n3483 6
R7674 VDD.n3701 VDD.n3697 6
R7675 VDD.n3724 VDD.n3720 6
R7676 VDD.n3938 VDD.n3934 6
R7677 VDD.n3962 VDD.n3958 6
R7678 VDD.n4176 VDD.n4172 6
R7679 VDD.n4199 VDD.n4195 6
R7680 VDD.n4413 VDD.n4409 6
R7681 VDD.n4437 VDD.n4433 6
R7682 VDD.n11131 VDD.n11130 5.92
R7683 VDD.n10341 VDD.n10340 5.721
R7684 VDD.n2137 VDD.n2136 5.538
R7685 VDD.n2186 VDD.n2185 5.538
R7686 VDD.n2368 VDD.n2367 5.538
R7687 VDD.n2417 VDD.n2416 5.538
R7688 VDD.n5196 VDD.n5195 5.538
R7689 VDD.n5263 VDD.n5262 5.538
R7690 VDD.n5021 VDD.n5020 5.538
R7691 VDD.n4972 VDD.n4971 5.538
R7692 VDD.n4790 VDD.n4789 5.538
R7693 VDD.n4741 VDD.n4740 5.538
R7694 VDD.n5481 VDD.n5480 5.458
R7695 VDD.n5842 VDD.n5841 5.458
R7696 VDD.n6204 VDD.n6203 5.458
R7697 VDD.n6566 VDD.n6565 5.458
R7698 VDD.n6928 VDD.n6927 5.458
R7699 VDD.n7290 VDD.n7289 5.458
R7700 VDD.n7652 VDD.n7651 5.458
R7701 VDD.n8014 VDD.n8013 5.458
R7702 VDD.n8376 VDD.n8375 5.458
R7703 VDD.n8738 VDD.n8737 5.458
R7704 VDD.n9100 VDD.n9099 5.458
R7705 VDD.n9462 VDD.n9461 5.458
R7706 VDD.n9824 VDD.n9823 5.458
R7707 VDD.n80 VDD.n78 5.454
R7708 VDD.n46 VDD.n44 5.454
R7709 VDD.n11403 VDD.n11402 5.454
R7710 VDD.n11205 VDD.n11203 5.454
R7711 VDD.n11892 VDD.n11891 5.454
R7712 VDD.n12311 VDD.n12309 5.454
R7713 VDD.n12277 VDD.n12275 5.454
R7714 VDD.n5231 VDD.n5230 5.415
R7715 VDD.n11354 VDD.n11353 5.299
R7716 VDD.n11683 VDD.n11682 5.299
R7717 VDD.n11631 VDD.n11630 5.299
R7718 VDD.n11682 VDD.n11681 5.299
R7719 VDD.n11630 VDD.n11629 5.299
R7720 VDD.n11353 VDD.n11352 5.299
R7721 VDD.n5524 VDD.n5523 5.081
R7722 VDD.n5885 VDD.n5884 5.081
R7723 VDD.n6247 VDD.n6246 5.081
R7724 VDD.n6609 VDD.n6608 5.081
R7725 VDD.n6971 VDD.n6970 5.081
R7726 VDD.n7333 VDD.n7332 5.081
R7727 VDD.n7695 VDD.n7694 5.081
R7728 VDD.n8057 VDD.n8056 5.081
R7729 VDD.n8419 VDD.n8418 5.081
R7730 VDD.n8781 VDD.n8780 5.081
R7731 VDD.n9143 VDD.n9142 5.081
R7732 VDD.n9505 VDD.n9504 5.081
R7733 VDD.n9867 VDD.n9866 5.081
R7734 VDD.n11434 VDD.n11433 5.052
R7735 VDD.n11236 VDD.n11235 5.052
R7736 VDD.n12172 VDD.n12171 5.052
R7737 VDD.n11968 VDD.n11967 5.052
R7738 VDD.n12206 VDD.n12205 5.052
R7739 VDD.n12002 VDD.n12001 5.052
R7740 VDD.n11111 VDD.n11110 5.052
R7741 VDD.n11162 VDD.n11161 5.052
R7742 VDD.n11920 VDD.n11919 5.052
R7743 VDD.n2021 VDD.n2020 4.818
R7744 VDD.n4498 VDD.n4497 4.731
R7745 VDD.n2856 VDD.n2855 4.731
R7746 VDD.n202 VDD.n201 4.698
R7747 VDD.n2794 VDD.n2793 4.65
R7748 VDD.n3118 VDD.n3117 4.65
R7749 VDD.n3356 VDD.n3355 4.65
R7750 VDD.n3593 VDD.n3592 4.65
R7751 VDD.n3831 VDD.n3830 4.65
R7752 VDD.n4068 VDD.n4067 4.65
R7753 VDD.n4306 VDD.n4305 4.65
R7754 VDD.n542 VDD.n541 4.65
R7755 VDD.n776 VDD.n775 4.65
R7756 VDD.n1009 VDD.n1008 4.65
R7757 VDD.n1243 VDD.n1242 4.65
R7758 VDD.n1476 VDD.n1475 4.65
R7759 VDD.n1710 VDD.n1709 4.65
R7760 VDD.n225 VDD.n224 4.65
R7761 VDD.n215 VDD.n214 4.65
R7762 VDD.n256 VDD.n255 4.65
R7763 VDD.n279 VDD.n278 4.65
R7764 VDD.n310 VDD.n309 4.65
R7765 VDD.n328 VDD.n327 4.65
R7766 VDD.n379 VDD.n378 4.65
R7767 VDD.n393 VDD.n392 4.65
R7768 VDD.n407 VDD.n406 4.65
R7769 VDD.n422 VDD.n421 4.65
R7770 VDD.n434 VDD.n433 4.65
R7771 VDD.n448 VDD.n447 4.65
R7772 VDD.n462 VDD.n461 4.65
R7773 VDD.n476 VDD.n475 4.65
R7774 VDD.n490 VDD.n489 4.65
R7775 VDD.n504 VDD.n503 4.65
R7776 VDD.n518 VDD.n517 4.65
R7777 VDD.n532 VDD.n531 4.65
R7778 VDD.n556 VDD.n555 4.65
R7779 VDD.n571 VDD.n570 4.65
R7780 VDD.n585 VDD.n584 4.65
R7781 VDD.n599 VDD.n598 4.65
R7782 VDD.n613 VDD.n612 4.65
R7783 VDD.n627 VDD.n626 4.65
R7784 VDD.n641 VDD.n640 4.65
R7785 VDD.n655 VDD.n654 4.65
R7786 VDD.n667 VDD.n666 4.65
R7787 VDD.n681 VDD.n680 4.65
R7788 VDD.n695 VDD.n694 4.65
R7789 VDD.n709 VDD.n708 4.65
R7790 VDD.n723 VDD.n722 4.65
R7791 VDD.n738 VDD.n737 4.65
R7792 VDD.n752 VDD.n751 4.65
R7793 VDD.n766 VDD.n765 4.65
R7794 VDD.n790 VDD.n789 4.65
R7795 VDD.n804 VDD.n803 4.65
R7796 VDD.n818 VDD.n817 4.65
R7797 VDD.n832 VDD.n831 4.65
R7798 VDD.n846 VDD.n845 4.65
R7799 VDD.n860 VDD.n859 4.65
R7800 VDD.n874 VDD.n873 4.65
R7801 VDD.n889 VDD.n888 4.65
R7802 VDD.n901 VDD.n900 4.65
R7803 VDD.n915 VDD.n914 4.65
R7804 VDD.n929 VDD.n928 4.65
R7805 VDD.n943 VDD.n942 4.65
R7806 VDD.n957 VDD.n956 4.65
R7807 VDD.n971 VDD.n970 4.65
R7808 VDD.n985 VDD.n984 4.65
R7809 VDD.n999 VDD.n998 4.65
R7810 VDD.n1023 VDD.n1022 4.65
R7811 VDD.n1038 VDD.n1037 4.65
R7812 VDD.n1052 VDD.n1051 4.65
R7813 VDD.n1066 VDD.n1065 4.65
R7814 VDD.n1080 VDD.n1079 4.65
R7815 VDD.n1094 VDD.n1093 4.65
R7816 VDD.n1108 VDD.n1107 4.65
R7817 VDD.n1122 VDD.n1121 4.65
R7818 VDD.n1134 VDD.n1133 4.65
R7819 VDD.n1148 VDD.n1147 4.65
R7820 VDD.n1162 VDD.n1161 4.65
R7821 VDD.n1176 VDD.n1175 4.65
R7822 VDD.n1190 VDD.n1189 4.65
R7823 VDD.n1205 VDD.n1204 4.65
R7824 VDD.n1219 VDD.n1218 4.65
R7825 VDD.n1233 VDD.n1232 4.65
R7826 VDD.n1257 VDD.n1256 4.65
R7827 VDD.n1271 VDD.n1270 4.65
R7828 VDD.n1285 VDD.n1284 4.65
R7829 VDD.n1299 VDD.n1298 4.65
R7830 VDD.n1313 VDD.n1312 4.65
R7831 VDD.n1327 VDD.n1326 4.65
R7832 VDD.n1341 VDD.n1340 4.65
R7833 VDD.n1356 VDD.n1355 4.65
R7834 VDD.n1368 VDD.n1367 4.65
R7835 VDD.n1382 VDD.n1381 4.65
R7836 VDD.n1396 VDD.n1395 4.65
R7837 VDD.n1410 VDD.n1409 4.65
R7838 VDD.n1424 VDD.n1423 4.65
R7839 VDD.n1438 VDD.n1437 4.65
R7840 VDD.n1452 VDD.n1451 4.65
R7841 VDD.n1466 VDD.n1465 4.65
R7842 VDD.n1490 VDD.n1489 4.65
R7843 VDD.n1505 VDD.n1504 4.65
R7844 VDD.n1519 VDD.n1518 4.65
R7845 VDD.n1533 VDD.n1532 4.65
R7846 VDD.n1547 VDD.n1546 4.65
R7847 VDD.n1561 VDD.n1560 4.65
R7848 VDD.n1575 VDD.n1574 4.65
R7849 VDD.n1589 VDD.n1588 4.65
R7850 VDD.n1601 VDD.n1600 4.65
R7851 VDD.n1615 VDD.n1614 4.65
R7852 VDD.n1629 VDD.n1628 4.65
R7853 VDD.n1643 VDD.n1642 4.65
R7854 VDD.n1657 VDD.n1656 4.65
R7855 VDD.n1672 VDD.n1671 4.65
R7856 VDD.n1686 VDD.n1685 4.65
R7857 VDD.n1700 VDD.n1699 4.65
R7858 VDD.n1724 VDD.n1723 4.65
R7859 VDD.n1738 VDD.n1737 4.65
R7860 VDD.n1752 VDD.n1751 4.65
R7861 VDD.n1766 VDD.n1765 4.65
R7862 VDD.n1780 VDD.n1779 4.65
R7863 VDD.n1794 VDD.n1793 4.65
R7864 VDD.n1808 VDD.n1807 4.65
R7865 VDD.n1823 VDD.n1822 4.65
R7866 VDD.n1835 VDD.n1834 4.65
R7867 VDD.n1849 VDD.n1848 4.65
R7868 VDD.n1885 VDD.n1884 4.65
R7869 VDD.n1904 VDD.n1903 4.65
R7870 VDD.n1923 VDD.n1922 4.65
R7871 VDD.n1867 VDD.n1866 4.65
R7872 VDD.n1945 VDD.n1944 4.65
R7873 VDD.n2018 VDD.n2017 4.65
R7874 VDD.n2976 VDD.n2975 4.65
R7875 VDD.n2990 VDD.n2989 4.65
R7876 VDD.n3002 VDD.n3001 4.65
R7877 VDD.n3129 VDD.n3128 4.65
R7878 VDD.n3143 VDD.n3142 4.65
R7879 VDD.n3158 VDD.n3157 4.65
R7880 VDD.n3172 VDD.n3171 4.65
R7881 VDD.n3186 VDD.n3185 4.65
R7882 VDD.n3200 VDD.n3199 4.65
R7883 VDD.n3214 VDD.n3213 4.65
R7884 VDD.n3228 VDD.n3227 4.65
R7885 VDD.n3239 VDD.n3238 4.65
R7886 VDD.n3367 VDD.n3366 4.65
R7887 VDD.n3381 VDD.n3380 4.65
R7888 VDD.n3395 VDD.n3394 4.65
R7889 VDD.n3409 VDD.n3408 4.65
R7890 VDD.n3423 VDD.n3422 4.65
R7891 VDD.n3437 VDD.n3436 4.65
R7892 VDD.n3451 VDD.n3450 4.65
R7893 VDD.n3465 VDD.n3464 4.65
R7894 VDD.n3477 VDD.n3476 4.65
R7895 VDD.n3604 VDD.n3603 4.65
R7896 VDD.n3618 VDD.n3617 4.65
R7897 VDD.n3633 VDD.n3632 4.65
R7898 VDD.n3647 VDD.n3646 4.65
R7899 VDD.n3661 VDD.n3660 4.65
R7900 VDD.n3675 VDD.n3674 4.65
R7901 VDD.n3689 VDD.n3688 4.65
R7902 VDD.n3703 VDD.n3702 4.65
R7903 VDD.n3714 VDD.n3713 4.65
R7904 VDD.n3842 VDD.n3841 4.65
R7905 VDD.n3856 VDD.n3855 4.65
R7906 VDD.n3870 VDD.n3869 4.65
R7907 VDD.n3884 VDD.n3883 4.65
R7908 VDD.n3898 VDD.n3897 4.65
R7909 VDD.n3912 VDD.n3911 4.65
R7910 VDD.n3926 VDD.n3925 4.65
R7911 VDD.n3940 VDD.n3939 4.65
R7912 VDD.n3952 VDD.n3951 4.65
R7913 VDD.n4079 VDD.n4078 4.65
R7914 VDD.n4093 VDD.n4092 4.65
R7915 VDD.n4108 VDD.n4107 4.65
R7916 VDD.n4122 VDD.n4121 4.65
R7917 VDD.n4136 VDD.n4135 4.65
R7918 VDD.n4150 VDD.n4149 4.65
R7919 VDD.n4164 VDD.n4163 4.65
R7920 VDD.n4178 VDD.n4177 4.65
R7921 VDD.n4189 VDD.n4188 4.65
R7922 VDD.n4317 VDD.n4316 4.65
R7923 VDD.n4331 VDD.n4330 4.65
R7924 VDD.n4345 VDD.n4344 4.65
R7925 VDD.n4359 VDD.n4358 4.65
R7926 VDD.n4373 VDD.n4372 4.65
R7927 VDD.n4387 VDD.n4386 4.65
R7928 VDD.n4401 VDD.n4400 4.65
R7929 VDD.n4415 VDD.n4414 4.65
R7930 VDD.n4427 VDD.n4426 4.65
R7931 VDD.n4560 VDD.n4559 4.65
R7932 VDD.n4512 VDD.n4511 4.65
R7933 VDD.n2962 VDD.n2961 4.65
R7934 VDD.n2915 VDD.n2914 4.65
R7935 VDD.n2896 VDD.n2895 4.65
R7936 VDD.n2866 VDD.n2865 4.65
R7937 VDD.n2840 VDD.n2839 4.65
R7938 VDD.n2808 VDD.n2807 4.65
R7939 VDD.n2787 VDD.n2786 4.65
R7940 VDD.n3014 VDD.n3013 4.65
R7941 VDD.n3028 VDD.n3027 4.65
R7942 VDD.n3042 VDD.n3041 4.65
R7943 VDD.n3056 VDD.n3055 4.65
R7944 VDD.n3070 VDD.n3069 4.65
R7945 VDD.n3084 VDD.n3083 4.65
R7946 VDD.n3098 VDD.n3097 4.65
R7947 VDD.n3112 VDD.n3111 4.65
R7948 VDD.n3251 VDD.n3250 4.65
R7949 VDD.n3265 VDD.n3264 4.65
R7950 VDD.n3279 VDD.n3278 4.65
R7951 VDD.n3293 VDD.n3292 4.65
R7952 VDD.n3307 VDD.n3306 4.65
R7953 VDD.n3322 VDD.n3321 4.65
R7954 VDD.n3336 VDD.n3335 4.65
R7955 VDD.n3350 VDD.n3349 4.65
R7956 VDD.n3489 VDD.n3488 4.65
R7957 VDD.n3503 VDD.n3502 4.65
R7958 VDD.n3517 VDD.n3516 4.65
R7959 VDD.n3531 VDD.n3530 4.65
R7960 VDD.n3545 VDD.n3544 4.65
R7961 VDD.n3559 VDD.n3558 4.65
R7962 VDD.n3573 VDD.n3572 4.65
R7963 VDD.n3587 VDD.n3586 4.65
R7964 VDD.n3726 VDD.n3725 4.65
R7965 VDD.n3740 VDD.n3739 4.65
R7966 VDD.n3754 VDD.n3753 4.65
R7967 VDD.n3768 VDD.n3767 4.65
R7968 VDD.n3782 VDD.n3781 4.65
R7969 VDD.n3797 VDD.n3796 4.65
R7970 VDD.n3811 VDD.n3810 4.65
R7971 VDD.n3825 VDD.n3824 4.65
R7972 VDD.n3964 VDD.n3963 4.65
R7973 VDD.n3978 VDD.n3977 4.65
R7974 VDD.n3992 VDD.n3991 4.65
R7975 VDD.n4006 VDD.n4005 4.65
R7976 VDD.n4020 VDD.n4019 4.65
R7977 VDD.n4034 VDD.n4033 4.65
R7978 VDD.n4048 VDD.n4047 4.65
R7979 VDD.n4062 VDD.n4061 4.65
R7980 VDD.n4201 VDD.n4200 4.65
R7981 VDD.n4215 VDD.n4214 4.65
R7982 VDD.n4229 VDD.n4228 4.65
R7983 VDD.n4243 VDD.n4242 4.65
R7984 VDD.n4257 VDD.n4256 4.65
R7985 VDD.n4272 VDD.n4271 4.65
R7986 VDD.n4286 VDD.n4285 4.65
R7987 VDD.n4300 VDD.n4299 4.65
R7988 VDD.n4439 VDD.n4438 4.65
R7989 VDD.n4453 VDD.n4452 4.65
R7990 VDD.n4472 VDD.n4471 4.65
R7991 VDD.n4492 VDD.n4491 4.65
R7992 VDD.n4532 VDD.n4531 4.65
R7993 VDD.n4623 VDD.n4622 4.65
R7994 VDD.n4884 VDD.n4883 4.65
R7995 VDD.n4653 VDD.n4652 4.65
R7996 VDD.n2049 VDD.n2048 4.65
R7997 VDD.n2280 VDD.n2279 4.65
R7998 VDD.n5633 VDD.n5632 4.65
R7999 VDD.n5601 VDD.n5600 4.65
R8000 VDD.n5994 VDD.n5993 4.65
R8001 VDD.n5962 VDD.n5961 4.65
R8002 VDD.n6356 VDD.n6355 4.65
R8003 VDD.n6324 VDD.n6323 4.65
R8004 VDD.n6718 VDD.n6717 4.65
R8005 VDD.n6686 VDD.n6685 4.65
R8006 VDD.n7080 VDD.n7079 4.65
R8007 VDD.n7048 VDD.n7047 4.65
R8008 VDD.n7442 VDD.n7441 4.65
R8009 VDD.n7410 VDD.n7409 4.65
R8010 VDD.n7804 VDD.n7803 4.65
R8011 VDD.n7772 VDD.n7771 4.65
R8012 VDD.n8166 VDD.n8165 4.65
R8013 VDD.n8134 VDD.n8133 4.65
R8014 VDD.n8528 VDD.n8527 4.65
R8015 VDD.n8496 VDD.n8495 4.65
R8016 VDD.n8890 VDD.n8889 4.65
R8017 VDD.n8858 VDD.n8857 4.65
R8018 VDD.n9252 VDD.n9251 4.65
R8019 VDD.n9220 VDD.n9219 4.65
R8020 VDD.n9614 VDD.n9613 4.65
R8021 VDD.n9582 VDD.n9581 4.65
R8022 VDD.n9976 VDD.n9975 4.65
R8023 VDD.n9944 VDD.n9943 4.65
R8024 VDD.n10289 VDD.n10288 4.65
R8025 VDD.n10171 VDD.n10170 4.65
R8026 VDD.n10088 VDD.n10087 4.65
R8027 VDD.n10044 VDD.n10043 4.65
R8028 VDD.n10636 VDD.n10635 4.65
R8029 VDD.n10517 VDD.n10516 4.65
R8030 VDD.n11118 VDD.n11117 4.65
R8031 VDD.n10853 VDD.n10852 4.65
R8032 VDD.n10943 VDD.n10942 4.65
R8033 VDD.n11882 VDD.n11881 4.65
R8034 VDD.n11700 VDD.n11699 4.65
R8035 VDD.n11634 VDD.n11633 4.65
R8036 VDD.n12088 VDD.n12087 4.65
R8037 VDD.n11319 VDD.n11318 4.65
R8038 VDD.n2021 VDD.n202 4.533
R8039 VDD.n541 VDD.n537 4.533
R8040 VDD.n541 VDD.n540 4.533
R8041 VDD.n775 VDD.n771 4.533
R8042 VDD.n775 VDD.n774 4.533
R8043 VDD.n1008 VDD.n1004 4.533
R8044 VDD.n1008 VDD.n1007 4.533
R8045 VDD.n1242 VDD.n1238 4.533
R8046 VDD.n1242 VDD.n1241 4.533
R8047 VDD.n1475 VDD.n1471 4.533
R8048 VDD.n1475 VDD.n1474 4.533
R8049 VDD.n1709 VDD.n1705 4.533
R8050 VDD.n1709 VDD.n1708 4.533
R8051 VDD.n11698 VDD.n11697 4.523
R8052 VDD.n11600 VDD.n11599 4.523
R8053 VDD.n2825 VDD.n2824 4.5
R8054 VDD.n2850 VDD.n2849 4.5
R8055 VDD.n2881 VDD.n2880 4.5
R8056 VDD.n2951 VDD.n2950 4.5
R8057 VDD.n4622 VDD.n4615 4.5
R8058 VDD.n2010 VDD.n2009 4.5
R8059 VDD.n368 VDD.n367 4.5
R8060 VDD.n265 VDD.n264 4.5
R8061 VDD.n255 VDD.n248 4.5
R8062 VDD.n296 VDD.n295 4.5
R8063 VDD.n2496 VDD.n2495 4.5
R8064 VDD.n2723 VDD.n2722 4.5
R8065 VDD.n2688 VDD.n2687 4.5
R8066 VDD.n2645 VDD.n2644 4.5
R8067 VDD.n5249 VDD.n5248 4.5
R8068 VDD.n5270 VDD.n5269 4.5
R8069 VDD.n5289 VDD.n5288 4.5
R8070 VDD.n5232 VDD.n5231 4.5
R8071 VDD.n5294 VDD.n5293 4.5
R8072 VDD.n5224 VDD.n5223 4.5
R8073 VDD.n5205 VDD.n5204 4.5
R8074 VDD.n5184 VDD.n5183 4.5
R8075 VDD.n5165 VDD.n5164 4.5
R8076 VDD.n149 VDD.n148 4.5
R8077 VDD.n130 VDD.n129 4.5
R8078 VDD.n2563 VDD.n2562 4.5
R8079 VDD.n2574 VDD.n2573 4.5
R8080 VDD.n2542 VDD.n2541 4.5
R8081 VDD.n2587 VDD.n2586 4.5
R8082 VDD.n2526 VDD.n2524 4.5
R8083 VDD.n2516 VDD.n2515 4.5
R8084 VDD.n2669 VDD.n2668 4.5
R8085 VDD.n2741 VDD.n2740 4.5
R8086 VDD.n2747 VDD.n2746 4.5
R8087 VDD.n2752 VDD.n2751 4.5
R8088 VDD.n2764 VDD.n2763 4.5
R8089 VDD.n5120 VDD.n5119 4.5
R8090 VDD.n5100 VDD.n5099 4.5
R8091 VDD.n5648 VDD.n5647 4.5
R8092 VDD.n5629 VDD.n5628 4.5
R8093 VDD.n5621 VDD.n5620 4.5
R8094 VDD.n5607 VDD.n5606 4.5
R8095 VDD.n5528 VDD.n5516 4.5
R8096 VDD.n5508 VDD.n5507 4.5
R8097 VDD.n5498 VDD.n5497 4.5
R8098 VDD.n5488 VDD.n5487 4.5
R8099 VDD.n5476 VDD.n5475 4.5
R8100 VDD.n5359 VDD.n5325 4.5
R8101 VDD.n5352 VDD.n5328 4.5
R8102 VDD.n5367 VDD.n5322 4.5
R8103 VDD.n5376 VDD.n5319 4.5
R8104 VDD.n5346 VDD.n5331 4.5
R8105 VDD.n5343 VDD.n5335 4.5
R8106 VDD.n5339 VDD.n5338 4.5
R8107 VDD.n5615 VDD.n5614 4.5
R8108 VDD.n5659 VDD.n5658 4.5
R8109 VDD.n6009 VDD.n6008 4.5
R8110 VDD.n5990 VDD.n5989 4.5
R8111 VDD.n5982 VDD.n5981 4.5
R8112 VDD.n5968 VDD.n5967 4.5
R8113 VDD.n5889 VDD.n5877 4.5
R8114 VDD.n5869 VDD.n5868 4.5
R8115 VDD.n5859 VDD.n5858 4.5
R8116 VDD.n5849 VDD.n5848 4.5
R8117 VDD.n5837 VDD.n5836 4.5
R8118 VDD.n5720 VDD.n5686 4.5
R8119 VDD.n5713 VDD.n5689 4.5
R8120 VDD.n5728 VDD.n5683 4.5
R8121 VDD.n5737 VDD.n5680 4.5
R8122 VDD.n5707 VDD.n5692 4.5
R8123 VDD.n5704 VDD.n5696 4.5
R8124 VDD.n5700 VDD.n5699 4.5
R8125 VDD.n5976 VDD.n5975 4.5
R8126 VDD.n6020 VDD.n6019 4.5
R8127 VDD.n6371 VDD.n6370 4.5
R8128 VDD.n6352 VDD.n6351 4.5
R8129 VDD.n6344 VDD.n6343 4.5
R8130 VDD.n6330 VDD.n6329 4.5
R8131 VDD.n6251 VDD.n6239 4.5
R8132 VDD.n6231 VDD.n6230 4.5
R8133 VDD.n6221 VDD.n6220 4.5
R8134 VDD.n6211 VDD.n6210 4.5
R8135 VDD.n6199 VDD.n6198 4.5
R8136 VDD.n6082 VDD.n6048 4.5
R8137 VDD.n6075 VDD.n6051 4.5
R8138 VDD.n6090 VDD.n6045 4.5
R8139 VDD.n6099 VDD.n6042 4.5
R8140 VDD.n6069 VDD.n6054 4.5
R8141 VDD.n6066 VDD.n6058 4.5
R8142 VDD.n6062 VDD.n6061 4.5
R8143 VDD.n6338 VDD.n6337 4.5
R8144 VDD.n6382 VDD.n6381 4.5
R8145 VDD.n6733 VDD.n6732 4.5
R8146 VDD.n6714 VDD.n6713 4.5
R8147 VDD.n6706 VDD.n6705 4.5
R8148 VDD.n6692 VDD.n6691 4.5
R8149 VDD.n6613 VDD.n6601 4.5
R8150 VDD.n6593 VDD.n6592 4.5
R8151 VDD.n6583 VDD.n6582 4.5
R8152 VDD.n6573 VDD.n6572 4.5
R8153 VDD.n6561 VDD.n6560 4.5
R8154 VDD.n6444 VDD.n6410 4.5
R8155 VDD.n6437 VDD.n6413 4.5
R8156 VDD.n6452 VDD.n6407 4.5
R8157 VDD.n6461 VDD.n6404 4.5
R8158 VDD.n6431 VDD.n6416 4.5
R8159 VDD.n6428 VDD.n6420 4.5
R8160 VDD.n6424 VDD.n6423 4.5
R8161 VDD.n6700 VDD.n6699 4.5
R8162 VDD.n6744 VDD.n6743 4.5
R8163 VDD.n7095 VDD.n7094 4.5
R8164 VDD.n7076 VDD.n7075 4.5
R8165 VDD.n7068 VDD.n7067 4.5
R8166 VDD.n7054 VDD.n7053 4.5
R8167 VDD.n6975 VDD.n6963 4.5
R8168 VDD.n6955 VDD.n6954 4.5
R8169 VDD.n6945 VDD.n6944 4.5
R8170 VDD.n6935 VDD.n6934 4.5
R8171 VDD.n6923 VDD.n6922 4.5
R8172 VDD.n6806 VDD.n6772 4.5
R8173 VDD.n6799 VDD.n6775 4.5
R8174 VDD.n6814 VDD.n6769 4.5
R8175 VDD.n6823 VDD.n6766 4.5
R8176 VDD.n6793 VDD.n6778 4.5
R8177 VDD.n6790 VDD.n6782 4.5
R8178 VDD.n6786 VDD.n6785 4.5
R8179 VDD.n7062 VDD.n7061 4.5
R8180 VDD.n7106 VDD.n7105 4.5
R8181 VDD.n7457 VDD.n7456 4.5
R8182 VDD.n7438 VDD.n7437 4.5
R8183 VDD.n7430 VDD.n7429 4.5
R8184 VDD.n7416 VDD.n7415 4.5
R8185 VDD.n7337 VDD.n7325 4.5
R8186 VDD.n7317 VDD.n7316 4.5
R8187 VDD.n7307 VDD.n7306 4.5
R8188 VDD.n7297 VDD.n7296 4.5
R8189 VDD.n7285 VDD.n7284 4.5
R8190 VDD.n7168 VDD.n7134 4.5
R8191 VDD.n7161 VDD.n7137 4.5
R8192 VDD.n7176 VDD.n7131 4.5
R8193 VDD.n7185 VDD.n7128 4.5
R8194 VDD.n7155 VDD.n7140 4.5
R8195 VDD.n7152 VDD.n7144 4.5
R8196 VDD.n7148 VDD.n7147 4.5
R8197 VDD.n7424 VDD.n7423 4.5
R8198 VDD.n7468 VDD.n7467 4.5
R8199 VDD.n7819 VDD.n7818 4.5
R8200 VDD.n7800 VDD.n7799 4.5
R8201 VDD.n7792 VDD.n7791 4.5
R8202 VDD.n7778 VDD.n7777 4.5
R8203 VDD.n7699 VDD.n7687 4.5
R8204 VDD.n7679 VDD.n7678 4.5
R8205 VDD.n7669 VDD.n7668 4.5
R8206 VDD.n7659 VDD.n7658 4.5
R8207 VDD.n7647 VDD.n7646 4.5
R8208 VDD.n7530 VDD.n7496 4.5
R8209 VDD.n7523 VDD.n7499 4.5
R8210 VDD.n7538 VDD.n7493 4.5
R8211 VDD.n7547 VDD.n7490 4.5
R8212 VDD.n7517 VDD.n7502 4.5
R8213 VDD.n7514 VDD.n7506 4.5
R8214 VDD.n7510 VDD.n7509 4.5
R8215 VDD.n7786 VDD.n7785 4.5
R8216 VDD.n7830 VDD.n7829 4.5
R8217 VDD.n8181 VDD.n8180 4.5
R8218 VDD.n8162 VDD.n8161 4.5
R8219 VDD.n8154 VDD.n8153 4.5
R8220 VDD.n8140 VDD.n8139 4.5
R8221 VDD.n8061 VDD.n8049 4.5
R8222 VDD.n8041 VDD.n8040 4.5
R8223 VDD.n8031 VDD.n8030 4.5
R8224 VDD.n8021 VDD.n8020 4.5
R8225 VDD.n8009 VDD.n8008 4.5
R8226 VDD.n7892 VDD.n7858 4.5
R8227 VDD.n7885 VDD.n7861 4.5
R8228 VDD.n7900 VDD.n7855 4.5
R8229 VDD.n7909 VDD.n7852 4.5
R8230 VDD.n7879 VDD.n7864 4.5
R8231 VDD.n7876 VDD.n7868 4.5
R8232 VDD.n7872 VDD.n7871 4.5
R8233 VDD.n8148 VDD.n8147 4.5
R8234 VDD.n8192 VDD.n8191 4.5
R8235 VDD.n8543 VDD.n8542 4.5
R8236 VDD.n8524 VDD.n8523 4.5
R8237 VDD.n8516 VDD.n8515 4.5
R8238 VDD.n8502 VDD.n8501 4.5
R8239 VDD.n8423 VDD.n8411 4.5
R8240 VDD.n8403 VDD.n8402 4.5
R8241 VDD.n8393 VDD.n8392 4.5
R8242 VDD.n8383 VDD.n8382 4.5
R8243 VDD.n8371 VDD.n8370 4.5
R8244 VDD.n8254 VDD.n8220 4.5
R8245 VDD.n8247 VDD.n8223 4.5
R8246 VDD.n8262 VDD.n8217 4.5
R8247 VDD.n8271 VDD.n8214 4.5
R8248 VDD.n8241 VDD.n8226 4.5
R8249 VDD.n8238 VDD.n8230 4.5
R8250 VDD.n8234 VDD.n8233 4.5
R8251 VDD.n8510 VDD.n8509 4.5
R8252 VDD.n8554 VDD.n8553 4.5
R8253 VDD.n8905 VDD.n8904 4.5
R8254 VDD.n8886 VDD.n8885 4.5
R8255 VDD.n8878 VDD.n8877 4.5
R8256 VDD.n8864 VDD.n8863 4.5
R8257 VDD.n8785 VDD.n8773 4.5
R8258 VDD.n8765 VDD.n8764 4.5
R8259 VDD.n8755 VDD.n8754 4.5
R8260 VDD.n8745 VDD.n8744 4.5
R8261 VDD.n8733 VDD.n8732 4.5
R8262 VDD.n8616 VDD.n8582 4.5
R8263 VDD.n8609 VDD.n8585 4.5
R8264 VDD.n8624 VDD.n8579 4.5
R8265 VDD.n8633 VDD.n8576 4.5
R8266 VDD.n8603 VDD.n8588 4.5
R8267 VDD.n8600 VDD.n8592 4.5
R8268 VDD.n8596 VDD.n8595 4.5
R8269 VDD.n8872 VDD.n8871 4.5
R8270 VDD.n8916 VDD.n8915 4.5
R8271 VDD.n9267 VDD.n9266 4.5
R8272 VDD.n9248 VDD.n9247 4.5
R8273 VDD.n9240 VDD.n9239 4.5
R8274 VDD.n9226 VDD.n9225 4.5
R8275 VDD.n9147 VDD.n9135 4.5
R8276 VDD.n9127 VDD.n9126 4.5
R8277 VDD.n9117 VDD.n9116 4.5
R8278 VDD.n9107 VDD.n9106 4.5
R8279 VDD.n9095 VDD.n9094 4.5
R8280 VDD.n8978 VDD.n8944 4.5
R8281 VDD.n8971 VDD.n8947 4.5
R8282 VDD.n8986 VDD.n8941 4.5
R8283 VDD.n8995 VDD.n8938 4.5
R8284 VDD.n8965 VDD.n8950 4.5
R8285 VDD.n8962 VDD.n8954 4.5
R8286 VDD.n8958 VDD.n8957 4.5
R8287 VDD.n9234 VDD.n9233 4.5
R8288 VDD.n9278 VDD.n9277 4.5
R8289 VDD.n9629 VDD.n9628 4.5
R8290 VDD.n9610 VDD.n9609 4.5
R8291 VDD.n9602 VDD.n9601 4.5
R8292 VDD.n9588 VDD.n9587 4.5
R8293 VDD.n9509 VDD.n9497 4.5
R8294 VDD.n9489 VDD.n9488 4.5
R8295 VDD.n9479 VDD.n9478 4.5
R8296 VDD.n9469 VDD.n9468 4.5
R8297 VDD.n9457 VDD.n9456 4.5
R8298 VDD.n9340 VDD.n9306 4.5
R8299 VDD.n9333 VDD.n9309 4.5
R8300 VDD.n9348 VDD.n9303 4.5
R8301 VDD.n9357 VDD.n9300 4.5
R8302 VDD.n9327 VDD.n9312 4.5
R8303 VDD.n9324 VDD.n9316 4.5
R8304 VDD.n9320 VDD.n9319 4.5
R8305 VDD.n9596 VDD.n9595 4.5
R8306 VDD.n9640 VDD.n9639 4.5
R8307 VDD.n9991 VDD.n9990 4.5
R8308 VDD.n9972 VDD.n9971 4.5
R8309 VDD.n9964 VDD.n9963 4.5
R8310 VDD.n9950 VDD.n9949 4.5
R8311 VDD.n9871 VDD.n9859 4.5
R8312 VDD.n9851 VDD.n9850 4.5
R8313 VDD.n9841 VDD.n9840 4.5
R8314 VDD.n9831 VDD.n9830 4.5
R8315 VDD.n9819 VDD.n9818 4.5
R8316 VDD.n9702 VDD.n9668 4.5
R8317 VDD.n9695 VDD.n9671 4.5
R8318 VDD.n9710 VDD.n9665 4.5
R8319 VDD.n9719 VDD.n9662 4.5
R8320 VDD.n9689 VDD.n9674 4.5
R8321 VDD.n9686 VDD.n9678 4.5
R8322 VDD.n9682 VDD.n9681 4.5
R8323 VDD.n9958 VDD.n9957 4.5
R8324 VDD.n10002 VDD.n10001 4.5
R8325 VDD.n10759 VDD.n10758 4.5
R8326 VDD.n10768 VDD.n10767 4.5
R8327 VDD.n10872 VDD.n10871 4.5
R8328 VDD.n10858 VDD.n10857 4.5
R8329 VDD.n11101 VDD.n11099 4.5
R8330 VDD.n11105 VDD.n11096 4.5
R8331 VDD.n11087 VDD.n11086 4.5
R8332 VDD.n11014 VDD.n10984 4.5
R8333 VDD.n11073 VDD.n11016 4.5
R8334 VDD.n11069 VDD.n11068 4.5
R8335 VDD.n11053 VDD.n11052 4.5
R8336 VDD.n10909 VDD.n10908 4.5
R8337 VDD.n10952 VDD.n10921 4.5
R8338 VDD.n10946 VDD.n10931 4.5
R8339 VDD.n11036 VDD.n11035 4.5
R8340 VDD.n10956 VDD.n10918 4.5
R8341 VDD.n11010 VDD.n11009 4.5
R8342 VDD.n10997 VDD.n10995 4.5
R8343 VDD.n11166 VDD.n11165 4.5
R8344 VDD.n11180 VDD.n11179 4.5
R8345 VDD.n11152 VDD.n11151 4.5
R8346 VDD.n11138 VDD.n11116 4.5
R8347 VDD.n10840 VDD.n10839 4.5
R8348 VDD.n10824 VDD.n10819 4.5
R8349 VDD.n10744 VDD.n10743 4.5
R8350 VDD.n10781 VDD.n10780 4.5
R8351 VDD.n10724 VDD.n10700 4.5
R8352 VDD.n11538 VDD.n11537 4.5
R8353 VDD.n11529 VDD.n11528 4.5
R8354 VDD.n11721 VDD.n11720 4.5
R8355 VDD.n11677 VDD.n11676 4.5
R8356 VDD.n11712 VDD.n11711 4.5
R8357 VDD.n11803 VDD.n11802 4.5
R8358 VDD.n11819 VDD.n11818 4.5
R8359 VDD.n11725 VDD.n11686 4.5
R8360 VDD.n11643 VDD.n11588 4.5
R8361 VDD.n11639 VDD.n11638 4.5
R8362 VDD.n11619 VDD.n11618 4.5
R8363 VDD.n11604 VDD.n11603 4.5
R8364 VDD.n11515 VDD.n11514 4.5
R8365 VDD.n11494 VDD.n11472 4.5
R8366 VDD.n11551 VDD.n11550 4.5
R8367 VDD.n11841 VDD.n11840 4.5
R8368 VDD.n11835 VDD.n11834 4.5
R8369 VDD.n11854 VDD.n11853 4.5
R8370 VDD.n11778 VDD.n11777 4.5
R8371 VDD.n11765 VDD.n11764 4.5
R8372 VDD.n11924 VDD.n11923 4.5
R8373 VDD.n11937 VDD.n11936 4.5
R8374 VDD.n11910 VDD.n11909 4.5
R8375 VDD.n11782 VDD.n11753 4.5
R8376 VDD.n11897 VDD.n11896 4.5
R8377 VDD.n11879 VDD.n11871 4.5
R8378 VDD.n11875 VDD.n11874 4.5
R8379 VDD.n10165 VDD.n10164 4.444
R8380 VDD.n10095 VDD.n10093 4.444
R8381 VDD.n10038 VDD.n10036 4.444
R8382 VDD.n10283 VDD.n10281 4.363
R8383 VDD.n10630 VDD.n10628 4.363
R8384 VDD.n10511 VDD.n10510 4.363
R8385 VDD.n5328 VDD.n5326 4.325
R8386 VDD.n5689 VDD.n5687 4.325
R8387 VDD.n6051 VDD.n6049 4.325
R8388 VDD.n6413 VDD.n6411 4.325
R8389 VDD.n6775 VDD.n6773 4.325
R8390 VDD.n7137 VDD.n7135 4.325
R8391 VDD.n7499 VDD.n7497 4.325
R8392 VDD.n7861 VDD.n7859 4.325
R8393 VDD.n8223 VDD.n8221 4.325
R8394 VDD.n8585 VDD.n8583 4.325
R8395 VDD.n8947 VDD.n8945 4.325
R8396 VDD.n9309 VDD.n9307 4.325
R8397 VDD.n9671 VDD.n9669 4.325
R8398 VDD.n5664 VDD.t18 4.289
R8399 VDD.n6025 VDD.t33 4.289
R8400 VDD.n6387 VDD.t14 4.289
R8401 VDD.n6749 VDD.t31 4.289
R8402 VDD.n7111 VDD.t42 4.289
R8403 VDD.n7473 VDD.t16 4.289
R8404 VDD.n7835 VDD.t53 4.289
R8405 VDD.n8197 VDD.t12 4.289
R8406 VDD.n8559 VDD.t49 4.289
R8407 VDD.n8921 VDD.t38 4.289
R8408 VDD.n9283 VDD.t47 4.289
R8409 VDD.n9645 VDD.t51 4.289
R8410 VDD.n10007 VDD.t59 4.289
R8411 VDD.n10237 VDD.n10235 4.252
R8412 VDD.n10120 VDD.n10118 4.252
R8413 VDD.n10584 VDD.n10582 4.25
R8414 VDD.n10466 VDD.n10464 4.25
R8415 VDD.n10176 VDD.n10175 4.137
R8416 VDD.n10081 VDD.n10080 4.137
R8417 VDD.n10049 VDD.n10048 4.137
R8418 VDD.n250 VDD.n249 4.137
R8419 VDD.n526 VDD.n525 4.137
R8420 VDD.n550 VDD.n549 4.137
R8421 VDD.n760 VDD.n759 4.137
R8422 VDD.n784 VDD.n783 4.137
R8423 VDD.n993 VDD.n992 4.137
R8424 VDD.n1017 VDD.n1016 4.137
R8425 VDD.n1227 VDD.n1226 4.137
R8426 VDD.n1251 VDD.n1250 4.137
R8427 VDD.n1460 VDD.n1459 4.137
R8428 VDD.n1484 VDD.n1483 4.137
R8429 VDD.n1694 VDD.n1693 4.137
R8430 VDD.n1718 VDD.n1717 4.137
R8431 VDD.n2012 VDD.n2011 4.137
R8432 VDD.n224 VDD.n219 4.136
R8433 VDD.n10687 VDD.n10575 4.113
R8434 VDD.n10566 VDD.n10457 4.113
R8435 VDD.n10340 VDD.n10228 4.113
R8436 VDD.n10220 VDD.n10111 4.113
R8437 VDD.n10294 VDD.n10293 4.063
R8438 VDD.n10641 VDD.n10640 4.063
R8439 VDD.n10522 VDD.n10521 4.063
R8440 VDD.n12226 VDD.n11949 4.013
R8441 VDD.n11459 VDD.n11458 4.013
R8442 VDD.n2857 VDD.n2856 4.013
R8443 VDD.n4499 VDD.n4498 4.013
R8444 VDD.n5335 VDD.n5332 3.95
R8445 VDD.n5696 VDD.n5693 3.95
R8446 VDD.n6058 VDD.n6055 3.95
R8447 VDD.n6420 VDD.n6417 3.95
R8448 VDD.n6782 VDD.n6779 3.95
R8449 VDD.n7144 VDD.n7141 3.95
R8450 VDD.n7506 VDD.n7503 3.95
R8451 VDD.n7868 VDD.n7865 3.95
R8452 VDD.n8230 VDD.n8227 3.95
R8453 VDD.n8592 VDD.n8589 3.95
R8454 VDD.n8954 VDD.n8951 3.95
R8455 VDD.n9316 VDD.n9313 3.95
R8456 VDD.n9678 VDD.n9675 3.95
R8457 VDD.n5628 VDD.n5627 3.948
R8458 VDD.n5989 VDD.n5988 3.948
R8459 VDD.n6351 VDD.n6350 3.948
R8460 VDD.n6713 VDD.n6712 3.948
R8461 VDD.n7075 VDD.n7074 3.948
R8462 VDD.n7437 VDD.n7436 3.948
R8463 VDD.n7799 VDD.n7798 3.948
R8464 VDD.n8161 VDD.n8160 3.948
R8465 VDD.n8523 VDD.n8522 3.948
R8466 VDD.n8885 VDD.n8884 3.948
R8467 VDD.n9247 VDD.n9246 3.948
R8468 VDD.n9609 VDD.n9608 3.948
R8469 VDD.n9971 VDD.n9970 3.948
R8470 VDD.n2156 VDD.n2149 3.938
R8471 VDD.n2177 VDD.n2169 3.938
R8472 VDD.n2387 VDD.n2380 3.938
R8473 VDD.n2408 VDD.n2400 3.938
R8474 VDD.n5221 VDD.n5214 3.938
R8475 VDD.n5287 VDD.n5280 3.938
R8476 VDD.n5012 VDD.n5004 3.938
R8477 VDD.n4991 VDD.n4984 3.938
R8478 VDD.n4781 VDD.n4773 3.938
R8479 VDD.n4760 VDD.n4753 3.938
R8480 VDD.n2033 VDD.n2031 3.894
R8481 VDD.n4637 VDD.n4635 3.894
R8482 VDD.n10074 VDD.n10072 3.869
R8483 VDD.n10029 VDD.n10027 3.867
R8484 VDD.n37 VDD.n35 3.783
R8485 VDD.n12268 VDD.n12266 3.781
R8486 VDD.n10057 VDD.n10020 3.734
R8487 VDD.n10102 VDD.n10065 3.734
R8488 VDD.n87 VDD.n29 3.692
R8489 VDD.n12318 VDD.n12260 3.692
R8490 VDD.n2043 VDD.n2039 3.692
R8491 VDD.n2057 VDD.n2053 3.692
R8492 VDD.n2274 VDD.n2270 3.692
R8493 VDD.n2288 VDD.n2284 3.692
R8494 VDD.n2513 VDD.n2509 3.692
R8495 VDD.n2583 VDD.n2579 3.692
R8496 VDD.n2738 VDD.n2734 3.692
R8497 VDD.n5116 VDD.n5112 3.692
R8498 VDD.n4892 VDD.n4888 3.692
R8499 VDD.n4878 VDD.n4874 3.692
R8500 VDD.n4661 VDD.n4657 3.692
R8501 VDD.n4647 VDD.n4643 3.692
R8502 VDD.n2037 VDD.n2036 3.692
R8503 VDD.n2051 VDD.n2050 3.692
R8504 VDD.n2268 VDD.n2267 3.692
R8505 VDD.n2282 VDD.n2281 3.692
R8506 VDD.n4886 VDD.n4885 3.692
R8507 VDD.n4872 VDD.n4871 3.692
R8508 VDD.n4655 VDD.n4654 3.692
R8509 VDD.n4641 VDD.n4640 3.692
R8510 VDD.n11307 VDD.n11306 3.636
R8511 VDD.n12096 VDD.n12095 3.636
R8512 VDD.n12076 VDD.n12075 3.636
R8513 VDD.n10939 VDD.n10938 3.636
R8514 VDD.n11031 VDD.n11030 3.636
R8515 VDD.n10814 VDD.n10813 3.636
R8516 VDD.n10739 VDD.n10738 3.636
R8517 VDD.n11798 VDD.n11797 3.636
R8518 VDD.n11510 VDD.n11509 3.636
R8519 VDD.n5614 VDD.n5613 3.573
R8520 VDD.n5975 VDD.n5974 3.573
R8521 VDD.n6337 VDD.n6336 3.573
R8522 VDD.n6699 VDD.n6698 3.573
R8523 VDD.n7061 VDD.n7060 3.573
R8524 VDD.n7423 VDD.n7422 3.573
R8525 VDD.n7785 VDD.n7784 3.573
R8526 VDD.n8147 VDD.n8146 3.573
R8527 VDD.n8509 VDD.n8508 3.573
R8528 VDD.n8871 VDD.n8870 3.573
R8529 VDD.n9233 VDD.n9232 3.573
R8530 VDD.n9595 VDD.n9594 3.573
R8531 VDD.n9957 VDD.n9956 3.573
R8532 VDD.n11342 VDD.n11341 3.566
R8533 VDD.n12108 VDD.n12107 3.566
R8534 VDD.n12064 VDD.n12063 3.566
R8535 VDD.n12109 VDD.n12108 3.566
R8536 VDD.n12063 VDD.n12062 3.566
R8537 VDD.n10924 VDD.n10923 3.566
R8538 VDD.n11048 VDD.n11047 3.566
R8539 VDD.n10833 VDD.n10832 3.566
R8540 VDD.n10752 VDD.n10751 3.566
R8541 VDD.n10925 VDD.n10924 3.566
R8542 VDD.n10834 VDD.n10833 3.566
R8543 VDD.n11047 VDD.n11046 3.566
R8544 VDD.n10751 VDD.n10750 3.566
R8545 VDD.n11706 VDD.n11705 3.566
R8546 VDD.n11614 VDD.n11613 3.566
R8547 VDD.n11705 VDD.n11704 3.566
R8548 VDD.n11613 VDD.n11612 3.566
R8549 VDD.n11341 VDD.n11340 3.566
R8550 VDD.n10291 VDD.n10290 3.555
R8551 VDD.n10278 VDD.n10277 3.555
R8552 VDD.n10173 VDD.n10172 3.555
R8553 VDD.n10161 VDD.n10160 3.555
R8554 VDD.n10090 VDD.n10089 3.555
R8555 VDD.n10078 VDD.n10077 3.555
R8556 VDD.n10046 VDD.n10045 3.555
R8557 VDD.n10033 VDD.n10032 3.555
R8558 VDD.n10638 VDD.n10637 3.555
R8559 VDD.n10625 VDD.n10624 3.555
R8560 VDD.n10519 VDD.n10518 3.555
R8561 VDD.n10507 VDD.n10506 3.555
R8562 VDD.n10129 VDD.n10128 3.51
R8563 VDD.n10095 VDD.n10094 3.51
R8564 VDD.n10038 VDD.n10037 3.51
R8565 VDD.n10283 VDD.n10282 3.47
R8566 VDD.n10258 VDD.n10257 3.47
R8567 VDD.n10333 VDD.n10332 3.47
R8568 VDD.n10308 VDD.n10307 3.47
R8569 VDD.n10630 VDD.n10629 3.47
R8570 VDD.n10605 VDD.n10604 3.47
R8571 VDD.n10680 VDD.n10679 3.47
R8572 VDD.n10655 VDD.n10654 3.47
R8573 VDD.n10475 VDD.n10474 3.47
R8574 VDD.n2142 VDD.n2135 3.446
R8575 VDD.n2191 VDD.n2184 3.446
R8576 VDD.n2373 VDD.n2366 3.446
R8577 VDD.n2422 VDD.n2415 3.446
R8578 VDD.n5201 VDD.n5194 3.446
R8579 VDD.n5268 VDD.n5261 3.446
R8580 VDD.n5026 VDD.n5019 3.446
R8581 VDD.n4977 VDD.n4970 3.446
R8582 VDD.n4795 VDD.n4788 3.446
R8583 VDD.n4746 VDD.n4739 3.446
R8584 VDD.n10449 VDD.n10103 3.361
R8585 VDD.n10169 VDD.n10168 3.347
R8586 VDD.n10042 VDD.n10041 3.347
R8587 VDD.n10086 VDD.n10085 3.347
R8588 VDD.n2804 VDD.n2803 3.321
R8589 VDD.n3108 VDD.n3107 3.321
R8590 VDD.n3125 VDD.n3124 3.321
R8591 VDD.n3346 VDD.n3345 3.321
R8592 VDD.n3363 VDD.n3362 3.321
R8593 VDD.n3583 VDD.n3582 3.321
R8594 VDD.n3600 VDD.n3599 3.321
R8595 VDD.n3821 VDD.n3820 3.321
R8596 VDD.n3838 VDD.n3837 3.321
R8597 VDD.n4058 VDD.n4057 3.321
R8598 VDD.n4075 VDD.n4074 3.321
R8599 VDD.n4296 VDD.n4295 3.321
R8600 VDD.n4313 VDD.n4312 3.321
R8601 VDD.n4619 VDD.n4618 3.321
R8602 VDD.n4631 VDD.n4630 3.321
R8603 VDD.n2153 VDD.n2152 3.321
R8604 VDD.n2174 VDD.n2173 3.321
R8605 VDD.n2384 VDD.n2383 3.321
R8606 VDD.n2405 VDD.n2404 3.321
R8607 VDD.n5218 VDD.n5217 3.321
R8608 VDD.n5284 VDD.n5283 3.321
R8609 VDD.n5008 VDD.n5007 3.321
R8610 VDD.n4988 VDD.n4987 3.321
R8611 VDD.n4777 VDD.n4776 3.321
R8612 VDD.n4757 VDD.n4756 3.321
R8613 VDD.n419 VDD.n418 3.321
R8614 VDD.n431 VDD.n430 3.321
R8615 VDD.n652 VDD.n651 3.321
R8616 VDD.n664 VDD.n663 3.321
R8617 VDD.n886 VDD.n885 3.321
R8618 VDD.n898 VDD.n897 3.321
R8619 VDD.n1033 VDD.n1032 3.321
R8620 VDD.n1119 VDD.n1118 3.321
R8621 VDD.n1131 VDD.n1130 3.321
R8622 VDD.n1353 VDD.n1352 3.321
R8623 VDD.n1365 VDD.n1364 3.321
R8624 VDD.n1586 VDD.n1585 3.321
R8625 VDD.n1598 VDD.n1597 3.321
R8626 VDD.n1820 VDD.n1819 3.321
R8627 VDD.n1832 VDD.n1831 3.321
R8628 VDD.n10515 VDD.n10514 3.309
R8629 VDD.n10287 VDD.n10286 3.309
R8630 VDD.n10634 VDD.n10633 3.309
R8631 VDD.n3001 VDD.n2995 3.247
R8632 VDD.n3238 VDD.n3233 3.247
R8633 VDD.n3476 VDD.n3470 3.247
R8634 VDD.n3713 VDD.n3708 3.247
R8635 VDD.n3951 VDD.n3945 3.247
R8636 VDD.n4188 VDD.n4183 3.247
R8637 VDD.n4426 VDD.n4420 3.247
R8638 VDD.n197 VDD.n196 3.2
R8639 VDD.n2065 VDD.n2064 3.2
R8640 VDD.n2254 VDD.n2253 3.2
R8641 VDD.n2296 VDD.n2295 3.2
R8642 VDD.n4900 VDD.n4899 3.2
R8643 VDD.n4858 VDD.n4857 3.2
R8644 VDD.n4669 VDD.n4668 3.2
R8645 VDD.n2766 VDD.n2765 3.2
R8646 VDD.n62 VDD.n61 3.103
R8647 VDD.n54 VDD.n53 3.103
R8648 VDD.n12190 VDD.n12189 3.103
R8649 VDD.n12181 VDD.n12180 3.103
R8650 VDD.n11986 VDD.n11985 3.103
R8651 VDD.n11977 VDD.n11976 3.103
R8652 VDD.n11068 VDD.n11067 3.103
R8653 VDD.n10992 VDD.n10986 3.103
R8654 VDD.n11165 VDD.n11157 3.103
R8655 VDD.n11179 VDD.n11170 3.103
R8656 VDD.n11172 VDD.n11171 3.103
R8657 VDD.n11143 VDD.n11142 3.103
R8658 VDD.n11151 VDD.n11150 3.103
R8659 VDD.n10743 VDD.n10742 3.103
R8660 VDD.n10757 VDD.n10756 3.103
R8661 VDD.n11834 VDD.n11833 3.103
R8662 VDD.n11761 VDD.n11756 3.103
R8663 VDD.n11923 VDD.n11915 3.103
R8664 VDD.n11936 VDD.n11928 3.103
R8665 VDD.n11930 VDD.n11929 3.103
R8666 VDD.n11902 VDD.n11901 3.103
R8667 VDD.n11909 VDD.n11908 3.103
R8668 VDD.n11514 VDD.n11513 3.103
R8669 VDD.n11527 VDD.n11526 3.103
R8670 VDD.n11419 VDD.n11418 3.103
R8671 VDD.n11411 VDD.n11410 3.103
R8672 VDD.n11221 VDD.n11220 3.103
R8673 VDD.n11213 VDD.n11212 3.103
R8674 VDD.n12293 VDD.n12292 3.103
R8675 VDD.n12285 VDD.n12284 3.103
R8676 VDD.n46 VDD.n45 3.084
R8677 VDD.n80 VDD.n79 3.084
R8678 VDD.n12186 VDD.n12185 3.084
R8679 VDD.n12161 VDD.n12160 3.084
R8680 VDD.n12136 VDD.n12135 3.084
R8681 VDD.n12111 VDD.n12110 3.084
R8682 VDD.n11982 VDD.n11981 3.084
R8683 VDD.n10880 VDD.n10879 3.084
R8684 VDD.n10904 VDD.n10903 3.084
R8685 VDD.n10927 VDD.n10926 3.084
R8686 VDD.n11148 VDD.n11147 3.084
R8687 VDD.n11132 VDD.n11131 3.084
R8688 VDD.n10869 VDD.n10868 3.084
R8689 VDD.n10836 VDD.n10835 3.084
R8690 VDD.n10696 VDD.n10695 3.084
R8691 VDD.n10754 VDD.n10753 3.084
R8692 VDD.n11050 VDD.n11049 3.084
R8693 VDD.n11082 VDD.n11081 3.084
R8694 VDD.n10991 VDD.n10990 3.084
R8695 VDD.n11177 VDD.n11176 3.084
R8696 VDD.n10706 VDD.n10705 3.084
R8697 VDD.n12195 VDD.n12194 3.084
R8698 VDD.n12066 VDD.n12065 3.084
R8699 VDD.n12041 VDD.n12040 3.084
R8700 VDD.n12016 VDD.n12015 3.084
R8701 VDD.n11991 VDD.n11990 3.084
R8702 VDD.n11331 VDD.n11330 3.084
R8703 VDD.n11205 VDD.n11204 3.084
R8704 VDD.n12277 VDD.n12276 3.084
R8705 VDD.n12311 VDD.n12310 3.084
R8706 VDD.n10303 VDD.n10302 3.081
R8707 VDD.n10266 VDD.n10265 3.081
R8708 VDD.n10185 VDD.n10184 3.081
R8709 VDD.n10149 VDD.n10148 3.081
R8710 VDD.n10059 VDD.n10058 3.081
R8711 VDD.n10067 VDD.n10066 3.081
R8712 VDD.n10014 VDD.n10013 3.081
R8713 VDD.n10022 VDD.n10021 3.081
R8714 VDD.n10650 VDD.n10649 3.081
R8715 VDD.n10613 VDD.n10612 3.081
R8716 VDD.n10531 VDD.n10530 3.081
R8717 VDD.n10495 VDD.n10494 3.081
R8718 VDD.n2786 VDD.n2776 3.056
R8719 VDD.n2994 VDD.n2993 3.056
R8720 VDD.n3006 VDD.n3005 3.056
R8721 VDD.n3111 VDD.n3102 3.056
R8722 VDD.n3128 VDD.n3120 3.056
R8723 VDD.n3232 VDD.n3231 3.056
R8724 VDD.n3243 VDD.n3242 3.056
R8725 VDD.n3349 VDD.n3340 3.056
R8726 VDD.n3366 VDD.n3358 3.056
R8727 VDD.n3469 VDD.n3468 3.056
R8728 VDD.n3481 VDD.n3480 3.056
R8729 VDD.n3586 VDD.n3577 3.056
R8730 VDD.n3603 VDD.n3595 3.056
R8731 VDD.n3707 VDD.n3706 3.056
R8732 VDD.n3718 VDD.n3717 3.056
R8733 VDD.n3824 VDD.n3815 3.056
R8734 VDD.n3841 VDD.n3833 3.056
R8735 VDD.n3944 VDD.n3943 3.056
R8736 VDD.n3956 VDD.n3955 3.056
R8737 VDD.n4061 VDD.n4052 3.056
R8738 VDD.n4078 VDD.n4070 3.056
R8739 VDD.n4182 VDD.n4181 3.056
R8740 VDD.n4193 VDD.n4192 3.056
R8741 VDD.n4299 VDD.n4290 3.056
R8742 VDD.n4316 VDD.n4308 3.056
R8743 VDD.n4419 VDD.n4418 3.056
R8744 VDD.n4431 VDD.n4430 3.056
R8745 VDD.n5519 VDD.n5517 3.033
R8746 VDD.n5637 VDD.n5636 3.033
R8747 VDD.n5880 VDD.n5878 3.033
R8748 VDD.n5998 VDD.n5997 3.033
R8749 VDD.n6242 VDD.n6240 3.033
R8750 VDD.n6360 VDD.n6359 3.033
R8751 VDD.n6604 VDD.n6602 3.033
R8752 VDD.n6722 VDD.n6721 3.033
R8753 VDD.n6966 VDD.n6964 3.033
R8754 VDD.n7084 VDD.n7083 3.033
R8755 VDD.n7328 VDD.n7326 3.033
R8756 VDD.n7446 VDD.n7445 3.033
R8757 VDD.n7690 VDD.n7688 3.033
R8758 VDD.n7808 VDD.n7807 3.033
R8759 VDD.n8052 VDD.n8050 3.033
R8760 VDD.n8170 VDD.n8169 3.033
R8761 VDD.n8414 VDD.n8412 3.033
R8762 VDD.n8532 VDD.n8531 3.033
R8763 VDD.n8776 VDD.n8774 3.033
R8764 VDD.n8894 VDD.n8893 3.033
R8765 VDD.n9138 VDD.n9136 3.033
R8766 VDD.n9256 VDD.n9255 3.033
R8767 VDD.n9500 VDD.n9498 3.033
R8768 VDD.n9618 VDD.n9617 3.033
R8769 VDD.n9862 VDD.n9860 3.033
R8770 VDD.n9980 VDD.n9979 3.033
R8771 VDD.n10935 VDD.n10932 3.033
R8772 VDD.n11021 VDD.n11020 3.033
R8773 VDD.n10845 VDD.n10810 3.033
R8774 VDD.n10729 VDD.n10728 3.033
R8775 VDD.n11134 VDD.n11133 3.033
R8776 VDD.n11690 VDD.n11689 3.033
R8777 VDD.n11788 VDD.n11787 3.033
R8778 VDD.n11626 VDD.n11625 3.033
R8779 VDD.n11500 VDD.n11499 3.033
R8780 VDD.n11883 VDD.n11863 3.033
R8781 VDD.n2905 VDD.n2904 3
R8782 VDD.n4539 VDD.n4538 3
R8783 VDD.n2802 VDD.n2801 3
R8784 VDD.n3106 VDD.n3105 3
R8785 VDD.n3122 VDD.n3121 3
R8786 VDD.n3344 VDD.n3343 3
R8787 VDD.n3360 VDD.n3359 3
R8788 VDD.n3581 VDD.n3580 3
R8789 VDD.n3597 VDD.n3596 3
R8790 VDD.n3819 VDD.n3818 3
R8791 VDD.n3835 VDD.n3834 3
R8792 VDD.n4056 VDD.n4055 3
R8793 VDD.n4072 VDD.n4071 3
R8794 VDD.n4294 VDD.n4293 3
R8795 VDD.n4310 VDD.n4309 3
R8796 VDD.n4617 VDD.n4616 3
R8797 VDD.n2128 VDD.n2121 2.953
R8798 VDD.n2205 VDD.n2198 2.953
R8799 VDD.n2359 VDD.n2352 2.953
R8800 VDD.n2436 VDD.n2429 2.953
R8801 VDD.n2495 VDD.n2484 2.953
R8802 VDD.n5180 VDD.n5173 2.953
R8803 VDD.n5247 VDD.n5240 2.953
R8804 VDD.n5040 VDD.n5033 2.953
R8805 VDD.n4963 VDD.n4956 2.953
R8806 VDD.n4809 VDD.n4802 2.953
R8807 VDD.n4732 VDD.n4725 2.953
R8808 VDD.n12099 VDD.n12094 2.909
R8809 VDD.n12079 VDD.n12074 2.909
R8810 VDD.n10930 VDD.n10929 2.909
R8811 VDD.n10942 VDD.n10937 2.909
R8812 VDD.n11035 VDD.n11034 2.909
R8813 VDD.n11034 VDD.n11029 2.909
R8814 VDD.n11116 VDD.n11115 2.909
R8815 VDD.n10839 VDD.n10837 2.909
R8816 VDD.n10817 VDD.n10812 2.909
R8817 VDD.n10819 VDD.n10817 2.909
R8818 VDD.n11710 VDD.n11709 2.909
R8819 VDD.n11699 VDD.n11692 2.909
R8820 VDD.n11802 VDD.n11801 2.909
R8821 VDD.n11801 VDD.n11796 2.909
R8822 VDD.n11896 VDD.n11895 2.909
R8823 VDD.n11618 VDD.n11616 2.909
R8824 VDD.n11601 VDD.n11594 2.909
R8825 VDD.n11603 VDD.n11601 2.909
R8826 VDD.n11332 VDD.n11325 2.909
R8827 VDD.n11310 VDD.n11305 2.909
R8828 VDD.n2786 VDD.n2778 2.865
R8829 VDD.n2982 VDD.n2981 2.865
R8830 VDD.n3004 VDD.n3003 2.865
R8831 VDD.n3111 VDD.n3104 2.865
R8832 VDD.n3142 VDD.n3133 2.865
R8833 VDD.n3220 VDD.n3219 2.865
R8834 VDD.n3241 VDD.n3240 2.865
R8835 VDD.n3349 VDD.n3342 2.865
R8836 VDD.n3380 VDD.n3371 2.865
R8837 VDD.n3457 VDD.n3456 2.865
R8838 VDD.n3479 VDD.n3478 2.865
R8839 VDD.n3586 VDD.n3579 2.865
R8840 VDD.n3617 VDD.n3608 2.865
R8841 VDD.n3695 VDD.n3694 2.865
R8842 VDD.n3716 VDD.n3715 2.865
R8843 VDD.n3824 VDD.n3817 2.865
R8844 VDD.n3855 VDD.n3846 2.865
R8845 VDD.n3932 VDD.n3931 2.865
R8846 VDD.n3954 VDD.n3953 2.865
R8847 VDD.n4061 VDD.n4054 2.865
R8848 VDD.n4092 VDD.n4083 2.865
R8849 VDD.n4170 VDD.n4169 2.865
R8850 VDD.n4191 VDD.n4190 2.865
R8851 VDD.n4299 VDD.n4292 2.865
R8852 VDD.n4330 VDD.n4321 2.865
R8853 VDD.n4407 VDD.n4406 2.865
R8854 VDD.n4429 VDD.n4428 2.865
R8855 VDD.n11461 VDD.n11460 2.859
R8856 VDD.n12228 VDD.n12227 2.851
R8857 VDD.n11194 VDD.n11193 2.793
R8858 VDD.n11959 VDD.n11958 2.793
R8859 VDD.n1932 VDD.n1931 2.787
R8860 VDD.n75 VDD.n74 2.715
R8861 VDD.n41 VDD.n40 2.715
R8862 VDD.n12203 VDD.n12202 2.715
R8863 VDD.n12169 VDD.n12168 2.715
R8864 VDD.n11999 VDD.n11998 2.715
R8865 VDD.n11965 VDD.n11964 2.715
R8866 VDD.n11052 VDD.n11051 2.715
R8867 VDD.n11159 VDD.n11158 2.715
R8868 VDD.n11108 VDD.n11107 2.715
R8869 VDD.n10737 VDD.n10736 2.715
R8870 VDD.n11818 VDD.n11817 2.715
R8871 VDD.n11917 VDD.n11916 2.715
R8872 VDD.n11888 VDD.n11887 2.715
R8873 VDD.n11508 VDD.n11507 2.715
R8874 VDD.n11431 VDD.n11430 2.715
R8875 VDD.n11399 VDD.n11398 2.715
R8876 VDD.n11233 VDD.n11232 2.715
R8877 VDD.n11200 VDD.n11199 2.715
R8878 VDD.n12306 VDD.n12305 2.715
R8879 VDD.n12272 VDD.n12271 2.715
R8880 VDD.n2079 VDD.n2078 2.707
R8881 VDD.n2240 VDD.n2239 2.707
R8882 VDD.n2310 VDD.n2309 2.707
R8883 VDD.n2471 VDD.n2470 2.707
R8884 VDD.n5183 VDD.n5180 2.707
R8885 VDD.n5182 VDD.n5181 2.707
R8886 VDD.n5288 VDD.n5278 2.707
R8887 VDD.n2740 VDD.n2739 2.707
R8888 VDD.n5099 VDD.n5098 2.707
R8889 VDD.n5075 VDD.n5074 2.707
R8890 VDD.n4914 VDD.n4913 2.707
R8891 VDD.n4844 VDD.n4843 2.707
R8892 VDD.n4683 VDD.n4682 2.707
R8893 VDD.n1933 VDD.n1929 2.695
R8894 VDD.n318 VDD.n317 2.695
R8895 VDD.n2980 VDD.n2979 2.674
R8896 VDD.n3020 VDD.n3019 2.674
R8897 VDD.n3097 VDD.n3088 2.674
R8898 VDD.n3142 VDD.n3135 2.674
R8899 VDD.n3218 VDD.n3217 2.674
R8900 VDD.n3257 VDD.n3256 2.674
R8901 VDD.n3335 VDD.n3326 2.674
R8902 VDD.n3380 VDD.n3373 2.674
R8903 VDD.n3455 VDD.n3454 2.674
R8904 VDD.n3495 VDD.n3494 2.674
R8905 VDD.n3572 VDD.n3563 2.674
R8906 VDD.n3617 VDD.n3610 2.674
R8907 VDD.n3693 VDD.n3692 2.674
R8908 VDD.n3732 VDD.n3731 2.674
R8909 VDD.n3810 VDD.n3801 2.674
R8910 VDD.n3855 VDD.n3848 2.674
R8911 VDD.n3930 VDD.n3929 2.674
R8912 VDD.n3970 VDD.n3969 2.674
R8913 VDD.n4047 VDD.n4038 2.674
R8914 VDD.n4092 VDD.n4085 2.674
R8915 VDD.n4168 VDD.n4167 2.674
R8916 VDD.n4207 VDD.n4206 2.674
R8917 VDD.n4285 VDD.n4276 2.674
R8918 VDD.n4330 VDD.n4323 2.674
R8919 VDD.n4405 VDD.n4404 2.674
R8920 VDD.n4445 VDD.n4444 2.674
R8921 VDD.n10316 VDD.n10315 2.607
R8922 VDD.n10253 VDD.n10252 2.607
R8923 VDD.n10197 VDD.n10196 2.607
R8924 VDD.n10137 VDD.n10136 2.607
R8925 VDD.n10663 VDD.n10662 2.607
R8926 VDD.n10600 VDD.n10599 2.607
R8927 VDD.n10543 VDD.n10542 2.607
R8928 VDD.n10483 VDD.n10482 2.607
R8929 VDD.n10890 VDD.n10883 2.601
R8930 VDD.n10716 VDD.n10709 2.601
R8931 VDD.n11659 VDD.n11652 2.601
R8932 VDD.n11486 VDD.n11479 2.601
R8933 VDD.n12112 VDD.n12106 2.521
R8934 VDD.n12067 VDD.n12061 2.521
R8935 VDD.n10928 VDD.n10922 2.521
R8936 VDD.n10755 VDD.n10749 2.521
R8937 VDD.n11708 VDD.n11703 2.521
R8938 VDD.n11525 VDD.n11520 2.521
R8939 VDD.n11344 VDD.n11339 2.521
R8940 VDD.n11298 VDD.n11293 2.521
R8941 VDD.n2968 VDD.n2967 2.483
R8942 VDD.n3018 VDD.n3017 2.483
R8943 VDD.n3097 VDD.n3090 2.483
R8944 VDD.n3157 VDD.n3147 2.483
R8945 VDD.n3206 VDD.n3205 2.483
R8946 VDD.n3255 VDD.n3254 2.483
R8947 VDD.n3335 VDD.n3328 2.483
R8948 VDD.n3394 VDD.n3385 2.483
R8949 VDD.n3443 VDD.n3442 2.483
R8950 VDD.n3493 VDD.n3492 2.483
R8951 VDD.n3572 VDD.n3565 2.483
R8952 VDD.n3632 VDD.n3622 2.483
R8953 VDD.n3681 VDD.n3680 2.483
R8954 VDD.n3730 VDD.n3729 2.483
R8955 VDD.n3810 VDD.n3803 2.483
R8956 VDD.n3869 VDD.n3860 2.483
R8957 VDD.n3918 VDD.n3917 2.483
R8958 VDD.n3968 VDD.n3967 2.483
R8959 VDD.n4047 VDD.n4040 2.483
R8960 VDD.n4107 VDD.n4097 2.483
R8961 VDD.n4156 VDD.n4155 2.483
R8962 VDD.n4205 VDD.n4204 2.483
R8963 VDD.n4285 VDD.n4278 2.483
R8964 VDD.n4344 VDD.n4335 2.483
R8965 VDD.n4393 VDD.n4392 2.483
R8966 VDD.n4443 VDD.n4442 2.483
R8967 VDD.n2114 VDD.n2107 2.461
R8968 VDD.n2219 VDD.n2212 2.461
R8969 VDD.n2345 VDD.n2338 2.461
R8970 VDD.n2450 VDD.n2443 2.461
R8971 VDD.n2515 VDD.n2504 2.461
R8972 VDD.n2541 VDD.n2540 2.461
R8973 VDD.n2552 VDD.n2551 2.461
R8974 VDD.n2562 VDD.n2560 2.461
R8975 VDD.n5162 VDD.n5155 2.461
R8976 VDD.n5164 VDD.n5162 2.461
R8977 VDD.n5223 VDD.n5222 2.461
R8978 VDD.n5231 VDD.n5227 2.461
R8979 VDD.n5238 VDD.n5237 2.461
R8980 VDD.n5248 VDD.n5247 2.461
R8981 VDD.n2644 VDD.n2643 2.461
R8982 VDD.n2643 VDD.n2636 2.461
R8983 VDD.n2668 VDD.n2657 2.461
R8984 VDD.n2746 VDD.n2744 2.461
R8985 VDD.n2763 VDD.n2762 2.461
R8986 VDD.n5054 VDD.n5047 2.461
R8987 VDD.n4949 VDD.n4942 2.461
R8988 VDD.n4823 VDD.n4816 2.461
R8989 VDD.n4718 VDD.n4711 2.461
R8990 VDD.n12230 VDD.n5307 2.387
R8991 VDD.n10228 VDD.n10222 2.37
R8992 VDD.n10235 VDD.n10230 2.37
R8993 VDD.n10111 VDD.n10105 2.37
R8994 VDD.n10118 VDD.n10113 2.37
R8995 VDD.n10575 VDD.n10569 2.37
R8996 VDD.n10582 VDD.n10577 2.37
R8997 VDD.n10457 VDD.n10451 2.37
R8998 VDD.n10464 VDD.n10459 2.37
R8999 VDD.n24 VDD.n23 2.327
R9000 VDD.n31 VDD.n30 2.327
R9001 VDD.n12215 VDD.n12214 2.327
R9002 VDD.n12156 VDD.n12155 2.327
R9003 VDD.n12011 VDD.n12010 2.327
R9004 VDD.n11953 VDD.n11952 2.327
R9005 VDD.n10994 VDD.n10993 2.327
R9006 VDD.n11120 VDD.n11119 2.327
R9007 VDD.n10699 VDD.n10698 2.327
R9008 VDD.n11763 VDD.n11762 2.327
R9009 VDD.n11857 VDD.n11856 2.327
R9010 VDD.n11471 VDD.n11470 2.327
R9011 VDD.n11443 VDD.n11442 2.327
R9012 VDD.n11387 VDD.n11386 2.327
R9013 VDD.n11245 VDD.n11244 2.327
R9014 VDD.n11189 VDD.n11188 2.327
R9015 VDD.n12255 VDD.n12254 2.327
R9016 VDD.n12262 VDD.n12261 2.327
R9017 VDD.n2966 VDD.n2965 2.292
R9018 VDD.n3034 VDD.n3033 2.292
R9019 VDD.n3083 VDD.n3074 2.292
R9020 VDD.n3157 VDD.n3149 2.292
R9021 VDD.n3204 VDD.n3203 2.292
R9022 VDD.n3271 VDD.n3270 2.292
R9023 VDD.n3321 VDD.n3311 2.292
R9024 VDD.n3394 VDD.n3387 2.292
R9025 VDD.n3441 VDD.n3440 2.292
R9026 VDD.n3509 VDD.n3508 2.292
R9027 VDD.n3558 VDD.n3549 2.292
R9028 VDD.n3632 VDD.n3624 2.292
R9029 VDD.n3679 VDD.n3678 2.292
R9030 VDD.n3746 VDD.n3745 2.292
R9031 VDD.n3796 VDD.n3786 2.292
R9032 VDD.n3869 VDD.n3862 2.292
R9033 VDD.n3916 VDD.n3915 2.292
R9034 VDD.n3984 VDD.n3983 2.292
R9035 VDD.n4033 VDD.n4024 2.292
R9036 VDD.n4107 VDD.n4099 2.292
R9037 VDD.n4154 VDD.n4153 2.292
R9038 VDD.n4221 VDD.n4220 2.292
R9039 VDD.n4271 VDD.n4261 2.292
R9040 VDD.n4344 VDD.n4337 2.292
R9041 VDD.n4391 VDD.n4390 2.292
R9042 VDD.n2858 VDD.n2857 2.26
R9043 VDD.n2906 VDD.n2905 2.26
R9044 VDD.n4500 VDD.n4499 2.26
R9045 VDD.n4540 VDD.n4539 2.26
R9046 VDD.n2832 VDD.n2831 2.26
R9047 VDD.n2887 VDD.n2886 2.26
R9048 VDD.n4480 VDD.n4479 2.26
R9049 VDD.n4521 VDD.n4520 2.26
R9050 VDD.n5334 VDD.n5333 2.258
R9051 VDD.n5612 VDD.n5611 2.258
R9052 VDD.n5695 VDD.n5694 2.258
R9053 VDD.n5973 VDD.n5972 2.258
R9054 VDD.n6057 VDD.n6056 2.258
R9055 VDD.n6335 VDD.n6334 2.258
R9056 VDD.n6419 VDD.n6418 2.258
R9057 VDD.n6697 VDD.n6696 2.258
R9058 VDD.n6781 VDD.n6780 2.258
R9059 VDD.n7059 VDD.n7058 2.258
R9060 VDD.n7143 VDD.n7142 2.258
R9061 VDD.n7421 VDD.n7420 2.258
R9062 VDD.n7505 VDD.n7504 2.258
R9063 VDD.n7783 VDD.n7782 2.258
R9064 VDD.n7867 VDD.n7866 2.258
R9065 VDD.n8145 VDD.n8144 2.258
R9066 VDD.n8229 VDD.n8228 2.258
R9067 VDD.n8507 VDD.n8506 2.258
R9068 VDD.n8591 VDD.n8590 2.258
R9069 VDD.n8869 VDD.n8868 2.258
R9070 VDD.n8953 VDD.n8952 2.258
R9071 VDD.n9231 VDD.n9230 2.258
R9072 VDD.n9315 VDD.n9314 2.258
R9073 VDD.n9593 VDD.n9592 2.258
R9074 VDD.n9677 VDD.n9676 2.258
R9075 VDD.n9955 VDD.n9954 2.258
R9076 VDD.n2093 VDD.n2092 2.215
R9077 VDD.n2226 VDD.n2225 2.215
R9078 VDD.n2324 VDD.n2323 2.215
R9079 VDD.n2457 VDD.n2456 2.215
R9080 VDD.n2524 VDD.n2523 2.215
R9081 VDD.n2586 VDD.n2585 2.215
R9082 VDD.n129 VDD.n128 2.215
R9083 VDD.n139 VDD.n138 2.215
R9084 VDD.n148 VDD.n147 2.215
R9085 VDD.n5204 VDD.n5201 2.215
R9086 VDD.n5203 VDD.n5202 2.215
R9087 VDD.n5293 VDD.n5292 2.215
R9088 VDD.n5269 VDD.n5259 2.215
R9089 VDD.n2687 VDD.n2677 2.215
R9090 VDD.n2679 VDD.n2678 2.215
R9091 VDD.n2722 VDD.n2721 2.215
R9092 VDD.n2713 VDD.n2712 2.215
R9093 VDD.n2751 VDD.n2750 2.215
R9094 VDD.n5119 VDD.n5118 2.215
R9095 VDD.n5061 VDD.n5060 2.215
R9096 VDD.n4928 VDD.n4927 2.215
R9097 VDD.n4830 VDD.n4829 2.215
R9098 VDD.n4697 VDD.n4696 2.215
R9099 VDD.n2784 VDD.n2783 2.203
R9100 VDD.n411 VDD.n410 2.133
R9101 VDD.n413 VDD.n412 2.133
R9102 VDD.n424 VDD.n423 2.133
R9103 VDD.n426 VDD.n425 2.133
R9104 VDD.n645 VDD.n644 2.133
R9105 VDD.n647 VDD.n646 2.133
R9106 VDD.n657 VDD.n656 2.133
R9107 VDD.n659 VDD.n658 2.133
R9108 VDD.n878 VDD.n877 2.133
R9109 VDD.n880 VDD.n879 2.133
R9110 VDD.n891 VDD.n890 2.133
R9111 VDD.n893 VDD.n892 2.133
R9112 VDD.n1112 VDD.n1111 2.133
R9113 VDD.n1114 VDD.n1113 2.133
R9114 VDD.n1124 VDD.n1123 2.133
R9115 VDD.n1126 VDD.n1125 2.133
R9116 VDD.n1345 VDD.n1344 2.133
R9117 VDD.n1347 VDD.n1346 2.133
R9118 VDD.n1358 VDD.n1357 2.133
R9119 VDD.n1360 VDD.n1359 2.133
R9120 VDD.n1579 VDD.n1578 2.133
R9121 VDD.n1581 VDD.n1580 2.133
R9122 VDD.n1591 VDD.n1590 2.133
R9123 VDD.n1593 VDD.n1592 2.133
R9124 VDD.n1812 VDD.n1811 2.133
R9125 VDD.n1814 VDD.n1813 2.133
R9126 VDD.n1825 VDD.n1824 2.133
R9127 VDD.n1827 VDD.n1826 2.133
R9128 VDD.n10328 VDD.n10327 2.133
R9129 VDD.n10241 VDD.n10240 2.133
R9130 VDD.n10209 VDD.n10208 2.133
R9131 VDD.n10124 VDD.n10123 2.133
R9132 VDD.n10675 VDD.n10674 2.133
R9133 VDD.n10588 VDD.n10587 2.133
R9134 VDD.n10555 VDD.n10554 2.133
R9135 VDD.n10470 VDD.n10469 2.133
R9136 VDD.n12124 VDD.n12119 2.133
R9137 VDD.n12054 VDD.n12049 2.133
R9138 VDD.n10907 VDD.n10906 2.133
R9139 VDD.n10852 VDD.n10847 2.133
R9140 VDD.n10831 VDD.n10830 2.133
R9141 VDD.n11675 VDD.n11674 2.133
R9142 VDD.n11633 VDD.n11628 2.133
R9143 VDD.n11611 VDD.n11610 2.133
R9144 VDD.n11356 VDD.n11351 2.133
R9145 VDD.n11286 VDD.n11281 2.133
R9146 VDD.n3032 VDD.n3031 2.101
R9147 VDD.n3083 VDD.n3076 2.101
R9148 VDD.n3171 VDD.n3162 2.101
R9149 VDD.n3192 VDD.n3191 2.101
R9150 VDD.n3269 VDD.n3268 2.101
R9151 VDD.n3321 VDD.n3313 2.101
R9152 VDD.n3408 VDD.n3399 2.101
R9153 VDD.n3429 VDD.n3428 2.101
R9154 VDD.n3507 VDD.n3506 2.101
R9155 VDD.n3558 VDD.n3551 2.101
R9156 VDD.n3646 VDD.n3637 2.101
R9157 VDD.n3667 VDD.n3666 2.101
R9158 VDD.n3744 VDD.n3743 2.101
R9159 VDD.n3796 VDD.n3788 2.101
R9160 VDD.n3883 VDD.n3874 2.101
R9161 VDD.n3904 VDD.n3903 2.101
R9162 VDD.n3982 VDD.n3981 2.101
R9163 VDD.n4033 VDD.n4026 2.101
R9164 VDD.n4121 VDD.n4112 2.101
R9165 VDD.n4142 VDD.n4141 2.101
R9166 VDD.n4219 VDD.n4218 2.101
R9167 VDD.n4271 VDD.n4263 2.101
R9168 VDD.n4358 VDD.n4349 2.101
R9169 VDD.n4379 VDD.n4378 2.101
R9170 VDD.n1934 VDD.n1933 2.082
R9171 VDD.n1873 VDD.n1872 2.082
R9172 VDD.n1892 VDD.n1891 2.082
R9173 VDD.n1912 VDD.n1911 2.082
R9174 VDD.n235 VDD.n234 2.082
R9175 VDD.n271 VDD.n270 2.082
R9176 VDD.n301 VDD.n300 2.082
R9177 VDD.n319 VDD.n318 2.082
R9178 VDD.n420 VDD.n415 2.068
R9179 VDD.n432 VDD.n428 2.068
R9180 VDD.n653 VDD.n649 2.068
R9181 VDD.n665 VDD.n661 2.068
R9182 VDD.n887 VDD.n882 2.068
R9183 VDD.n899 VDD.n895 2.068
R9184 VDD.n1120 VDD.n1116 2.068
R9185 VDD.n1132 VDD.n1128 2.068
R9186 VDD.n1354 VDD.n1349 2.068
R9187 VDD.n1366 VDD.n1362 2.068
R9188 VDD.n1587 VDD.n1583 2.068
R9189 VDD.n1599 VDD.n1595 2.068
R9190 VDD.n1821 VDD.n1816 2.068
R9191 VDD.n1833 VDD.n1829 2.068
R9192 VDD.n208 VDD.n207 2.046
R9193 VDD.n209 VDD.n208 2.046
R9194 VDD.n531 VDD.n522 2
R9195 VDD.n531 VDD.n524 2
R9196 VDD.n555 VDD.n546 2
R9197 VDD.n555 VDD.n548 2
R9198 VDD.n765 VDD.n756 2
R9199 VDD.n765 VDD.n758 2
R9200 VDD.n789 VDD.n780 2
R9201 VDD.n789 VDD.n782 2
R9202 VDD.n998 VDD.n989 2
R9203 VDD.n998 VDD.n991 2
R9204 VDD.n1022 VDD.n1013 2
R9205 VDD.n1022 VDD.n1015 2
R9206 VDD.n1232 VDD.n1223 2
R9207 VDD.n1232 VDD.n1225 2
R9208 VDD.n1256 VDD.n1247 2
R9209 VDD.n1256 VDD.n1249 2
R9210 VDD.n1465 VDD.n1456 2
R9211 VDD.n1465 VDD.n1458 2
R9212 VDD.n1489 VDD.n1480 2
R9213 VDD.n1489 VDD.n1482 2
R9214 VDD.n1699 VDD.n1690 2
R9215 VDD.n1699 VDD.n1692 2
R9216 VDD.n1723 VDD.n1714 2
R9217 VDD.n1723 VDD.n1716 2
R9218 VDD.n214 VDD.n204 2
R9219 VDD.n214 VDD.n206 2
R9220 VDD.n2100 VDD.n2093 1.969
R9221 VDD.n2233 VDD.n2226 1.969
R9222 VDD.n2331 VDD.n2324 1.969
R9223 VDD.n2464 VDD.n2457 1.969
R9224 VDD.n2487 VDD.n2486 1.969
R9225 VDD.n2507 VDD.n2506 1.969
R9226 VDD.n119 VDD.n118 1.969
R9227 VDD.n129 VDD.n127 1.969
R9228 VDD.n146 VDD.n139 1.969
R9229 VDD.n148 VDD.n146 1.969
R9230 VDD.n5204 VDD.n5203 1.969
R9231 VDD.n5259 VDD.n5258 1.969
R9232 VDD.n5269 VDD.n5268 1.969
R9233 VDD.n2687 VDD.n2686 1.969
R9234 VDD.n2686 VDD.n2679 1.969
R9235 VDD.n2722 VDD.n2711 1.969
R9236 VDD.n5109 VDD.n5108 1.969
R9237 VDD.n5119 VDD.n5117 1.969
R9238 VDD.n5068 VDD.n5061 1.969
R9239 VDD.n4935 VDD.n4928 1.969
R9240 VDD.n4837 VDD.n4830 1.969
R9241 VDD.n4704 VDD.n4697 1.969
R9242 VDD.n12144 VDD.n12143 1.939
R9243 VDD.n12024 VDD.n12023 1.939
R9244 VDD.n11045 VDD.n11044 1.939
R9245 VDD.n11062 VDD.n11061 1.939
R9246 VDD.n11008 VDD.n11007 1.939
R9247 VDD.n11090 VDD.n11089 1.939
R9248 VDD.n11812 VDD.n11811 1.939
R9249 VDD.n11828 VDD.n11827 1.939
R9250 VDD.n11776 VDD.n11775 1.939
R9251 VDD.n11865 VDD.n11864 1.939
R9252 VDD.n11375 VDD.n11374 1.939
R9253 VDD.n11257 VDD.n11256 1.939
R9254 VDD.n3048 VDD.n3047 1.91
R9255 VDD.n3069 VDD.n3060 1.91
R9256 VDD.n3171 VDD.n3164 1.91
R9257 VDD.n3190 VDD.n3189 1.91
R9258 VDD.n3285 VDD.n3284 1.91
R9259 VDD.n3306 VDD.n3297 1.91
R9260 VDD.n3408 VDD.n3401 1.91
R9261 VDD.n3427 VDD.n3426 1.91
R9262 VDD.n3523 VDD.n3522 1.91
R9263 VDD.n3544 VDD.n3535 1.91
R9264 VDD.n3646 VDD.n3639 1.91
R9265 VDD.n3665 VDD.n3664 1.91
R9266 VDD.n3760 VDD.n3759 1.91
R9267 VDD.n3781 VDD.n3772 1.91
R9268 VDD.n3883 VDD.n3876 1.91
R9269 VDD.n3902 VDD.n3901 1.91
R9270 VDD.n3998 VDD.n3997 1.91
R9271 VDD.n4019 VDD.n4010 1.91
R9272 VDD.n4121 VDD.n4114 1.91
R9273 VDD.n4140 VDD.n4139 1.91
R9274 VDD.n4235 VDD.n4234 1.91
R9275 VDD.n4256 VDD.n4247 1.91
R9276 VDD.n4358 VDD.n4351 1.91
R9277 VDD.n4377 VDD.n4376 1.91
R9278 VDD.n4626 VDD.n4625 1.901
R9279 VDD.n10334 VDD.n10328 1.896
R9280 VDD.n10246 VDD.n10241 1.896
R9281 VDD.n10214 VDD.n10209 1.896
R9282 VDD.n10130 VDD.n10124 1.896
R9283 VDD.n10681 VDD.n10675 1.896
R9284 VDD.n10593 VDD.n10588 1.896
R9285 VDD.n10560 VDD.n10555 1.896
R9286 VDD.n10476 VDD.n10470 1.896
R9287 VDD.n5330 VDD.n5329 1.882
R9288 VDD.n5331 VDD.n5330 1.882
R9289 VDD.n5619 VDD.n5618 1.882
R9290 VDD.n5691 VDD.n5690 1.882
R9291 VDD.n5692 VDD.n5691 1.882
R9292 VDD.n5980 VDD.n5979 1.882
R9293 VDD.n6053 VDD.n6052 1.882
R9294 VDD.n6054 VDD.n6053 1.882
R9295 VDD.n6342 VDD.n6341 1.882
R9296 VDD.n6415 VDD.n6414 1.882
R9297 VDD.n6416 VDD.n6415 1.882
R9298 VDD.n6704 VDD.n6703 1.882
R9299 VDD.n6777 VDD.n6776 1.882
R9300 VDD.n6778 VDD.n6777 1.882
R9301 VDD.n7066 VDD.n7065 1.882
R9302 VDD.n7139 VDD.n7138 1.882
R9303 VDD.n7140 VDD.n7139 1.882
R9304 VDD.n7428 VDD.n7427 1.882
R9305 VDD.n7501 VDD.n7500 1.882
R9306 VDD.n7502 VDD.n7501 1.882
R9307 VDD.n7790 VDD.n7789 1.882
R9308 VDD.n7863 VDD.n7862 1.882
R9309 VDD.n7864 VDD.n7863 1.882
R9310 VDD.n8152 VDD.n8151 1.882
R9311 VDD.n8225 VDD.n8224 1.882
R9312 VDD.n8226 VDD.n8225 1.882
R9313 VDD.n8514 VDD.n8513 1.882
R9314 VDD.n8587 VDD.n8586 1.882
R9315 VDD.n8588 VDD.n8587 1.882
R9316 VDD.n8876 VDD.n8875 1.882
R9317 VDD.n8949 VDD.n8948 1.882
R9318 VDD.n8950 VDD.n8949 1.882
R9319 VDD.n9238 VDD.n9237 1.882
R9320 VDD.n9311 VDD.n9310 1.882
R9321 VDD.n9312 VDD.n9311 1.882
R9322 VDD.n9600 VDD.n9599 1.882
R9323 VDD.n9673 VDD.n9672 1.882
R9324 VDD.n9674 VDD.n9673 1.882
R9325 VDD.n9962 VDD.n9961 1.882
R9326 VDD.n397 VDD.n396 1.866
R9327 VDD.n399 VDD.n398 1.866
R9328 VDD.n438 VDD.n437 1.866
R9329 VDD.n440 VDD.n439 1.866
R9330 VDD.n631 VDD.n630 1.866
R9331 VDD.n633 VDD.n632 1.866
R9332 VDD.n671 VDD.n670 1.866
R9333 VDD.n673 VDD.n672 1.866
R9334 VDD.n864 VDD.n863 1.866
R9335 VDD.n866 VDD.n865 1.866
R9336 VDD.n905 VDD.n904 1.866
R9337 VDD.n907 VDD.n906 1.866
R9338 VDD.n1098 VDD.n1097 1.866
R9339 VDD.n1100 VDD.n1099 1.866
R9340 VDD.n1138 VDD.n1137 1.866
R9341 VDD.n1140 VDD.n1139 1.866
R9342 VDD.n1331 VDD.n1330 1.866
R9343 VDD.n1333 VDD.n1332 1.866
R9344 VDD.n1372 VDD.n1371 1.866
R9345 VDD.n1374 VDD.n1373 1.866
R9346 VDD.n1565 VDD.n1564 1.866
R9347 VDD.n1567 VDD.n1566 1.866
R9348 VDD.n1605 VDD.n1604 1.866
R9349 VDD.n1607 VDD.n1606 1.866
R9350 VDD.n1798 VDD.n1797 1.866
R9351 VDD.n1800 VDD.n1799 1.866
R9352 VDD.n1839 VDD.n1838 1.866
R9353 VDD.n1841 VDD.n1840 1.866
R9354 VDD.n2151 VDD.n2150 1.846
R9355 VDD.n2171 VDD.n2170 1.846
R9356 VDD.n2382 VDD.n2381 1.846
R9357 VDD.n2402 VDD.n2401 1.846
R9358 VDD.n5216 VDD.n5215 1.846
R9359 VDD.n5282 VDD.n5281 1.846
R9360 VDD.n5006 VDD.n5005 1.846
R9361 VDD.n4986 VDD.n4985 1.846
R9362 VDD.n4775 VDD.n4774 1.846
R9363 VDD.n4755 VDD.n4754 1.846
R9364 VDD.n5665 VDD.n5664 1.844
R9365 VDD.n6026 VDD.n6025 1.844
R9366 VDD.n6388 VDD.n6387 1.844
R9367 VDD.n6750 VDD.n6749 1.844
R9368 VDD.n7112 VDD.n7111 1.844
R9369 VDD.n7474 VDD.n7473 1.844
R9370 VDD.n7836 VDD.n7835 1.844
R9371 VDD.n8198 VDD.n8197 1.844
R9372 VDD.n8560 VDD.n8559 1.844
R9373 VDD.n8922 VDD.n8921 1.844
R9374 VDD.n9284 VDD.n9283 1.844
R9375 VDD.n9646 VDD.n9645 1.844
R9376 VDD.n10008 VDD.n10007 1.844
R9377 VDD.n11415 VDD.n11414 1.818
R9378 VDD.n11217 VDD.n11216 1.818
R9379 VDD.n12195 VDD.n12193 1.818
R9380 VDD.n12186 VDD.n12184 1.818
R9381 VDD.n11991 VDD.n11989 1.818
R9382 VDD.n11982 VDD.n11980 1.818
R9383 VDD.n11177 VDD.n11175 1.818
R9384 VDD.n11148 VDD.n11146 1.818
R9385 VDD.n11906 VDD.n11905 1.818
R9386 VDD.n212 VDD.n211 1.806
R9387 VDD.n11328 VDD.n11327 1.801
R9388 VDD.n11695 VDD.n11694 1.801
R9389 VDD.n11597 VDD.n11596 1.801
R9390 VDD.n11694 VDD.n11693 1.801
R9391 VDD.n11596 VDD.n11595 1.801
R9392 VDD.n11327 VDD.n11326 1.801
R9393 VDD.n12137 VDD.n12131 1.745
R9394 VDD.n12042 VDD.n12036 1.745
R9395 VDD.n10905 VDD.n10899 1.745
R9396 VDD.n10918 VDD.n10911 1.745
R9397 VDD.n10697 VDD.n10691 1.745
R9398 VDD.n11673 VDD.n11668 1.745
R9399 VDD.n11686 VDD.n11679 1.745
R9400 VDD.n11469 VDD.n11464 1.745
R9401 VDD.n11368 VDD.n11363 1.745
R9402 VDD.n11274 VDD.n11269 1.745
R9403 VDD.n517 VDD.n508 1.733
R9404 VDD.n517 VDD.n510 1.733
R9405 VDD.n570 VDD.n560 1.733
R9406 VDD.n570 VDD.n562 1.733
R9407 VDD.n751 VDD.n742 1.733
R9408 VDD.n751 VDD.n744 1.733
R9409 VDD.n803 VDD.n794 1.733
R9410 VDD.n803 VDD.n796 1.733
R9411 VDD.n984 VDD.n975 1.733
R9412 VDD.n984 VDD.n977 1.733
R9413 VDD.n1037 VDD.n1027 1.733
R9414 VDD.n1037 VDD.n1029 1.733
R9415 VDD.n1218 VDD.n1209 1.733
R9416 VDD.n1218 VDD.n1211 1.733
R9417 VDD.n1270 VDD.n1261 1.733
R9418 VDD.n1270 VDD.n1263 1.733
R9419 VDD.n1451 VDD.n1442 1.733
R9420 VDD.n1451 VDD.n1444 1.733
R9421 VDD.n1504 VDD.n1494 1.733
R9422 VDD.n1504 VDD.n1496 1.733
R9423 VDD.n1685 VDD.n1676 1.733
R9424 VDD.n1685 VDD.n1678 1.733
R9425 VDD.n1737 VDD.n1728 1.733
R9426 VDD.n1737 VDD.n1730 1.733
R9427 VDD.n2107 VDD.n2106 1.723
R9428 VDD.n2212 VDD.n2211 1.723
R9429 VDD.n2338 VDD.n2337 1.723
R9430 VDD.n2443 VDD.n2442 1.723
R9431 VDD.n2515 VDD.n2514 1.723
R9432 VDD.n2506 VDD.n2505 1.723
R9433 VDD.n2562 VDD.n2561 1.723
R9434 VDD.n5155 VDD.n5154 1.723
R9435 VDD.n5164 VDD.n5163 1.723
R9436 VDD.n5223 VDD.n5221 1.723
R9437 VDD.n5248 VDD.n5238 1.723
R9438 VDD.n2644 VDD.n2634 1.723
R9439 VDD.n2636 VDD.n2635 1.723
R9440 VDD.n2668 VDD.n2667 1.723
R9441 VDD.n2659 VDD.n2658 1.723
R9442 VDD.n5110 VDD.n5109 1.723
R9443 VDD.n5090 VDD.n5089 1.723
R9444 VDD.n5047 VDD.n5046 1.723
R9445 VDD.n4942 VDD.n4941 1.723
R9446 VDD.n4816 VDD.n4815 1.723
R9447 VDD.n4711 VDD.n4710 1.723
R9448 VDD.n3046 VDD.n3045 1.719
R9449 VDD.n3069 VDD.n3062 1.719
R9450 VDD.n3185 VDD.n3176 1.719
R9451 VDD.n3178 VDD.n3177 1.719
R9452 VDD.n3283 VDD.n3282 1.719
R9453 VDD.n3306 VDD.n3299 1.719
R9454 VDD.n3422 VDD.n3413 1.719
R9455 VDD.n3415 VDD.n3414 1.719
R9456 VDD.n3521 VDD.n3520 1.719
R9457 VDD.n3544 VDD.n3537 1.719
R9458 VDD.n3660 VDD.n3651 1.719
R9459 VDD.n3653 VDD.n3652 1.719
R9460 VDD.n3758 VDD.n3757 1.719
R9461 VDD.n3781 VDD.n3774 1.719
R9462 VDD.n3897 VDD.n3888 1.719
R9463 VDD.n3890 VDD.n3889 1.719
R9464 VDD.n3996 VDD.n3995 1.719
R9465 VDD.n4019 VDD.n4012 1.719
R9466 VDD.n4135 VDD.n4126 1.719
R9467 VDD.n4128 VDD.n4127 1.719
R9468 VDD.n4233 VDD.n4232 1.719
R9469 VDD.n4256 VDD.n4249 1.719
R9470 VDD.n4372 VDD.n4363 1.719
R9471 VDD.n4365 VDD.n4364 1.719
R9472 VDD.n57 VDD.n56 1.715
R9473 VDD.n66 VDD.n65 1.715
R9474 VDD.n11422 VDD.n11421 1.715
R9475 VDD.n11224 VDD.n11223 1.715
R9476 VDD.n11933 VDD.n11932 1.715
R9477 VDD.n12288 VDD.n12287 1.715
R9478 VDD.n12297 VDD.n12296 1.715
R9479 VDD.n10222 VDD.n10221 1.659
R9480 VDD.n10230 VDD.n10229 1.659
R9481 VDD.n10105 VDD.n10104 1.659
R9482 VDD.n10113 VDD.n10112 1.659
R9483 VDD.n10569 VDD.n10568 1.659
R9484 VDD.n10577 VDD.n10576 1.659
R9485 VDD.n10451 VDD.n10450 1.659
R9486 VDD.n10459 VDD.n10458 1.659
R9487 VDD.n383 VDD.n382 1.6
R9488 VDD.n385 VDD.n384 1.6
R9489 VDD.n452 VDD.n451 1.6
R9490 VDD.n454 VDD.n453 1.6
R9491 VDD.n617 VDD.n616 1.6
R9492 VDD.n619 VDD.n618 1.6
R9493 VDD.n685 VDD.n684 1.6
R9494 VDD.n687 VDD.n686 1.6
R9495 VDD.n850 VDD.n849 1.6
R9496 VDD.n852 VDD.n851 1.6
R9497 VDD.n919 VDD.n918 1.6
R9498 VDD.n921 VDD.n920 1.6
R9499 VDD.n1084 VDD.n1083 1.6
R9500 VDD.n1086 VDD.n1085 1.6
R9501 VDD.n1152 VDD.n1151 1.6
R9502 VDD.n1154 VDD.n1153 1.6
R9503 VDD.n1317 VDD.n1316 1.6
R9504 VDD.n1319 VDD.n1318 1.6
R9505 VDD.n1386 VDD.n1385 1.6
R9506 VDD.n1388 VDD.n1387 1.6
R9507 VDD.n1551 VDD.n1550 1.6
R9508 VDD.n1553 VDD.n1552 1.6
R9509 VDD.n1619 VDD.n1618 1.6
R9510 VDD.n1621 VDD.n1620 1.6
R9511 VDD.n1784 VDD.n1783 1.6
R9512 VDD.n1786 VDD.n1785 1.6
R9513 VDD.n12131 VDD.n12130 1.551
R9514 VDD.n12036 VDD.n12035 1.551
R9515 VDD.n10899 VDD.n10898 1.551
R9516 VDD.n11085 VDD.n11084 1.551
R9517 VDD.n10863 VDD.n10862 1.551
R9518 VDD.n10780 VDD.n10779 1.551
R9519 VDD.n10691 VDD.n10690 1.551
R9520 VDD.n11668 VDD.n11667 1.551
R9521 VDD.n11852 VDD.n11851 1.551
R9522 VDD.n11581 VDD.n11580 1.551
R9523 VDD.n11550 VDD.n11549 1.551
R9524 VDD.n11464 VDD.n11463 1.551
R9525 VDD.n11363 VDD.n11362 1.551
R9526 VDD.n11269 VDD.n11268 1.551
R9527 VDD.n3055 VDD.n3046 1.528
R9528 VDD.n3062 VDD.n3061 1.528
R9529 VDD.n3176 VDD.n3175 1.528
R9530 VDD.n3185 VDD.n3178 1.528
R9531 VDD.n3292 VDD.n3283 1.528
R9532 VDD.n3299 VDD.n3298 1.528
R9533 VDD.n3413 VDD.n3412 1.528
R9534 VDD.n3422 VDD.n3415 1.528
R9535 VDD.n3530 VDD.n3521 1.528
R9536 VDD.n3537 VDD.n3536 1.528
R9537 VDD.n3651 VDD.n3650 1.528
R9538 VDD.n3660 VDD.n3653 1.528
R9539 VDD.n3767 VDD.n3758 1.528
R9540 VDD.n3774 VDD.n3773 1.528
R9541 VDD.n3888 VDD.n3887 1.528
R9542 VDD.n3897 VDD.n3890 1.528
R9543 VDD.n4005 VDD.n3996 1.528
R9544 VDD.n4012 VDD.n4011 1.528
R9545 VDD.n4126 VDD.n4125 1.528
R9546 VDD.n4135 VDD.n4128 1.528
R9547 VDD.n4242 VDD.n4233 1.528
R9548 VDD.n4249 VDD.n4248 1.528
R9549 VDD.n4363 VDD.n4362 1.528
R9550 VDD.n4372 VDD.n4365 1.528
R9551 VDD.n5614 VDD.n5612 1.505
R9552 VDD.n5620 VDD.n5619 1.505
R9553 VDD.n5975 VDD.n5973 1.505
R9554 VDD.n5981 VDD.n5980 1.505
R9555 VDD.n6337 VDD.n6335 1.505
R9556 VDD.n6343 VDD.n6342 1.505
R9557 VDD.n6699 VDD.n6697 1.505
R9558 VDD.n6705 VDD.n6704 1.505
R9559 VDD.n7061 VDD.n7059 1.505
R9560 VDD.n7067 VDD.n7066 1.505
R9561 VDD.n7423 VDD.n7421 1.505
R9562 VDD.n7429 VDD.n7428 1.505
R9563 VDD.n7785 VDD.n7783 1.505
R9564 VDD.n7791 VDD.n7790 1.505
R9565 VDD.n8147 VDD.n8145 1.505
R9566 VDD.n8153 VDD.n8152 1.505
R9567 VDD.n8509 VDD.n8507 1.505
R9568 VDD.n8515 VDD.n8514 1.505
R9569 VDD.n8871 VDD.n8869 1.505
R9570 VDD.n8877 VDD.n8876 1.505
R9571 VDD.n9233 VDD.n9231 1.505
R9572 VDD.n9239 VDD.n9238 1.505
R9573 VDD.n9595 VDD.n9593 1.505
R9574 VDD.n9601 VDD.n9600 1.505
R9575 VDD.n9957 VDD.n9955 1.505
R9576 VDD.n9963 VDD.n9962 1.505
R9577 VDD.n5126 VDD.n5125 1.5
R9578 VDD.n2528 VDD.n2527 1.5
R9579 VDD.n2590 VDD.n2589 1.5
R9580 VDD.n156 VDD.n155 1.5
R9581 VDD.n2690 VDD.n2689 1.5
R9582 VDD.n2755 VDD.n2754 1.5
R9583 VDD.n10873 VDD.n10872 1.5
R9584 VDD.n11644 VDD.n11643 1.5
R9585 VDD.n11183 VDD.n11106 1.49
R9586 VDD.n2769 VDD.n2768 1.489
R9587 VDD.n2780 VDD.n2779 1.488
R9588 VDD.n2781 VDD.n2780 1.488
R9589 VDD.n2768 VDD.n2767 1.488
R9590 VDD.n2086 VDD.n2079 1.476
R9591 VDD.n2247 VDD.n2240 1.476
R9592 VDD.n2317 VDD.n2310 1.476
R9593 VDD.n2478 VDD.n2471 1.476
R9594 VDD.n2586 VDD.n2577 1.476
R9595 VDD.n127 VDD.n120 1.476
R9596 VDD.n5183 VDD.n5182 1.476
R9597 VDD.n5288 VDD.n5287 1.476
R9598 VDD.n2667 VDD.n2660 1.476
R9599 VDD.n2740 VDD.n2732 1.476
R9600 VDD.n5089 VDD.n5088 1.476
R9601 VDD.n5099 VDD.n5097 1.476
R9602 VDD.n5082 VDD.n5075 1.476
R9603 VDD.n4921 VDD.n4914 1.476
R9604 VDD.n4851 VDD.n4844 1.476
R9605 VDD.n4690 VDD.n4683 1.476
R9606 VDD.n503 VDD.n494 1.466
R9607 VDD.n503 VDD.n496 1.466
R9608 VDD.n584 VDD.n575 1.466
R9609 VDD.n584 VDD.n577 1.466
R9610 VDD.n737 VDD.n727 1.466
R9611 VDD.n737 VDD.n729 1.466
R9612 VDD.n817 VDD.n808 1.466
R9613 VDD.n817 VDD.n810 1.466
R9614 VDD.n970 VDD.n961 1.466
R9615 VDD.n970 VDD.n963 1.466
R9616 VDD.n1051 VDD.n1042 1.466
R9617 VDD.n1051 VDD.n1044 1.466
R9618 VDD.n1204 VDD.n1194 1.466
R9619 VDD.n1204 VDD.n1196 1.466
R9620 VDD.n1284 VDD.n1275 1.466
R9621 VDD.n1284 VDD.n1277 1.466
R9622 VDD.n1437 VDD.n1428 1.466
R9623 VDD.n1437 VDD.n1430 1.466
R9624 VDD.n1518 VDD.n1509 1.466
R9625 VDD.n1518 VDD.n1511 1.466
R9626 VDD.n1671 VDD.n1661 1.466
R9627 VDD.n1671 VDD.n1663 1.466
R9628 VDD.n1751 VDD.n1742 1.466
R9629 VDD.n1751 VDD.n1744 1.466
R9630 VDD.n10437 VDD.n10436 1.439
R9631 VDD.n10401 VDD.n10399 1.439
R9632 VDD.n10374 VDD.n10372 1.439
R9633 VDD.n10357 VDD.n10355 1.439
R9634 VDD.n10321 VDD.n10316 1.422
R9635 VDD.n10259 VDD.n10253 1.422
R9636 VDD.n10202 VDD.n10197 1.422
R9637 VDD.n10142 VDD.n10137 1.422
R9638 VDD.n10668 VDD.n10663 1.422
R9639 VDD.n10606 VDD.n10600 1.422
R9640 VDD.n10548 VDD.n10543 1.422
R9641 VDD.n10488 VDD.n10483 1.422
R9642 VDD.n12149 VDD.n12144 1.357
R9643 VDD.n12029 VDD.n12024 1.357
R9644 VDD.n10889 VDD.n10884 1.357
R9645 VDD.n10917 VDD.n10912 1.357
R9646 VDD.n10777 VDD.n10772 1.357
R9647 VDD.n10715 VDD.n10710 1.357
R9648 VDD.n11658 VDD.n11653 1.357
R9649 VDD.n11685 VDD.n11680 1.357
R9650 VDD.n11547 VDD.n11542 1.357
R9651 VDD.n11485 VDD.n11480 1.357
R9652 VDD.n11380 VDD.n11375 1.357
R9653 VDD.n11262 VDD.n11257 1.357
R9654 VDD.n10431 VDD.n10430 1.355
R9655 VDD.n10405 VDD.n10404 1.355
R9656 VDD.n10378 VDD.n10377 1.355
R9657 VDD.n10349 VDD.n10348 1.355
R9658 VDD.n3055 VDD.n3048 1.337
R9659 VDD.n3060 VDD.n3059 1.337
R9660 VDD.n3164 VDD.n3163 1.337
R9661 VDD.n3199 VDD.n3190 1.337
R9662 VDD.n3292 VDD.n3285 1.337
R9663 VDD.n3297 VDD.n3296 1.337
R9664 VDD.n3401 VDD.n3400 1.337
R9665 VDD.n3436 VDD.n3427 1.337
R9666 VDD.n3530 VDD.n3523 1.337
R9667 VDD.n3535 VDD.n3534 1.337
R9668 VDD.n3639 VDD.n3638 1.337
R9669 VDD.n3674 VDD.n3665 1.337
R9670 VDD.n3767 VDD.n3760 1.337
R9671 VDD.n3772 VDD.n3771 1.337
R9672 VDD.n3876 VDD.n3875 1.337
R9673 VDD.n3911 VDD.n3902 1.337
R9674 VDD.n4005 VDD.n3998 1.337
R9675 VDD.n4010 VDD.n4009 1.337
R9676 VDD.n4114 VDD.n4113 1.337
R9677 VDD.n4149 VDD.n4140 1.337
R9678 VDD.n4242 VDD.n4235 1.337
R9679 VDD.n4247 VDD.n4246 1.337
R9680 VDD.n4351 VDD.n4350 1.337
R9681 VDD.n4386 VDD.n4377 1.337
R9682 VDD.n466 VDD.n465 1.333
R9683 VDD.n468 VDD.n467 1.333
R9684 VDD.n603 VDD.n602 1.333
R9685 VDD.n605 VDD.n604 1.333
R9686 VDD.n699 VDD.n698 1.333
R9687 VDD.n701 VDD.n700 1.333
R9688 VDD.n836 VDD.n835 1.333
R9689 VDD.n838 VDD.n837 1.333
R9690 VDD.n933 VDD.n932 1.333
R9691 VDD.n935 VDD.n934 1.333
R9692 VDD.n1070 VDD.n1069 1.333
R9693 VDD.n1072 VDD.n1071 1.333
R9694 VDD.n1166 VDD.n1165 1.333
R9695 VDD.n1168 VDD.n1167 1.333
R9696 VDD.n1303 VDD.n1302 1.333
R9697 VDD.n1305 VDD.n1304 1.333
R9698 VDD.n1400 VDD.n1399 1.333
R9699 VDD.n1402 VDD.n1401 1.333
R9700 VDD.n1537 VDD.n1536 1.333
R9701 VDD.n1539 VDD.n1538 1.333
R9702 VDD.n1633 VDD.n1632 1.333
R9703 VDD.n1635 VDD.n1634 1.333
R9704 VDD.n1770 VDD.n1769 1.333
R9705 VDD.n1772 VDD.n1771 1.333
R9706 VDD.n5 VDD.n3 1.248
R9707 VDD.n12236 VDD.n12234 1.248
R9708 VDD.n2121 VDD.n2120 1.23
R9709 VDD.n2198 VDD.n2197 1.23
R9710 VDD.n2352 VDD.n2351 1.23
R9711 VDD.n2429 VDD.n2428 1.23
R9712 VDD.n2495 VDD.n2494 1.23
R9713 VDD.n2486 VDD.n2485 1.23
R9714 VDD.n2573 VDD.n2572 1.23
R9715 VDD.n5173 VDD.n5172 1.23
R9716 VDD.n5240 VDD.n5239 1.23
R9717 VDD.n2746 VDD.n2745 1.23
R9718 VDD.n5033 VDD.n5032 1.23
R9719 VDD.n4956 VDD.n4955 1.23
R9720 VDD.n4802 VDD.n4801 1.23
R9721 VDD.n4725 VDD.n4724 1.23
R9722 VDD.n10883 VDD.n10881 1.211
R9723 VDD.n10709 VDD.n10707 1.211
R9724 VDD.n11652 VDD.n11650 1.211
R9725 VDD.n11479 VDD.n11477 1.211
R9726 VDD.n4627 VDD.n4626 1.21
R9727 VDD.n489 VDD.n480 1.2
R9728 VDD.n489 VDD.n482 1.2
R9729 VDD.n598 VDD.n589 1.2
R9730 VDD.n598 VDD.n591 1.2
R9731 VDD.n722 VDD.n713 1.2
R9732 VDD.n722 VDD.n715 1.2
R9733 VDD.n831 VDD.n822 1.2
R9734 VDD.n831 VDD.n824 1.2
R9735 VDD.n956 VDD.n947 1.2
R9736 VDD.n956 VDD.n949 1.2
R9737 VDD.n1065 VDD.n1056 1.2
R9738 VDD.n1065 VDD.n1058 1.2
R9739 VDD.n1189 VDD.n1180 1.2
R9740 VDD.n1189 VDD.n1182 1.2
R9741 VDD.n1298 VDD.n1289 1.2
R9742 VDD.n1298 VDD.n1291 1.2
R9743 VDD.n1423 VDD.n1414 1.2
R9744 VDD.n1423 VDD.n1416 1.2
R9745 VDD.n1532 VDD.n1523 1.2
R9746 VDD.n1532 VDD.n1525 1.2
R9747 VDD.n1656 VDD.n1647 1.2
R9748 VDD.n1656 VDD.n1649 1.2
R9749 VDD.n1765 VDD.n1756 1.2
R9750 VDD.n1765 VDD.n1758 1.2
R9751 VDD.n6030 VDD.n5668 1.182
R9752 VDD.n12119 VDD.n12118 1.163
R9753 VDD.n12049 VDD.n12048 1.163
R9754 VDD.n10906 VDD.n10905 1.163
R9755 VDD.n10908 VDD.n10907 1.163
R9756 VDD.n10911 VDD.n10910 1.163
R9757 VDD.n11061 VDD.n11060 1.163
R9758 VDD.n10983 VDD.n10982 1.163
R9759 VDD.n11098 VDD.n11097 1.163
R9760 VDD.n10847 VDD.n10846 1.163
R9761 VDD.n10779 VDD.n10778 1.163
R9762 VDD.n11674 VDD.n11673 1.163
R9763 VDD.n11676 VDD.n11675 1.163
R9764 VDD.n11679 VDD.n11678 1.163
R9765 VDD.n11827 VDD.n11826 1.163
R9766 VDD.n11752 VDD.n11751 1.163
R9767 VDD.n11873 VDD.n11872 1.163
R9768 VDD.n11628 VDD.n11627 1.163
R9769 VDD.n11549 VDD.n11548 1.163
R9770 VDD.n11351 VDD.n11350 1.163
R9771 VDD.n11281 VDD.n11280 1.163
R9772 VDD.n3041 VDD.n3032 1.146
R9773 VDD.n3076 VDD.n3075 1.146
R9774 VDD.n3162 VDD.n3161 1.146
R9775 VDD.n3199 VDD.n3192 1.146
R9776 VDD.n3278 VDD.n3269 1.146
R9777 VDD.n3313 VDD.n3312 1.146
R9778 VDD.n3399 VDD.n3398 1.146
R9779 VDD.n3436 VDD.n3429 1.146
R9780 VDD.n3516 VDD.n3507 1.146
R9781 VDD.n3551 VDD.n3550 1.146
R9782 VDD.n3637 VDD.n3636 1.146
R9783 VDD.n3674 VDD.n3667 1.146
R9784 VDD.n3753 VDD.n3744 1.146
R9785 VDD.n3788 VDD.n3787 1.146
R9786 VDD.n3874 VDD.n3873 1.146
R9787 VDD.n3911 VDD.n3904 1.146
R9788 VDD.n3991 VDD.n3982 1.146
R9789 VDD.n4026 VDD.n4025 1.146
R9790 VDD.n4112 VDD.n4111 1.146
R9791 VDD.n4149 VDD.n4142 1.146
R9792 VDD.n4228 VDD.n4219 1.146
R9793 VDD.n4263 VDD.n4262 1.146
R9794 VDD.n4349 VDD.n4348 1.146
R9795 VDD.n4386 VDD.n4379 1.146
R9796 VDD.n12078 VDD.n12077 1.145
R9797 VDD.n11033 VDD.n11032 1.145
R9798 VDD.n10741 VDD.n10740 1.145
R9799 VDD.n10816 VDD.n10815 1.145
R9800 VDD.n10941 VDD.n10940 1.145
R9801 VDD.n11800 VDD.n11799 1.145
R9802 VDD.n11512 VDD.n11511 1.145
R9803 VDD.n12098 VDD.n12097 1.145
R9804 VDD.n11309 VDD.n11308 1.145
R9805 VDD.n10432 VDD.n10431 1.144
R9806 VDD.n10406 VDD.n10405 1.142
R9807 VDD.n10379 VDD.n10378 1.142
R9808 VDD.n14 VDD.n13 1.141
R9809 VDD.n12245 VDD.n12244 1.141
R9810 VDD.n21 VDD.n20 1.138
R9811 VDD.n12324 VDD.n12323 1.138
R9812 VDD.n90 VDD.n89 1.137
R9813 VDD.n18 VDD.n17 1.137
R9814 VDD.n5583 VDD.n5582 1.137
R9815 VDD.n5591 VDD.n5590 1.137
R9816 VDD.n5541 VDD.n5540 1.137
R9817 VDD.n5434 VDD.n5433 1.137
R9818 VDD.n5406 VDD.n5405 1.137
R9819 VDD.n5392 VDD.n5391 1.137
R9820 VDD.n5398 VDD.n5397 1.137
R9821 VDD.n5415 VDD.n5414 1.137
R9822 VDD.n5430 VDD.n5429 1.137
R9823 VDD.n5423 VDD.n5422 1.137
R9824 VDD.n5441 VDD.n5440 1.137
R9825 VDD.n5451 VDD.n5450 1.137
R9826 VDD.n5537 VDD.n5536 1.137
R9827 VDD.n5460 VDD.n5459 1.137
R9828 VDD.n5530 VDD.n5529 1.137
R9829 VDD.n5548 VDD.n5547 1.137
R9830 VDD.n5558 VDD.n5557 1.137
R9831 VDD.n5564 VDD.n5563 1.137
R9832 VDD.n5579 VDD.n5578 1.137
R9833 VDD.n5572 VDD.n5571 1.137
R9834 VDD.n5668 VDD.n5667 1.137
R9835 VDD.n5944 VDD.n5943 1.137
R9836 VDD.n5952 VDD.n5951 1.137
R9837 VDD.n5902 VDD.n5901 1.137
R9838 VDD.n5795 VDD.n5794 1.137
R9839 VDD.n5767 VDD.n5766 1.137
R9840 VDD.n5753 VDD.n5752 1.137
R9841 VDD.n5759 VDD.n5758 1.137
R9842 VDD.n5776 VDD.n5775 1.137
R9843 VDD.n5791 VDD.n5790 1.137
R9844 VDD.n5784 VDD.n5783 1.137
R9845 VDD.n5802 VDD.n5801 1.137
R9846 VDD.n5812 VDD.n5811 1.137
R9847 VDD.n5898 VDD.n5897 1.137
R9848 VDD.n5821 VDD.n5820 1.137
R9849 VDD.n5891 VDD.n5890 1.137
R9850 VDD.n5909 VDD.n5908 1.137
R9851 VDD.n5919 VDD.n5918 1.137
R9852 VDD.n5925 VDD.n5924 1.137
R9853 VDD.n5940 VDD.n5939 1.137
R9854 VDD.n5933 VDD.n5932 1.137
R9855 VDD.n6029 VDD.n6028 1.137
R9856 VDD.n6306 VDD.n6305 1.137
R9857 VDD.n6314 VDD.n6313 1.137
R9858 VDD.n6264 VDD.n6263 1.137
R9859 VDD.n6157 VDD.n6156 1.137
R9860 VDD.n6129 VDD.n6128 1.137
R9861 VDD.n6115 VDD.n6114 1.137
R9862 VDD.n6121 VDD.n6120 1.137
R9863 VDD.n6138 VDD.n6137 1.137
R9864 VDD.n6153 VDD.n6152 1.137
R9865 VDD.n6146 VDD.n6145 1.137
R9866 VDD.n6164 VDD.n6163 1.137
R9867 VDD.n6174 VDD.n6173 1.137
R9868 VDD.n6260 VDD.n6259 1.137
R9869 VDD.n6183 VDD.n6182 1.137
R9870 VDD.n6253 VDD.n6252 1.137
R9871 VDD.n6271 VDD.n6270 1.137
R9872 VDD.n6281 VDD.n6280 1.137
R9873 VDD.n6287 VDD.n6286 1.137
R9874 VDD.n6302 VDD.n6301 1.137
R9875 VDD.n6295 VDD.n6294 1.137
R9876 VDD.n6391 VDD.n6390 1.137
R9877 VDD.n6668 VDD.n6667 1.137
R9878 VDD.n6676 VDD.n6675 1.137
R9879 VDD.n6626 VDD.n6625 1.137
R9880 VDD.n6519 VDD.n6518 1.137
R9881 VDD.n6491 VDD.n6490 1.137
R9882 VDD.n6477 VDD.n6476 1.137
R9883 VDD.n6483 VDD.n6482 1.137
R9884 VDD.n6500 VDD.n6499 1.137
R9885 VDD.n6515 VDD.n6514 1.137
R9886 VDD.n6508 VDD.n6507 1.137
R9887 VDD.n6526 VDD.n6525 1.137
R9888 VDD.n6536 VDD.n6535 1.137
R9889 VDD.n6622 VDD.n6621 1.137
R9890 VDD.n6545 VDD.n6544 1.137
R9891 VDD.n6615 VDD.n6614 1.137
R9892 VDD.n6633 VDD.n6632 1.137
R9893 VDD.n6643 VDD.n6642 1.137
R9894 VDD.n6649 VDD.n6648 1.137
R9895 VDD.n6664 VDD.n6663 1.137
R9896 VDD.n6657 VDD.n6656 1.137
R9897 VDD.n6753 VDD.n6752 1.137
R9898 VDD.n7030 VDD.n7029 1.137
R9899 VDD.n7038 VDD.n7037 1.137
R9900 VDD.n6988 VDD.n6987 1.137
R9901 VDD.n6881 VDD.n6880 1.137
R9902 VDD.n6853 VDD.n6852 1.137
R9903 VDD.n6839 VDD.n6838 1.137
R9904 VDD.n6845 VDD.n6844 1.137
R9905 VDD.n6862 VDD.n6861 1.137
R9906 VDD.n6877 VDD.n6876 1.137
R9907 VDD.n6870 VDD.n6869 1.137
R9908 VDD.n6888 VDD.n6887 1.137
R9909 VDD.n6898 VDD.n6897 1.137
R9910 VDD.n6984 VDD.n6983 1.137
R9911 VDD.n6907 VDD.n6906 1.137
R9912 VDD.n6977 VDD.n6976 1.137
R9913 VDD.n6995 VDD.n6994 1.137
R9914 VDD.n7005 VDD.n7004 1.137
R9915 VDD.n7011 VDD.n7010 1.137
R9916 VDD.n7026 VDD.n7025 1.137
R9917 VDD.n7019 VDD.n7018 1.137
R9918 VDD.n7115 VDD.n7114 1.137
R9919 VDD.n7392 VDD.n7391 1.137
R9920 VDD.n7400 VDD.n7399 1.137
R9921 VDD.n7350 VDD.n7349 1.137
R9922 VDD.n7243 VDD.n7242 1.137
R9923 VDD.n7215 VDD.n7214 1.137
R9924 VDD.n7201 VDD.n7200 1.137
R9925 VDD.n7207 VDD.n7206 1.137
R9926 VDD.n7224 VDD.n7223 1.137
R9927 VDD.n7239 VDD.n7238 1.137
R9928 VDD.n7232 VDD.n7231 1.137
R9929 VDD.n7250 VDD.n7249 1.137
R9930 VDD.n7260 VDD.n7259 1.137
R9931 VDD.n7346 VDD.n7345 1.137
R9932 VDD.n7269 VDD.n7268 1.137
R9933 VDD.n7339 VDD.n7338 1.137
R9934 VDD.n7357 VDD.n7356 1.137
R9935 VDD.n7367 VDD.n7366 1.137
R9936 VDD.n7373 VDD.n7372 1.137
R9937 VDD.n7388 VDD.n7387 1.137
R9938 VDD.n7381 VDD.n7380 1.137
R9939 VDD.n7477 VDD.n7476 1.137
R9940 VDD.n7754 VDD.n7753 1.137
R9941 VDD.n7762 VDD.n7761 1.137
R9942 VDD.n7712 VDD.n7711 1.137
R9943 VDD.n7605 VDD.n7604 1.137
R9944 VDD.n7577 VDD.n7576 1.137
R9945 VDD.n7563 VDD.n7562 1.137
R9946 VDD.n7569 VDD.n7568 1.137
R9947 VDD.n7586 VDD.n7585 1.137
R9948 VDD.n7601 VDD.n7600 1.137
R9949 VDD.n7594 VDD.n7593 1.137
R9950 VDD.n7612 VDD.n7611 1.137
R9951 VDD.n7622 VDD.n7621 1.137
R9952 VDD.n7708 VDD.n7707 1.137
R9953 VDD.n7631 VDD.n7630 1.137
R9954 VDD.n7701 VDD.n7700 1.137
R9955 VDD.n7719 VDD.n7718 1.137
R9956 VDD.n7729 VDD.n7728 1.137
R9957 VDD.n7735 VDD.n7734 1.137
R9958 VDD.n7750 VDD.n7749 1.137
R9959 VDD.n7743 VDD.n7742 1.137
R9960 VDD.n7839 VDD.n7838 1.137
R9961 VDD.n8116 VDD.n8115 1.137
R9962 VDD.n8124 VDD.n8123 1.137
R9963 VDD.n8074 VDD.n8073 1.137
R9964 VDD.n7967 VDD.n7966 1.137
R9965 VDD.n7939 VDD.n7938 1.137
R9966 VDD.n7925 VDD.n7924 1.137
R9967 VDD.n7931 VDD.n7930 1.137
R9968 VDD.n7948 VDD.n7947 1.137
R9969 VDD.n7963 VDD.n7962 1.137
R9970 VDD.n7956 VDD.n7955 1.137
R9971 VDD.n7974 VDD.n7973 1.137
R9972 VDD.n7984 VDD.n7983 1.137
R9973 VDD.n8070 VDD.n8069 1.137
R9974 VDD.n7993 VDD.n7992 1.137
R9975 VDD.n8063 VDD.n8062 1.137
R9976 VDD.n8081 VDD.n8080 1.137
R9977 VDD.n8091 VDD.n8090 1.137
R9978 VDD.n8097 VDD.n8096 1.137
R9979 VDD.n8112 VDD.n8111 1.137
R9980 VDD.n8105 VDD.n8104 1.137
R9981 VDD.n8201 VDD.n8200 1.137
R9982 VDD.n8478 VDD.n8477 1.137
R9983 VDD.n8486 VDD.n8485 1.137
R9984 VDD.n8436 VDD.n8435 1.137
R9985 VDD.n8329 VDD.n8328 1.137
R9986 VDD.n8301 VDD.n8300 1.137
R9987 VDD.n8287 VDD.n8286 1.137
R9988 VDD.n8293 VDD.n8292 1.137
R9989 VDD.n8310 VDD.n8309 1.137
R9990 VDD.n8325 VDD.n8324 1.137
R9991 VDD.n8318 VDD.n8317 1.137
R9992 VDD.n8336 VDD.n8335 1.137
R9993 VDD.n8346 VDD.n8345 1.137
R9994 VDD.n8432 VDD.n8431 1.137
R9995 VDD.n8355 VDD.n8354 1.137
R9996 VDD.n8425 VDD.n8424 1.137
R9997 VDD.n8443 VDD.n8442 1.137
R9998 VDD.n8453 VDD.n8452 1.137
R9999 VDD.n8459 VDD.n8458 1.137
R10000 VDD.n8474 VDD.n8473 1.137
R10001 VDD.n8467 VDD.n8466 1.137
R10002 VDD.n8563 VDD.n8562 1.137
R10003 VDD.n8840 VDD.n8839 1.137
R10004 VDD.n8848 VDD.n8847 1.137
R10005 VDD.n8798 VDD.n8797 1.137
R10006 VDD.n8691 VDD.n8690 1.137
R10007 VDD.n8663 VDD.n8662 1.137
R10008 VDD.n8649 VDD.n8648 1.137
R10009 VDD.n8655 VDD.n8654 1.137
R10010 VDD.n8672 VDD.n8671 1.137
R10011 VDD.n8687 VDD.n8686 1.137
R10012 VDD.n8680 VDD.n8679 1.137
R10013 VDD.n8698 VDD.n8697 1.137
R10014 VDD.n8708 VDD.n8707 1.137
R10015 VDD.n8794 VDD.n8793 1.137
R10016 VDD.n8717 VDD.n8716 1.137
R10017 VDD.n8787 VDD.n8786 1.137
R10018 VDD.n8805 VDD.n8804 1.137
R10019 VDD.n8815 VDD.n8814 1.137
R10020 VDD.n8821 VDD.n8820 1.137
R10021 VDD.n8836 VDD.n8835 1.137
R10022 VDD.n8829 VDD.n8828 1.137
R10023 VDD.n8925 VDD.n8924 1.137
R10024 VDD.n9202 VDD.n9201 1.137
R10025 VDD.n9210 VDD.n9209 1.137
R10026 VDD.n9160 VDD.n9159 1.137
R10027 VDD.n9053 VDD.n9052 1.137
R10028 VDD.n9025 VDD.n9024 1.137
R10029 VDD.n9011 VDD.n9010 1.137
R10030 VDD.n9017 VDD.n9016 1.137
R10031 VDD.n9034 VDD.n9033 1.137
R10032 VDD.n9049 VDD.n9048 1.137
R10033 VDD.n9042 VDD.n9041 1.137
R10034 VDD.n9060 VDD.n9059 1.137
R10035 VDD.n9070 VDD.n9069 1.137
R10036 VDD.n9156 VDD.n9155 1.137
R10037 VDD.n9079 VDD.n9078 1.137
R10038 VDD.n9149 VDD.n9148 1.137
R10039 VDD.n9167 VDD.n9166 1.137
R10040 VDD.n9177 VDD.n9176 1.137
R10041 VDD.n9183 VDD.n9182 1.137
R10042 VDD.n9198 VDD.n9197 1.137
R10043 VDD.n9191 VDD.n9190 1.137
R10044 VDD.n9287 VDD.n9286 1.137
R10045 VDD.n9564 VDD.n9563 1.137
R10046 VDD.n9572 VDD.n9571 1.137
R10047 VDD.n9522 VDD.n9521 1.137
R10048 VDD.n9415 VDD.n9414 1.137
R10049 VDD.n9387 VDD.n9386 1.137
R10050 VDD.n9373 VDD.n9372 1.137
R10051 VDD.n9379 VDD.n9378 1.137
R10052 VDD.n9396 VDD.n9395 1.137
R10053 VDD.n9411 VDD.n9410 1.137
R10054 VDD.n9404 VDD.n9403 1.137
R10055 VDD.n9422 VDD.n9421 1.137
R10056 VDD.n9432 VDD.n9431 1.137
R10057 VDD.n9518 VDD.n9517 1.137
R10058 VDD.n9441 VDD.n9440 1.137
R10059 VDD.n9511 VDD.n9510 1.137
R10060 VDD.n9529 VDD.n9528 1.137
R10061 VDD.n9539 VDD.n9538 1.137
R10062 VDD.n9545 VDD.n9544 1.137
R10063 VDD.n9560 VDD.n9559 1.137
R10064 VDD.n9553 VDD.n9552 1.137
R10065 VDD.n9649 VDD.n9648 1.137
R10066 VDD.n9926 VDD.n9925 1.137
R10067 VDD.n9934 VDD.n9933 1.137
R10068 VDD.n9884 VDD.n9883 1.137
R10069 VDD.n9777 VDD.n9776 1.137
R10070 VDD.n9749 VDD.n9748 1.137
R10071 VDD.n9735 VDD.n9734 1.137
R10072 VDD.n9741 VDD.n9740 1.137
R10073 VDD.n9758 VDD.n9757 1.137
R10074 VDD.n9773 VDD.n9772 1.137
R10075 VDD.n9766 VDD.n9765 1.137
R10076 VDD.n9784 VDD.n9783 1.137
R10077 VDD.n9794 VDD.n9793 1.137
R10078 VDD.n9880 VDD.n9879 1.137
R10079 VDD.n9803 VDD.n9802 1.137
R10080 VDD.n9873 VDD.n9872 1.137
R10081 VDD.n9891 VDD.n9890 1.137
R10082 VDD.n9901 VDD.n9900 1.137
R10083 VDD.n9907 VDD.n9906 1.137
R10084 VDD.n9922 VDD.n9921 1.137
R10085 VDD.n9915 VDD.n9914 1.137
R10086 VDD.n10011 VDD.n10010 1.137
R10087 VDD.n10443 VDD.n10442 1.137
R10088 VDD.n10425 VDD.n10424 1.137
R10089 VDD.n10438 VDD.n10437 1.137
R10090 VDD.n10402 VDD.n10401 1.137
R10091 VDD.n10412 VDD.n10411 1.137
R10092 VDD.n10417 VDD.n10416 1.137
R10093 VDD.n10375 VDD.n10374 1.137
R10094 VDD.n10385 VDD.n10384 1.137
R10095 VDD.n10390 VDD.n10389 1.137
R10096 VDD.n10358 VDD.n10357 1.137
R10097 VDD.n10350 VDD.n10349 1.137
R10098 VDD.n10344 VDD.n10343 1.137
R10099 VDD.n10363 VDD.n10362 1.137
R10100 VDD.n12321 VDD.n12320 1.137
R10101 VDD.n12252 VDD.n12251 1.137
R10102 VDD.n10433 VDD.n10432 1.137
R10103 VDD.n10352 VDD.n10351 1.136
R10104 VDD.n10446 VDD.n10445 1.136
R10105 VDD.n10366 VDD.n10365 1.136
R10106 VDD.n10393 VDD.n10392 1.136
R10107 VDD.n10420 VDD.n10419 1.136
R10108 VDD.n93 VDD.n92 1.135
R10109 VDD.n5322 VDD.n5321 1.129
R10110 VDD.n5335 VDD.n5334 1.129
R10111 VDD.n5338 VDD.n5337 1.129
R10112 VDD.n5683 VDD.n5682 1.129
R10113 VDD.n5696 VDD.n5695 1.129
R10114 VDD.n5699 VDD.n5698 1.129
R10115 VDD.n6045 VDD.n6044 1.129
R10116 VDD.n6058 VDD.n6057 1.129
R10117 VDD.n6061 VDD.n6060 1.129
R10118 VDD.n6407 VDD.n6406 1.129
R10119 VDD.n6420 VDD.n6419 1.129
R10120 VDD.n6423 VDD.n6422 1.129
R10121 VDD.n6769 VDD.n6768 1.129
R10122 VDD.n6782 VDD.n6781 1.129
R10123 VDD.n6785 VDD.n6784 1.129
R10124 VDD.n7131 VDD.n7130 1.129
R10125 VDD.n7144 VDD.n7143 1.129
R10126 VDD.n7147 VDD.n7146 1.129
R10127 VDD.n7493 VDD.n7492 1.129
R10128 VDD.n7506 VDD.n7505 1.129
R10129 VDD.n7509 VDD.n7508 1.129
R10130 VDD.n7855 VDD.n7854 1.129
R10131 VDD.n7868 VDD.n7867 1.129
R10132 VDD.n7871 VDD.n7870 1.129
R10133 VDD.n8217 VDD.n8216 1.129
R10134 VDD.n8230 VDD.n8229 1.129
R10135 VDD.n8233 VDD.n8232 1.129
R10136 VDD.n8579 VDD.n8578 1.129
R10137 VDD.n8592 VDD.n8591 1.129
R10138 VDD.n8595 VDD.n8594 1.129
R10139 VDD.n8941 VDD.n8940 1.129
R10140 VDD.n8954 VDD.n8953 1.129
R10141 VDD.n8957 VDD.n8956 1.129
R10142 VDD.n9303 VDD.n9302 1.129
R10143 VDD.n9316 VDD.n9315 1.129
R10144 VDD.n9319 VDD.n9318 1.129
R10145 VDD.n9665 VDD.n9664 1.129
R10146 VDD.n9678 VDD.n9677 1.129
R10147 VDD.n9681 VDD.n9680 1.129
R10148 VDD.n5297 VDD.n5296 1.125
R10149 VDD.n11183 VDD.n11088 1.11
R10150 VDD.n11940 VDD.n11855 1.11
R10151 VDD.n11940 VDD.n11939 1.101
R10152 VDD.n11183 VDD.n11182 1.101
R10153 VDD.n6030 VDD.n6029 1.09
R10154 VDD.n6392 VDD.n6391 1.09
R10155 VDD.n6754 VDD.n6753 1.09
R10156 VDD.n7116 VDD.n7115 1.09
R10157 VDD.n7478 VDD.n7477 1.09
R10158 VDD.n7840 VDD.n7839 1.09
R10159 VDD.n8202 VDD.n8201 1.09
R10160 VDD.n8564 VDD.n8563 1.09
R10161 VDD.n8926 VDD.n8925 1.09
R10162 VDD.n9288 VDD.n9287 1.09
R10163 VDD.n9650 VDD.n9649 1.09
R10164 VDD.n10012 VDD.n10011 1.09
R10165 VDD VDD.n12326 1.089
R10166 VDD.n5307 VDD.n94 1.074
R10167 VDD.n480 VDD.n479 1.066
R10168 VDD.n482 VDD.n481 1.066
R10169 VDD.n589 VDD.n588 1.066
R10170 VDD.n591 VDD.n590 1.066
R10171 VDD.n713 VDD.n712 1.066
R10172 VDD.n715 VDD.n714 1.066
R10173 VDD.n822 VDD.n821 1.066
R10174 VDD.n824 VDD.n823 1.066
R10175 VDD.n947 VDD.n946 1.066
R10176 VDD.n949 VDD.n948 1.066
R10177 VDD.n1056 VDD.n1055 1.066
R10178 VDD.n1058 VDD.n1057 1.066
R10179 VDD.n1180 VDD.n1179 1.066
R10180 VDD.n1182 VDD.n1181 1.066
R10181 VDD.n1289 VDD.n1288 1.066
R10182 VDD.n1291 VDD.n1290 1.066
R10183 VDD.n1414 VDD.n1413 1.066
R10184 VDD.n1416 VDD.n1415 1.066
R10185 VDD.n1523 VDD.n1522 1.066
R10186 VDD.n1525 VDD.n1524 1.066
R10187 VDD.n1647 VDD.n1646 1.066
R10188 VDD.n1649 VDD.n1648 1.066
R10189 VDD.n1756 VDD.n1755 1.066
R10190 VDD.n1758 VDD.n1757 1.066
R10191 VDD.n10689 VDD.n10012 1.047
R10192 VDD.n13 VDD.n12 1.043
R10193 VDD.n12244 VDD.n12243 1.043
R10194 VDD.n5529 VDD.n5528 1.042
R10195 VDD.n5890 VDD.n5889 1.042
R10196 VDD.n6252 VDD.n6251 1.042
R10197 VDD.n6614 VDD.n6613 1.042
R10198 VDD.n6976 VDD.n6975 1.042
R10199 VDD.n7338 VDD.n7337 1.042
R10200 VDD.n7700 VDD.n7699 1.042
R10201 VDD.n8062 VDD.n8061 1.042
R10202 VDD.n8424 VDD.n8423 1.042
R10203 VDD.n8786 VDD.n8785 1.042
R10204 VDD.n9148 VDD.n9147 1.042
R10205 VDD.n9510 VDD.n9509 1.042
R10206 VDD.n9872 VDD.n9871 1.042
R10207 VDD.n11816 VDD.n11815 1.009
R10208 VDD.n11524 VDD.n11523 1.009
R10209 VDD.n11297 VDD.n11296 1.009
R10210 VDD.n88 VDD.n87 1.008
R10211 VDD.n366 VDD.n365 1.003
R10212 VDD.n2008 VDD.n2007 1.003
R10213 VDD.n2817 VDD.n2816 1.003
R10214 VDD.n241 VDD.n240 1.003
R10215 VDD.n4614 VDD.n4613 1.002
R10216 VDD.n2949 VDD.n2948 1.002
R10217 VDD.n2031 VDD.n197 0.984
R10218 VDD.n2072 VDD.n2065 0.984
R10219 VDD.n2261 VDD.n2254 0.984
R10220 VDD.n2303 VDD.n2296 0.984
R10221 VDD.n2494 VDD.n2487 0.984
R10222 VDD.n2560 VDD.n2553 0.984
R10223 VDD.n2660 VDD.n2659 0.984
R10224 VDD.n2721 VDD.n2714 0.984
R10225 VDD.n2714 VDD.n2713 0.984
R10226 VDD.n5097 VDD.n5090 0.984
R10227 VDD.n4907 VDD.n4900 0.984
R10228 VDD.n4865 VDD.n4858 0.984
R10229 VDD.n4676 VDD.n4669 0.984
R10230 VDD.n4635 VDD.n2766 0.984
R10231 VDD.n29 VDD.n24 0.969
R10232 VDD.n35 VDD.n31 0.969
R10233 VDD.n12220 VDD.n12215 0.969
R10234 VDD.n12162 VDD.n12156 0.969
R10235 VDD.n12017 VDD.n12011 0.969
R10236 VDD.n11958 VDD.n11953 0.969
R10237 VDD.n10881 VDD.n10875 0.969
R10238 VDD.n11083 VDD.n11077 0.969
R10239 VDD.n11086 VDD.n11083 0.969
R10240 VDD.n11133 VDD.n11120 0.969
R10241 VDD.n11096 VDD.n11090 0.969
R10242 VDD.n10871 VDD.n10863 0.969
R10243 VDD.n10870 VDD.n10864 0.969
R10244 VDD.n10700 VDD.n10699 0.969
R10245 VDD.n10698 VDD.n10697 0.969
R10246 VDD.n10707 VDD.n10701 0.969
R10247 VDD.n11850 VDD.n11845 0.969
R10248 VDD.n11853 VDD.n11850 0.969
R10249 VDD.n11863 VDD.n11857 0.969
R10250 VDD.n11871 VDD.n11865 0.969
R10251 VDD.n11588 VDD.n11581 0.969
R10252 VDD.n11587 VDD.n11582 0.969
R10253 VDD.n11472 VDD.n11471 0.969
R10254 VDD.n11470 VDD.n11469 0.969
R10255 VDD.n11448 VDD.n11443 0.969
R10256 VDD.n11392 VDD.n11387 0.969
R10257 VDD.n11250 VDD.n11245 0.969
R10258 VDD.n11193 VDD.n11189 0.969
R10259 VDD.n12260 VDD.n12255 0.969
R10260 VDD.n12266 VDD.n12262 0.969
R10261 VDD.n2975 VDD.n2966 0.955
R10262 VDD.n3041 VDD.n3034 0.955
R10263 VDD.n3074 VDD.n3073 0.955
R10264 VDD.n3149 VDD.n3148 0.955
R10265 VDD.n3213 VDD.n3204 0.955
R10266 VDD.n3278 VDD.n3271 0.955
R10267 VDD.n3311 VDD.n3310 0.955
R10268 VDD.n3387 VDD.n3386 0.955
R10269 VDD.n3450 VDD.n3441 0.955
R10270 VDD.n3516 VDD.n3509 0.955
R10271 VDD.n3549 VDD.n3548 0.955
R10272 VDD.n3624 VDD.n3623 0.955
R10273 VDD.n3688 VDD.n3679 0.955
R10274 VDD.n3753 VDD.n3746 0.955
R10275 VDD.n3786 VDD.n3785 0.955
R10276 VDD.n3862 VDD.n3861 0.955
R10277 VDD.n3925 VDD.n3916 0.955
R10278 VDD.n3991 VDD.n3984 0.955
R10279 VDD.n4024 VDD.n4023 0.955
R10280 VDD.n4099 VDD.n4098 0.955
R10281 VDD.n4163 VDD.n4154 0.955
R10282 VDD.n4228 VDD.n4221 0.955
R10283 VDD.n4261 VDD.n4260 0.955
R10284 VDD.n4337 VDD.n4336 0.955
R10285 VDD.n4400 VDD.n4391 0.955
R10286 VDD.n10117 VDD.n10116 0.955
R10287 VDD.n10309 VDD.n10303 0.948
R10288 VDD.n10271 VDD.n10266 0.948
R10289 VDD.n10190 VDD.n10185 0.948
R10290 VDD.n10154 VDD.n10149 0.948
R10291 VDD.n10065 VDD.n10059 0.948
R10292 VDD.n10072 VDD.n10067 0.948
R10293 VDD.n10020 VDD.n10014 0.948
R10294 VDD.n10027 VDD.n10022 0.948
R10295 VDD.n10656 VDD.n10650 0.948
R10296 VDD.n10618 VDD.n10613 0.948
R10297 VDD.n10536 VDD.n10531 0.948
R10298 VDD.n10500 VDD.n10495 0.948
R10299 VDD.n10227 VDD.n10226 0.939
R10300 VDD.n10574 VDD.n10573 0.939
R10301 VDD.n10463 VDD.n10462 0.939
R10302 VDD.n475 VDD.n466 0.933
R10303 VDD.n475 VDD.n468 0.933
R10304 VDD.n612 VDD.n603 0.933
R10305 VDD.n612 VDD.n605 0.933
R10306 VDD.n708 VDD.n699 0.933
R10307 VDD.n708 VDD.n701 0.933
R10308 VDD.n845 VDD.n836 0.933
R10309 VDD.n845 VDD.n838 0.933
R10310 VDD.n942 VDD.n933 0.933
R10311 VDD.n942 VDD.n935 0.933
R10312 VDD.n1079 VDD.n1070 0.933
R10313 VDD.n1079 VDD.n1072 0.933
R10314 VDD.n1175 VDD.n1166 0.933
R10315 VDD.n1175 VDD.n1168 0.933
R10316 VDD.n1312 VDD.n1303 0.933
R10317 VDD.n1312 VDD.n1305 0.933
R10318 VDD.n1409 VDD.n1400 0.933
R10319 VDD.n1409 VDD.n1402 0.933
R10320 VDD.n1546 VDD.n1537 0.933
R10321 VDD.n1546 VDD.n1539 0.933
R10322 VDD.n1642 VDD.n1633 0.933
R10323 VDD.n1642 VDD.n1635 0.933
R10324 VDD.n1779 VDD.n1770 0.933
R10325 VDD.n1779 VDD.n1772 0.933
R10326 VDD.n11947 VDD.n11946 0.925
R10327 VDD.n12319 VDD.n12318 0.924
R10328 VDD.n5384 VDD.n5383 0.869
R10329 VDD.n5745 VDD.n5744 0.869
R10330 VDD.n6107 VDD.n6106 0.869
R10331 VDD.n6469 VDD.n6468 0.869
R10332 VDD.n6831 VDD.n6830 0.869
R10333 VDD.n7193 VDD.n7192 0.869
R10334 VDD.n7555 VDD.n7554 0.869
R10335 VDD.n7917 VDD.n7916 0.869
R10336 VDD.n8279 VDD.n8278 0.869
R10337 VDD.n8641 VDD.n8640 0.869
R10338 VDD.n9003 VDD.n9002 0.869
R10339 VDD.n9365 VDD.n9364 0.869
R10340 VDD.n9727 VDD.n9726 0.869
R10341 VDD.n12053 VDD.n12052 0.868
R10342 VDD.n11066 VDD.n11065 0.868
R10343 VDD.n10776 VDD.n10775 0.868
R10344 VDD.n10851 VDD.n10850 0.868
R10345 VDD.n10916 VDD.n10915 0.868
R10346 VDD.n11832 VDD.n11831 0.868
R10347 VDD.n11546 VDD.n11545 0.868
R10348 VDD.n12123 VDD.n12122 0.868
R10349 VDD.n11285 VDD.n11284 0.868
R10350 VDD.n5147 VDD.n2699 0.851
R10351 VDD.n5151 VDD.n2608 0.851
R10352 VDD.n2600 VDD.n109 0.851
R10353 VDD.n2599 VDD.n117 0.851
R10354 VDD.n2596 VDD.n180 0.851
R10355 VDD.n2601 VDD.n102 0.85
R10356 VDD.n2597 VDD.n173 0.85
R10357 VDD.n2598 VDD.n164 0.85
R10358 VDD.n5306 VDD.n5305 0.85
R10359 VDD.n494 VDD.n493 0.8
R10360 VDD.n496 VDD.n495 0.8
R10361 VDD.n575 VDD.n574 0.8
R10362 VDD.n577 VDD.n576 0.8
R10363 VDD.n727 VDD.n726 0.8
R10364 VDD.n729 VDD.n728 0.8
R10365 VDD.n808 VDD.n807 0.8
R10366 VDD.n810 VDD.n809 0.8
R10367 VDD.n961 VDD.n960 0.8
R10368 VDD.n963 VDD.n962 0.8
R10369 VDD.n1042 VDD.n1041 0.8
R10370 VDD.n1044 VDD.n1043 0.8
R10371 VDD.n1194 VDD.n1193 0.8
R10372 VDD.n1196 VDD.n1195 0.8
R10373 VDD.n1275 VDD.n1274 0.8
R10374 VDD.n1277 VDD.n1276 0.8
R10375 VDD.n1428 VDD.n1427 0.8
R10376 VDD.n1430 VDD.n1429 0.8
R10377 VDD.n1509 VDD.n1508 0.8
R10378 VDD.n1511 VDD.n1510 0.8
R10379 VDD.n1661 VDD.n1660 0.8
R10380 VDD.n1663 VDD.n1662 0.8
R10381 VDD.n1742 VDD.n1741 0.8
R10382 VDD.n1744 VDD.n1743 0.8
R10383 VDD.n10213 VDD.n10212 0.78
R10384 VDD.n12106 VDD.n12105 0.775
R10385 VDD.n12061 VDD.n12060 0.775
R10386 VDD.n10921 VDD.n10919 0.775
R10387 VDD.n11044 VDD.n11043 0.775
R10388 VDD.n11086 VDD.n11085 0.775
R10389 VDD.n11009 VDD.n11008 0.775
R10390 VDD.n10995 VDD.n10994 0.775
R10391 VDD.n11099 VDD.n11098 0.775
R10392 VDD.n10871 VDD.n10870 0.775
R10393 VDD.n11720 VDD.n11718 0.775
R10394 VDD.n11811 VDD.n11810 0.775
R10395 VDD.n11853 VDD.n11852 0.775
R10396 VDD.n11777 VDD.n11776 0.775
R10397 VDD.n11764 VDD.n11763 0.775
R10398 VDD.n11874 VDD.n11873 0.775
R10399 VDD.n11588 VDD.n11587 0.775
R10400 VDD.n11339 VDD.n11338 0.775
R10401 VDD.n11293 VDD.n11292 0.775
R10402 VDD.n10245 VDD.n10244 0.767
R10403 VDD.n10592 VDD.n10591 0.767
R10404 VDD.n10559 VDD.n10558 0.767
R10405 VDD.n2975 VDD.n2968 0.764
R10406 VDD.n3027 VDD.n3018 0.764
R10407 VDD.n3090 VDD.n3089 0.764
R10408 VDD.n3147 VDD.n3146 0.764
R10409 VDD.n3213 VDD.n3206 0.764
R10410 VDD.n3264 VDD.n3255 0.764
R10411 VDD.n3328 VDD.n3327 0.764
R10412 VDD.n3385 VDD.n3384 0.764
R10413 VDD.n3450 VDD.n3443 0.764
R10414 VDD.n3502 VDD.n3493 0.764
R10415 VDD.n3565 VDD.n3564 0.764
R10416 VDD.n3622 VDD.n3621 0.764
R10417 VDD.n3688 VDD.n3681 0.764
R10418 VDD.n3739 VDD.n3730 0.764
R10419 VDD.n3803 VDD.n3802 0.764
R10420 VDD.n3860 VDD.n3859 0.764
R10421 VDD.n3925 VDD.n3918 0.764
R10422 VDD.n3977 VDD.n3968 0.764
R10423 VDD.n4040 VDD.n4039 0.764
R10424 VDD.n4097 VDD.n4096 0.764
R10425 VDD.n4163 VDD.n4156 0.764
R10426 VDD.n4214 VDD.n4205 0.764
R10427 VDD.n4278 VDD.n4277 0.764
R10428 VDD.n4335 VDD.n4334 0.764
R10429 VDD.n4400 VDD.n4393 0.764
R10430 VDD.n4452 VDD.n4443 0.764
R10431 VDD.n5319 VDD.n5318 0.752
R10432 VDD.n5516 VDD.n5515 0.752
R10433 VDD.n5606 VDD.n5605 0.752
R10434 VDD.n5628 VDD.n5626 0.752
R10435 VDD.n5647 VDD.n5646 0.752
R10436 VDD.n5658 VDD.n5657 0.752
R10437 VDD.n5680 VDD.n5679 0.752
R10438 VDD.n5877 VDD.n5876 0.752
R10439 VDD.n5967 VDD.n5966 0.752
R10440 VDD.n5989 VDD.n5987 0.752
R10441 VDD.n6008 VDD.n6007 0.752
R10442 VDD.n6019 VDD.n6018 0.752
R10443 VDD.n6042 VDD.n6041 0.752
R10444 VDD.n6239 VDD.n6238 0.752
R10445 VDD.n6329 VDD.n6328 0.752
R10446 VDD.n6351 VDD.n6349 0.752
R10447 VDD.n6370 VDD.n6369 0.752
R10448 VDD.n6381 VDD.n6380 0.752
R10449 VDD.n6404 VDD.n6403 0.752
R10450 VDD.n6601 VDD.n6600 0.752
R10451 VDD.n6691 VDD.n6690 0.752
R10452 VDD.n6713 VDD.n6711 0.752
R10453 VDD.n6732 VDD.n6731 0.752
R10454 VDD.n6743 VDD.n6742 0.752
R10455 VDD.n6766 VDD.n6765 0.752
R10456 VDD.n6963 VDD.n6962 0.752
R10457 VDD.n7053 VDD.n7052 0.752
R10458 VDD.n7075 VDD.n7073 0.752
R10459 VDD.n7094 VDD.n7093 0.752
R10460 VDD.n7105 VDD.n7104 0.752
R10461 VDD.n7128 VDD.n7127 0.752
R10462 VDD.n7325 VDD.n7324 0.752
R10463 VDD.n7415 VDD.n7414 0.752
R10464 VDD.n7437 VDD.n7435 0.752
R10465 VDD.n7456 VDD.n7455 0.752
R10466 VDD.n7467 VDD.n7466 0.752
R10467 VDD.n7490 VDD.n7489 0.752
R10468 VDD.n7687 VDD.n7686 0.752
R10469 VDD.n7777 VDD.n7776 0.752
R10470 VDD.n7799 VDD.n7797 0.752
R10471 VDD.n7818 VDD.n7817 0.752
R10472 VDD.n7829 VDD.n7828 0.752
R10473 VDD.n7852 VDD.n7851 0.752
R10474 VDD.n8049 VDD.n8048 0.752
R10475 VDD.n8139 VDD.n8138 0.752
R10476 VDD.n8161 VDD.n8159 0.752
R10477 VDD.n8180 VDD.n8179 0.752
R10478 VDD.n8191 VDD.n8190 0.752
R10479 VDD.n8214 VDD.n8213 0.752
R10480 VDD.n8411 VDD.n8410 0.752
R10481 VDD.n8501 VDD.n8500 0.752
R10482 VDD.n8523 VDD.n8521 0.752
R10483 VDD.n8542 VDD.n8541 0.752
R10484 VDD.n8553 VDD.n8552 0.752
R10485 VDD.n8576 VDD.n8575 0.752
R10486 VDD.n8773 VDD.n8772 0.752
R10487 VDD.n8863 VDD.n8862 0.752
R10488 VDD.n8885 VDD.n8883 0.752
R10489 VDD.n8904 VDD.n8903 0.752
R10490 VDD.n8915 VDD.n8914 0.752
R10491 VDD.n8938 VDD.n8937 0.752
R10492 VDD.n9135 VDD.n9134 0.752
R10493 VDD.n9225 VDD.n9224 0.752
R10494 VDD.n9247 VDD.n9245 0.752
R10495 VDD.n9266 VDD.n9265 0.752
R10496 VDD.n9277 VDD.n9276 0.752
R10497 VDD.n9300 VDD.n9299 0.752
R10498 VDD.n9497 VDD.n9496 0.752
R10499 VDD.n9587 VDD.n9586 0.752
R10500 VDD.n9609 VDD.n9607 0.752
R10501 VDD.n9628 VDD.n9627 0.752
R10502 VDD.n9639 VDD.n9638 0.752
R10503 VDD.n9662 VDD.n9661 0.752
R10504 VDD.n9859 VDD.n9858 0.752
R10505 VDD.n9949 VDD.n9948 0.752
R10506 VDD.n9971 VDD.n9969 0.752
R10507 VDD.n9990 VDD.n9989 0.752
R10508 VDD.n10001 VDD.n10000 0.752
R10509 VDD.n11460 VDD.n11185 0.75
R10510 VDD.n16 VDD.n15 0.747
R10511 VDD.n2135 VDD.n2134 0.738
R10512 VDD.n2184 VDD.n2183 0.738
R10513 VDD.n2366 VDD.n2365 0.738
R10514 VDD.n2415 VDD.n2414 0.738
R10515 VDD.n2553 VDD.n2552 0.738
R10516 VDD.n120 VDD.n119 0.738
R10517 VDD.n5194 VDD.n5193 0.738
R10518 VDD.n5261 VDD.n5260 0.738
R10519 VDD.n5019 VDD.n5018 0.738
R10520 VDD.n4970 VDD.n4969 0.738
R10521 VDD.n4788 VDD.n4787 0.738
R10522 VDD.n4739 VDD.n4738 0.738
R10523 VDD.n5383 VDD.n5382 0.729
R10524 VDD.n5744 VDD.n5743 0.729
R10525 VDD.n6106 VDD.n6105 0.729
R10526 VDD.n6468 VDD.n6467 0.729
R10527 VDD.n6830 VDD.n6829 0.729
R10528 VDD.n7192 VDD.n7191 0.729
R10529 VDD.n7554 VDD.n7553 0.729
R10530 VDD.n7916 VDD.n7915 0.729
R10531 VDD.n8278 VDD.n8277 0.729
R10532 VDD.n8640 VDD.n8639 0.729
R10533 VDD.n9002 VDD.n9001 0.729
R10534 VDD.n9364 VDD.n9363 0.729
R10535 VDD.n9726 VDD.n9725 0.729
R10536 VDD.n5667 VDD.n5666 0.725
R10537 VDD.n6028 VDD.n6027 0.725
R10538 VDD.n6390 VDD.n6389 0.725
R10539 VDD.n6752 VDD.n6751 0.725
R10540 VDD.n7114 VDD.n7113 0.725
R10541 VDD.n7476 VDD.n7475 0.725
R10542 VDD.n7838 VDD.n7837 0.725
R10543 VDD.n8200 VDD.n8199 0.725
R10544 VDD.n8562 VDD.n8561 0.725
R10545 VDD.n8924 VDD.n8923 0.725
R10546 VDD.n9286 VDD.n9285 0.725
R10547 VDD.n9648 VDD.n9647 0.725
R10548 VDD.n10010 VDD.n10009 0.725
R10549 VDD.n11849 VDD.n11848 0.723
R10550 VDD.n11468 VDD.n11467 0.723
R10551 VDD.n11273 VDD.n11272 0.723
R10552 VDD.n10 VDD.n9 0.705
R10553 VDD.n12241 VDD.n12240 0.705
R10554 VDD.n10448 VDD.n10447 0.701
R10555 VDD.n12247 VDD.n12246 0.682
R10556 VDD.n335 VDD.n334 0.68
R10557 VDD.n12227 VDD.n11942 0.679
R10558 VDD.n5145 VDD.n5129 0.675
R10559 VDD.n5149 VDD.n2692 0.675
R10560 VDD.n195 VDD.n193 0.675
R10561 VDD.n5144 VDD.n5143 0.675
R10562 VDD.n2594 VDD.n2593 0.675
R10563 VDD.n392 VDD.n383 0.666
R10564 VDD.n392 VDD.n385 0.666
R10565 VDD.n461 VDD.n452 0.666
R10566 VDD.n461 VDD.n454 0.666
R10567 VDD.n626 VDD.n617 0.666
R10568 VDD.n626 VDD.n619 0.666
R10569 VDD.n694 VDD.n685 0.666
R10570 VDD.n694 VDD.n687 0.666
R10571 VDD.n859 VDD.n850 0.666
R10572 VDD.n859 VDD.n852 0.666
R10573 VDD.n928 VDD.n919 0.666
R10574 VDD.n928 VDD.n921 0.666
R10575 VDD.n1093 VDD.n1084 0.666
R10576 VDD.n1093 VDD.n1086 0.666
R10577 VDD.n1161 VDD.n1152 0.666
R10578 VDD.n1161 VDD.n1154 0.666
R10579 VDD.n1326 VDD.n1317 0.666
R10580 VDD.n1326 VDD.n1319 0.666
R10581 VDD.n1395 VDD.n1386 0.666
R10582 VDD.n1395 VDD.n1388 0.666
R10583 VDD.n1560 VDD.n1551 0.666
R10584 VDD.n1560 VDD.n1553 0.666
R10585 VDD.n1628 VDD.n1619 0.666
R10586 VDD.n1628 VDD.n1621 0.666
R10587 VDD.n1793 VDD.n1784 0.666
R10588 VDD.n1793 VDD.n1786 0.666
R10589 VDD.n1959 VDD.n1958 0.656
R10590 VDD.n11961 VDD.n11959 0.622
R10591 VDD.n11196 VDD.n11194 0.622
R10592 VDD.n11727 VDD.n11726 0.609
R10593 VDD.n10958 VDD.n10957 0.609
R10594 VDD.n11553 VDD.n11552 0.608
R10595 VDD.n10783 VDD.n10782 0.608
R10596 VDD.n2886 VDD.n2885 0.604
R10597 VDD.n4520 VDD.n4519 0.604
R10598 VDD.n10201 VDD.n10200 0.598
R10599 VDD.n10320 VDD.n10319 0.587
R10600 VDD.n10667 VDD.n10666 0.587
R10601 VDD.n10547 VDD.n10546 0.587
R10602 VDD.n81 VDD.n75 0.581
R10603 VDD.n47 VDD.n41 0.581
R10604 VDD.n12208 VDD.n12203 0.581
R10605 VDD.n12174 VDD.n12169 0.581
R10606 VDD.n12004 VDD.n11999 0.581
R10607 VDD.n11970 VDD.n11965 0.581
R10608 VDD.n11052 VDD.n11042 0.581
R10609 VDD.n11051 VDD.n11045 0.581
R10610 VDD.n10984 VDD.n10983 0.581
R10611 VDD.n11009 VDD.n11006 0.581
R10612 VDD.n11164 VDD.n11159 0.581
R10613 VDD.n11113 VDD.n11108 0.581
R10614 VDD.n10767 VDD.n10766 0.581
R10615 VDD.n10780 VDD.n10777 0.581
R10616 VDD.n11818 VDD.n11809 0.581
R10617 VDD.n11817 VDD.n11812 0.581
R10618 VDD.n11753 VDD.n11752 0.581
R10619 VDD.n11777 VDD.n11774 0.581
R10620 VDD.n11922 VDD.n11917 0.581
R10621 VDD.n11893 VDD.n11888 0.581
R10622 VDD.n11537 VDD.n11536 0.581
R10623 VDD.n11550 VDD.n11547 0.581
R10624 VDD.n11436 VDD.n11431 0.581
R10625 VDD.n11404 VDD.n11399 0.581
R10626 VDD.n11238 VDD.n11233 0.581
R10627 VDD.n11206 VDD.n11200 0.581
R10628 VDD.n12312 VDD.n12306 0.581
R10629 VDD.n12278 VDD.n12272 0.581
R10630 VDD.n2989 VDD.n2980 0.573
R10631 VDD.n3027 VDD.n3020 0.573
R10632 VDD.n3088 VDD.n3087 0.573
R10633 VDD.n3135 VDD.n3134 0.573
R10634 VDD.n3227 VDD.n3218 0.573
R10635 VDD.n3264 VDD.n3257 0.573
R10636 VDD.n3326 VDD.n3325 0.573
R10637 VDD.n3373 VDD.n3372 0.573
R10638 VDD.n3464 VDD.n3455 0.573
R10639 VDD.n3502 VDD.n3495 0.573
R10640 VDD.n3563 VDD.n3562 0.573
R10641 VDD.n3610 VDD.n3609 0.573
R10642 VDD.n3702 VDD.n3693 0.573
R10643 VDD.n3739 VDD.n3732 0.573
R10644 VDD.n3801 VDD.n3800 0.573
R10645 VDD.n3848 VDD.n3847 0.573
R10646 VDD.n3939 VDD.n3930 0.573
R10647 VDD.n3977 VDD.n3970 0.573
R10648 VDD.n4038 VDD.n4037 0.573
R10649 VDD.n4085 VDD.n4084 0.573
R10650 VDD.n4177 VDD.n4168 0.573
R10651 VDD.n4214 VDD.n4207 0.573
R10652 VDD.n4276 VDD.n4275 0.573
R10653 VDD.n4323 VDD.n4322 0.573
R10654 VDD.n4414 VDD.n4405 0.573
R10655 VDD.n4452 VDD.n4445 0.573
R10656 VDD.n12028 VDD.n12027 0.572
R10657 VDD.n11005 VDD.n11004 0.572
R10658 VDD.n10714 VDD.n10713 0.572
R10659 VDD.n11094 VDD.n11093 0.572
R10660 VDD.n10888 VDD.n10887 0.572
R10661 VDD.n11773 VDD.n11772 0.572
R10662 VDD.n11484 VDD.n11483 0.572
R10663 VDD.n12148 VDD.n12147 0.572
R10664 VDD.n11261 VDD.n11260 0.572
R10665 VDD.n4550 VDD.n4549 0.545
R10666 VDD.n508 VDD.n507 0.533
R10667 VDD.n510 VDD.n509 0.533
R10668 VDD.n560 VDD.n559 0.533
R10669 VDD.n562 VDD.n561 0.533
R10670 VDD.n742 VDD.n741 0.533
R10671 VDD.n744 VDD.n743 0.533
R10672 VDD.n794 VDD.n793 0.533
R10673 VDD.n796 VDD.n795 0.533
R10674 VDD.n975 VDD.n974 0.533
R10675 VDD.n977 VDD.n976 0.533
R10676 VDD.n1027 VDD.n1026 0.533
R10677 VDD.n1029 VDD.n1028 0.533
R10678 VDD.n1209 VDD.n1208 0.533
R10679 VDD.n1211 VDD.n1210 0.533
R10680 VDD.n1261 VDD.n1260 0.533
R10681 VDD.n1263 VDD.n1262 0.533
R10682 VDD.n1442 VDD.n1441 0.533
R10683 VDD.n1444 VDD.n1443 0.533
R10684 VDD.n1494 VDD.n1493 0.533
R10685 VDD.n1496 VDD.n1495 0.533
R10686 VDD.n1676 VDD.n1675 0.533
R10687 VDD.n1678 VDD.n1677 0.533
R10688 VDD.n1728 VDD.n1727 0.533
R10689 VDD.n1730 VDD.n1729 0.533
R10690 VDD.n2825 VDD.n2812 0.513
R10691 VDD.n255 VDD.n229 0.51
R10692 VDD.n2044 VDD.n2037 0.492
R10693 VDD.n2058 VDD.n2051 0.492
R10694 VDD.n2275 VDD.n2268 0.492
R10695 VDD.n2289 VDD.n2282 0.492
R10696 VDD.n2514 VDD.n2507 0.492
R10697 VDD.n2585 VDD.n2584 0.492
R10698 VDD.n5117 VDD.n5110 0.492
R10699 VDD.n4893 VDD.n4886 0.492
R10700 VDD.n4879 VDD.n4872 0.492
R10701 VDD.n4662 VDD.n4655 0.492
R10702 VDD.n4648 VDD.n4641 0.492
R10703 VDD.n10296 VDD.n10291 0.474
R10704 VDD.n10284 VDD.n10278 0.474
R10705 VDD.n10178 VDD.n10173 0.474
R10706 VDD.n10166 VDD.n10161 0.474
R10707 VDD.n10096 VDD.n10090 0.474
R10708 VDD.n10083 VDD.n10078 0.474
R10709 VDD.n10051 VDD.n10046 0.474
R10710 VDD.n10039 VDD.n10033 0.474
R10711 VDD.n10643 VDD.n10638 0.474
R10712 VDD.n10631 VDD.n10625 0.474
R10713 VDD.n10524 VDD.n10519 0.474
R10714 VDD.n10512 VDD.n10507 0.474
R10715 VDD.n4463 VDD.n4462 0.436
R10716 VDD.n10567 VDD.n10449 0.425
R10717 VDD.n11476 VDD.n11475 0.416
R10718 VDD.n11760 VDD.n11759 0.416
R10719 VDD.n11649 VDD.n11648 0.416
R10720 VDD.n11447 VDD.n11446 0.416
R10721 VDD.n11249 VDD.n11248 0.416
R10722 VDD.n10189 VDD.n10188 0.407
R10723 VDD.n10064 VDD.n10063 0.407
R10724 VDD.n10026 VDD.n10025 0.407
R10725 VDD.n10270 VDD.n10269 0.4
R10726 VDD.n10617 VDD.n10616 0.4
R10727 VDD.n10535 VDD.n10534 0.4
R10728 VDD.n4552 VDD.n4551 0.4
R10729 VDD.n406 VDD.n397 0.4
R10730 VDD.n406 VDD.n399 0.4
R10731 VDD.n447 VDD.n438 0.4
R10732 VDD.n447 VDD.n440 0.4
R10733 VDD.n640 VDD.n631 0.4
R10734 VDD.n640 VDD.n633 0.4
R10735 VDD.n680 VDD.n671 0.4
R10736 VDD.n680 VDD.n673 0.4
R10737 VDD.n873 VDD.n864 0.4
R10738 VDD.n873 VDD.n866 0.4
R10739 VDD.n914 VDD.n905 0.4
R10740 VDD.n914 VDD.n907 0.4
R10741 VDD.n1107 VDD.n1098 0.4
R10742 VDD.n1107 VDD.n1100 0.4
R10743 VDD.n1147 VDD.n1138 0.4
R10744 VDD.n1147 VDD.n1140 0.4
R10745 VDD.n1340 VDD.n1331 0.4
R10746 VDD.n1340 VDD.n1333 0.4
R10747 VDD.n1381 VDD.n1372 0.4
R10748 VDD.n1381 VDD.n1374 0.4
R10749 VDD.n1574 VDD.n1565 0.4
R10750 VDD.n1574 VDD.n1567 0.4
R10751 VDD.n1614 VDD.n1605 0.4
R10752 VDD.n1614 VDD.n1607 0.4
R10753 VDD.n1807 VDD.n1798 0.4
R10754 VDD.n1807 VDD.n1800 0.4
R10755 VDD.n1848 VDD.n1839 0.4
R10756 VDD.n1848 VDD.n1841 0.4
R10757 VDD.n1859 VDD.n1858 0.393
R10758 VDD.n12094 VDD.n12093 0.387
R10759 VDD.n12074 VDD.n12073 0.387
R10760 VDD.n10918 VDD.n10917 0.387
R10761 VDD.n10929 VDD.n10928 0.387
R10762 VDD.n10931 VDD.n10930 0.387
R10763 VDD.n10937 VDD.n10936 0.387
R10764 VDD.n11035 VDD.n11027 0.387
R10765 VDD.n11029 VDD.n11028 0.387
R10766 VDD.n11116 VDD.n11113 0.387
R10767 VDD.n11115 VDD.n11114 0.387
R10768 VDD.n11096 VDD.n11095 0.387
R10769 VDD.n10857 VDD.n10856 0.387
R10770 VDD.n10837 VDD.n10831 0.387
R10771 VDD.n10839 VDD.n10838 0.387
R10772 VDD.n10812 VDD.n10811 0.387
R10773 VDD.n10819 VDD.n10818 0.387
R10774 VDD.n10736 VDD.n10735 0.387
R10775 VDD.n11686 VDD.n11685 0.387
R10776 VDD.n11709 VDD.n11708 0.387
R10777 VDD.n11711 VDD.n11710 0.387
R10778 VDD.n11692 VDD.n11691 0.387
R10779 VDD.n11802 VDD.n11794 0.387
R10780 VDD.n11796 VDD.n11795 0.387
R10781 VDD.n11896 VDD.n11893 0.387
R10782 VDD.n11895 VDD.n11894 0.387
R10783 VDD.n11871 VDD.n11870 0.387
R10784 VDD.n11638 VDD.n11637 0.387
R10785 VDD.n11616 VDD.n11611 0.387
R10786 VDD.n11618 VDD.n11617 0.387
R10787 VDD.n11594 VDD.n11593 0.387
R10788 VDD.n11603 VDD.n11602 0.387
R10789 VDD.n11507 VDD.n11506 0.387
R10790 VDD.n11325 VDD.n11324 0.387
R10791 VDD.n11305 VDD.n11304 0.387
R10792 VDD.n2778 VDD.n2777 0.382
R10793 VDD.n2989 VDD.n2982 0.382
R10794 VDD.n3013 VDD.n3004 0.382
R10795 VDD.n3104 VDD.n3103 0.382
R10796 VDD.n3133 VDD.n3132 0.382
R10797 VDD.n3227 VDD.n3220 0.382
R10798 VDD.n3250 VDD.n3241 0.382
R10799 VDD.n3342 VDD.n3341 0.382
R10800 VDD.n3371 VDD.n3370 0.382
R10801 VDD.n3464 VDD.n3457 0.382
R10802 VDD.n3488 VDD.n3479 0.382
R10803 VDD.n3579 VDD.n3578 0.382
R10804 VDD.n3608 VDD.n3607 0.382
R10805 VDD.n3702 VDD.n3695 0.382
R10806 VDD.n3725 VDD.n3716 0.382
R10807 VDD.n3817 VDD.n3816 0.382
R10808 VDD.n3846 VDD.n3845 0.382
R10809 VDD.n3939 VDD.n3932 0.382
R10810 VDD.n3963 VDD.n3954 0.382
R10811 VDD.n4054 VDD.n4053 0.382
R10812 VDD.n4083 VDD.n4082 0.382
R10813 VDD.n4177 VDD.n4170 0.382
R10814 VDD.n4200 VDD.n4191 0.382
R10815 VDD.n4292 VDD.n4291 0.382
R10816 VDD.n4321 VDD.n4320 0.382
R10817 VDD.n4414 VDD.n4407 0.382
R10818 VDD.n4438 VDD.n4429 0.382
R10819 VDD.n5325 VDD.n5324 0.376
R10820 VDD.n5328 VDD.n5327 0.376
R10821 VDD.n5475 VDD.n5474 0.376
R10822 VDD.n5487 VDD.n5486 0.376
R10823 VDD.n5497 VDD.n5496 0.376
R10824 VDD.n5507 VDD.n5506 0.376
R10825 VDD.n5686 VDD.n5685 0.376
R10826 VDD.n5689 VDD.n5688 0.376
R10827 VDD.n5836 VDD.n5835 0.376
R10828 VDD.n5848 VDD.n5847 0.376
R10829 VDD.n5858 VDD.n5857 0.376
R10830 VDD.n5868 VDD.n5867 0.376
R10831 VDD.n6048 VDD.n6047 0.376
R10832 VDD.n6051 VDD.n6050 0.376
R10833 VDD.n6198 VDD.n6197 0.376
R10834 VDD.n6210 VDD.n6209 0.376
R10835 VDD.n6220 VDD.n6219 0.376
R10836 VDD.n6230 VDD.n6229 0.376
R10837 VDD.n6410 VDD.n6409 0.376
R10838 VDD.n6413 VDD.n6412 0.376
R10839 VDD.n6560 VDD.n6559 0.376
R10840 VDD.n6572 VDD.n6571 0.376
R10841 VDD.n6582 VDD.n6581 0.376
R10842 VDD.n6592 VDD.n6591 0.376
R10843 VDD.n6772 VDD.n6771 0.376
R10844 VDD.n6775 VDD.n6774 0.376
R10845 VDD.n6922 VDD.n6921 0.376
R10846 VDD.n6934 VDD.n6933 0.376
R10847 VDD.n6944 VDD.n6943 0.376
R10848 VDD.n6954 VDD.n6953 0.376
R10849 VDD.n7134 VDD.n7133 0.376
R10850 VDD.n7137 VDD.n7136 0.376
R10851 VDD.n7284 VDD.n7283 0.376
R10852 VDD.n7296 VDD.n7295 0.376
R10853 VDD.n7306 VDD.n7305 0.376
R10854 VDD.n7316 VDD.n7315 0.376
R10855 VDD.n7496 VDD.n7495 0.376
R10856 VDD.n7499 VDD.n7498 0.376
R10857 VDD.n7646 VDD.n7645 0.376
R10858 VDD.n7658 VDD.n7657 0.376
R10859 VDD.n7668 VDD.n7667 0.376
R10860 VDD.n7678 VDD.n7677 0.376
R10861 VDD.n7858 VDD.n7857 0.376
R10862 VDD.n7861 VDD.n7860 0.376
R10863 VDD.n8008 VDD.n8007 0.376
R10864 VDD.n8020 VDD.n8019 0.376
R10865 VDD.n8030 VDD.n8029 0.376
R10866 VDD.n8040 VDD.n8039 0.376
R10867 VDD.n8220 VDD.n8219 0.376
R10868 VDD.n8223 VDD.n8222 0.376
R10869 VDD.n8370 VDD.n8369 0.376
R10870 VDD.n8382 VDD.n8381 0.376
R10871 VDD.n8392 VDD.n8391 0.376
R10872 VDD.n8402 VDD.n8401 0.376
R10873 VDD.n8582 VDD.n8581 0.376
R10874 VDD.n8585 VDD.n8584 0.376
R10875 VDD.n8732 VDD.n8731 0.376
R10876 VDD.n8744 VDD.n8743 0.376
R10877 VDD.n8754 VDD.n8753 0.376
R10878 VDD.n8764 VDD.n8763 0.376
R10879 VDD.n8944 VDD.n8943 0.376
R10880 VDD.n8947 VDD.n8946 0.376
R10881 VDD.n9094 VDD.n9093 0.376
R10882 VDD.n9106 VDD.n9105 0.376
R10883 VDD.n9116 VDD.n9115 0.376
R10884 VDD.n9126 VDD.n9125 0.376
R10885 VDD.n9306 VDD.n9305 0.376
R10886 VDD.n9309 VDD.n9308 0.376
R10887 VDD.n9456 VDD.n9455 0.376
R10888 VDD.n9468 VDD.n9467 0.376
R10889 VDD.n9478 VDD.n9477 0.376
R10890 VDD.n9488 VDD.n9487 0.376
R10891 VDD.n9668 VDD.n9667 0.376
R10892 VDD.n9671 VDD.n9670 0.376
R10893 VDD.n9818 VDD.n9817 0.376
R10894 VDD.n9830 VDD.n9829 0.376
R10895 VDD.n9840 VDD.n9839 0.376
R10896 VDD.n9850 VDD.n9849 0.376
R10897 VDD.n223 VDD.n222 0.374
R10898 VDD.n265 VDD.n260 0.374
R10899 VDD.n2832 VDD.n2828 0.366
R10900 VDD.n2850 VDD.n2844 0.366
R10901 VDD.n2928 VDD.n2927 0.366
R10902 VDD.n4483 VDD.n4482 0.363
R10903 VDD.n4540 VDD.n4537 0.363
R10904 VDD.n4622 VDD.n4569 0.363
R10905 VDD.n4634 VDD.n4633 0.341
R10906 VDD.n235 VDD.n231 0.34
R10907 VDD.n347 VDD.n346 0.34
R10908 VDD.n2799 VDD.n2797 0.33
R10909 VDD.n1876 VDD.n1875 0.328
R10910 VDD.n1934 VDD.n1928 0.328
R10911 VDD.n1937 VDD.n1936 0.328
R10912 VDD.n4566 VDD.n4564 0.327
R10913 VDD.n327 VDD.n314 0.306
R10914 VDD.n327 VDD.n320 0.306
R10915 VDD.n1963 VDD.n1961 0.295
R10916 VDD.n2900 VDD.n2899 0.293
R10917 VDD.n2901 VDD.n2900 0.293
R10918 VDD.n2914 VDD.n2907 0.293
R10919 VDD.n4491 VDD.n4481 0.29
R10920 VDD.n4503 VDD.n4502 0.29
R10921 VDD.n10449 VDD.n10448 0.275
R10922 VDD.n224 VDD.n223 0.272
R10923 VDD.n314 VDD.n313 0.272
R10924 VDD.n350 VDD.n349 0.272
R10925 VDD.n522 VDD.n521 0.266
R10926 VDD.n524 VDD.n523 0.266
R10927 VDD.n546 VDD.n545 0.266
R10928 VDD.n548 VDD.n547 0.266
R10929 VDD.n756 VDD.n755 0.266
R10930 VDD.n758 VDD.n757 0.266
R10931 VDD.n780 VDD.n779 0.266
R10932 VDD.n782 VDD.n781 0.266
R10933 VDD.n989 VDD.n988 0.266
R10934 VDD.n991 VDD.n990 0.266
R10935 VDD.n1013 VDD.n1012 0.266
R10936 VDD.n1015 VDD.n1014 0.266
R10937 VDD.n1223 VDD.n1222 0.266
R10938 VDD.n1225 VDD.n1224 0.266
R10939 VDD.n1247 VDD.n1246 0.266
R10940 VDD.n1249 VDD.n1248 0.266
R10941 VDD.n1456 VDD.n1455 0.266
R10942 VDD.n1458 VDD.n1457 0.266
R10943 VDD.n1480 VDD.n1479 0.266
R10944 VDD.n1482 VDD.n1481 0.266
R10945 VDD.n1690 VDD.n1689 0.266
R10946 VDD.n1692 VDD.n1691 0.266
R10947 VDD.n1714 VDD.n1713 0.266
R10948 VDD.n1716 VDD.n1715 0.266
R10949 VDD.n204 VDD.n203 0.266
R10950 VDD.n206 VDD.n205 0.266
R10951 VDD.n1895 VDD.n1894 0.262
R10952 VDD.n2793 VDD.n2792 0.256
R10953 VDD.n2884 VDD.n2883 0.256
R10954 VDD.n2927 VDD.n2926 0.256
R10955 VDD.n2953 VDD.n2951 0.256
R10956 VDD.n2931 VDD.n2930 0.256
R10957 VDD.n12207 VDD.n12206 0.254
R10958 VDD.n12003 VDD.n12002 0.254
R10959 VDD.n11163 VDD.n11162 0.254
R10960 VDD.n11112 VDD.n11111 0.254
R10961 VDD.n11921 VDD.n11920 0.254
R10962 VDD.n12173 VDD.n12172 0.254
R10963 VDD.n11969 VDD.n11968 0.254
R10964 VDD.n11435 VDD.n11434 0.254
R10965 VDD.n11237 VDD.n11236 0.254
R10966 VDD.n4457 VDD.n4456 0.254
R10967 VDD.n4496 VDD.n4495 0.254
R10968 VDD.n4524 VDD.n4523 0.254
R10969 VDD.n4622 VDD.n4566 0.254
R10970 VDD.n2149 VDD.n2148 0.246
R10971 VDD.n2169 VDD.n2168 0.246
R10972 VDD.n2380 VDD.n2379 0.246
R10973 VDD.n2400 VDD.n2399 0.246
R10974 VDD.n5214 VDD.n5213 0.246
R10975 VDD.n5280 VDD.n5279 0.246
R10976 VDD.n5004 VDD.n5003 0.246
R10977 VDD.n4984 VDD.n4983 0.246
R10978 VDD.n4773 VDD.n4772 0.246
R10979 VDD.n4753 VDD.n4752 0.246
R10980 VDD.n278 VDD.n271 0.238
R10981 VDD.n296 VDD.n283 0.238
R10982 VDD.n378 VDD.n371 0.238
R10983 VDD.n370 VDD.n368 0.238
R10984 VDD.n10448 VDD.n10341 0.237
R10985 VDD.n1884 VDD.n1874 0.229
R10986 VDD.n1890 VDD.n1889 0.229
R10987 VDD.n1903 VDD.n1896 0.229
R10988 VDD.n2800 VDD.n2799 0.22
R10989 VDD.n2865 VDD.n2858 0.22
R10990 VDD.n2870 VDD.n2869 0.22
R10991 VDD.n2881 VDD.n2870 0.22
R10992 VDD.n2906 VDD.n2903 0.22
R10993 VDD.n2961 VDD.n2954 0.22
R10994 VDD.n4460 VDD.n4458 0.218
R10995 VDD.n4471 VDD.n4461 0.218
R10996 VDD.n4511 VDD.n4504 0.218
R10997 VDD.n4531 VDD.n4521 0.218
R10998 VDD.n4523 VDD.n4522 0.218
R10999 VDD.n10177 VDD.n10176 0.208
R11000 VDD.n10082 VDD.n10081 0.208
R11001 VDD.n10050 VDD.n10049 0.208
R11002 VDD.n10295 VDD.n10294 0.205
R11003 VDD.n10642 VDD.n10641 0.205
R11004 VDD.n10523 VDD.n10522 0.205
R11005 VDD.n222 VDD.n221 0.204
R11006 VDD.n283 VDD.n282 0.204
R11007 VDD.n299 VDD.n298 0.204
R11008 VDD.n319 VDD.n315 0.204
R11009 VDD.n346 VDD.n345 0.204
R11010 VDD.n1853 VDD.n1852 0.196
R11011 VDD.n1856 VDD.n1854 0.196
R11012 VDD.n1909 VDD.n1908 0.196
R11013 VDD.n1915 VDD.n1914 0.196
R11014 VDD.n1914 VDD.n1913 0.196
R11015 VDD.n2017 VDD.n1963 0.196
R11016 VDD.n68 VDD.n62 0.193
R11017 VDD.n59 VDD.n54 0.193
R11018 VDD.n12196 VDD.n12190 0.193
R11019 VDD.n12187 VDD.n12181 0.193
R11020 VDD.n11992 VDD.n11986 0.193
R11021 VDD.n11983 VDD.n11977 0.193
R11022 VDD.n11068 VDD.n11059 0.193
R11023 VDD.n11067 VDD.n11062 0.193
R11024 VDD.n11016 VDD.n11015 0.193
R11025 VDD.n10986 VDD.n10985 0.193
R11026 VDD.n10995 VDD.n10992 0.193
R11027 VDD.n11157 VDD.n11156 0.193
R11028 VDD.n11165 VDD.n11164 0.193
R11029 VDD.n11179 VDD.n11178 0.193
R11030 VDD.n11178 VDD.n11172 0.193
R11031 VDD.n11149 VDD.n11143 0.193
R11032 VDD.n11151 VDD.n11149 0.193
R11033 VDD.n10743 VDD.n10734 0.193
R11034 VDD.n10742 VDD.n10737 0.193
R11035 VDD.n10758 VDD.n10757 0.193
R11036 VDD.n10756 VDD.n10755 0.193
R11037 VDD.n11834 VDD.n11825 0.193
R11038 VDD.n11833 VDD.n11828 0.193
R11039 VDD.n11840 VDD.n11839 0.193
R11040 VDD.n11756 VDD.n11755 0.193
R11041 VDD.n11764 VDD.n11761 0.193
R11042 VDD.n11915 VDD.n11914 0.193
R11043 VDD.n11923 VDD.n11922 0.193
R11044 VDD.n11936 VDD.n11935 0.193
R11045 VDD.n11935 VDD.n11930 0.193
R11046 VDD.n11907 VDD.n11902 0.193
R11047 VDD.n11909 VDD.n11907 0.193
R11048 VDD.n11514 VDD.n11505 0.193
R11049 VDD.n11513 VDD.n11508 0.193
R11050 VDD.n11528 VDD.n11527 0.193
R11051 VDD.n11526 VDD.n11525 0.193
R11052 VDD.n11424 VDD.n11419 0.193
R11053 VDD.n11416 VDD.n11411 0.193
R11054 VDD.n11226 VDD.n11221 0.193
R11055 VDD.n11218 VDD.n11213 0.193
R11056 VDD.n12299 VDD.n12293 0.193
R11057 VDD.n12290 VDD.n12285 0.193
R11058 VDD.n2776 VDD.n2775 0.191
R11059 VDD.n3001 VDD.n2994 0.191
R11060 VDD.n3013 VDD.n3006 0.191
R11061 VDD.n3102 VDD.n3101 0.191
R11062 VDD.n3120 VDD.n3119 0.191
R11063 VDD.n3238 VDD.n3232 0.191
R11064 VDD.n3250 VDD.n3243 0.191
R11065 VDD.n3340 VDD.n3339 0.191
R11066 VDD.n3358 VDD.n3357 0.191
R11067 VDD.n3476 VDD.n3469 0.191
R11068 VDD.n3488 VDD.n3481 0.191
R11069 VDD.n3577 VDD.n3576 0.191
R11070 VDD.n3595 VDD.n3594 0.191
R11071 VDD.n3713 VDD.n3707 0.191
R11072 VDD.n3725 VDD.n3718 0.191
R11073 VDD.n3815 VDD.n3814 0.191
R11074 VDD.n3833 VDD.n3832 0.191
R11075 VDD.n3951 VDD.n3944 0.191
R11076 VDD.n3963 VDD.n3956 0.191
R11077 VDD.n4052 VDD.n4051 0.191
R11078 VDD.n4070 VDD.n4069 0.191
R11079 VDD.n4188 VDD.n4182 0.191
R11080 VDD.n4200 VDD.n4193 0.191
R11081 VDD.n4290 VDD.n4289 0.191
R11082 VDD.n4308 VDD.n4307 0.191
R11083 VDD.n4426 VDD.n4419 0.191
R11084 VDD.n4438 VDD.n4431 0.191
R11085 VDD.n5494 VDD.n5493 0.189
R11086 VDD.n5510 VDD.n5509 0.189
R11087 VDD.n5855 VDD.n5854 0.189
R11088 VDD.n5871 VDD.n5870 0.189
R11089 VDD.n6217 VDD.n6216 0.189
R11090 VDD.n6233 VDD.n6232 0.189
R11091 VDD.n6579 VDD.n6578 0.189
R11092 VDD.n6595 VDD.n6594 0.189
R11093 VDD.n6941 VDD.n6940 0.189
R11094 VDD.n6957 VDD.n6956 0.189
R11095 VDD.n7303 VDD.n7302 0.189
R11096 VDD.n7319 VDD.n7318 0.189
R11097 VDD.n7665 VDD.n7664 0.189
R11098 VDD.n7681 VDD.n7680 0.189
R11099 VDD.n8027 VDD.n8026 0.189
R11100 VDD.n8043 VDD.n8042 0.189
R11101 VDD.n8389 VDD.n8388 0.189
R11102 VDD.n8405 VDD.n8404 0.189
R11103 VDD.n8751 VDD.n8750 0.189
R11104 VDD.n8767 VDD.n8766 0.189
R11105 VDD.n9113 VDD.n9112 0.189
R11106 VDD.n9129 VDD.n9128 0.189
R11107 VDD.n9475 VDD.n9474 0.189
R11108 VDD.n9491 VDD.n9490 0.189
R11109 VDD.n9837 VDD.n9836 0.189
R11110 VDD.n9853 VDD.n9852 0.189
R11111 VDD.n12230 VDD.n12229 0.185
R11112 VDD.n2853 VDD.n2852 0.183
R11113 VDD.n2895 VDD.n2881 0.183
R11114 VDD.n4480 VDD.n4476 0.181
R11115 VDD.n4484 VDD.n4483 0.181
R11116 VDD.n4517 VDD.n4516 0.181
R11117 VDD.n4569 VDD.n4568 0.181
R11118 VDD.n255 VDD.n235 0.17
R11119 VDD.n309 VDD.n302 0.17
R11120 VDD.n348 VDD.n347 0.17
R11121 VDD.n5000 VDD.n4996 0.168
R11122 VDD.n4894 VDD.n4884 0.168
R11123 VDD.n4884 VDD.n4880 0.168
R11124 VDD.n4769 VDD.n4765 0.168
R11125 VDD.n4663 VDD.n4653 0.168
R11126 VDD.n4653 VDD.n4649 0.168
R11127 VDD.n2794 VDD.n2789 0.168
R11128 VDD.n3014 VDD.n3002 0.168
R11129 VDD.n3118 VDD.n3114 0.168
R11130 VDD.n3251 VDD.n3239 0.168
R11131 VDD.n3356 VDD.n3352 0.168
R11132 VDD.n3489 VDD.n3477 0.168
R11133 VDD.n3593 VDD.n3589 0.168
R11134 VDD.n3726 VDD.n3714 0.168
R11135 VDD.n3831 VDD.n3827 0.168
R11136 VDD.n3964 VDD.n3952 0.168
R11137 VDD.n4068 VDD.n4064 0.168
R11138 VDD.n4201 VDD.n4189 0.168
R11139 VDD.n4306 VDD.n4302 0.168
R11140 VDD.n4439 VDD.n4427 0.168
R11141 VDD.n225 VDD.n217 0.168
R11142 VDD.n226 VDD.n225 0.168
R11143 VDD.n434 VDD.n422 0.168
R11144 VDD.n542 VDD.n534 0.168
R11145 VDD.n543 VDD.n542 0.168
R11146 VDD.n667 VDD.n655 0.168
R11147 VDD.n776 VDD.n768 0.168
R11148 VDD.n777 VDD.n776 0.168
R11149 VDD.n901 VDD.n889 0.168
R11150 VDD.n1009 VDD.n1001 0.168
R11151 VDD.n1010 VDD.n1009 0.168
R11152 VDD.n1134 VDD.n1122 0.168
R11153 VDD.n1243 VDD.n1235 0.168
R11154 VDD.n1244 VDD.n1243 0.168
R11155 VDD.n1368 VDD.n1356 0.168
R11156 VDD.n1476 VDD.n1468 0.168
R11157 VDD.n1477 VDD.n1476 0.168
R11158 VDD.n1601 VDD.n1589 0.168
R11159 VDD.n1710 VDD.n1702 0.168
R11160 VDD.n1711 VDD.n1710 0.168
R11161 VDD.n1835 VDD.n1823 0.168
R11162 VDD.n2049 VDD.n2045 0.168
R11163 VDD.n2059 VDD.n2049 0.168
R11164 VDD.n2165 VDD.n2161 0.168
R11165 VDD.n2280 VDD.n2276 0.168
R11166 VDD.n2290 VDD.n2280 0.168
R11167 VDD.n2396 VDD.n2392 0.168
R11168 VDD.n5468 VDD.n5467 0.166
R11169 VDD.n5600 VDD.n5599 0.166
R11170 VDD.n5829 VDD.n5828 0.166
R11171 VDD.n5961 VDD.n5960 0.166
R11172 VDD.n6191 VDD.n6190 0.166
R11173 VDD.n6323 VDD.n6322 0.166
R11174 VDD.n6553 VDD.n6552 0.166
R11175 VDD.n6685 VDD.n6684 0.166
R11176 VDD.n6915 VDD.n6914 0.166
R11177 VDD.n7047 VDD.n7046 0.166
R11178 VDD.n7277 VDD.n7276 0.166
R11179 VDD.n7409 VDD.n7408 0.166
R11180 VDD.n7639 VDD.n7638 0.166
R11181 VDD.n7771 VDD.n7770 0.166
R11182 VDD.n8001 VDD.n8000 0.166
R11183 VDD.n8133 VDD.n8132 0.166
R11184 VDD.n8363 VDD.n8362 0.166
R11185 VDD.n8495 VDD.n8494 0.166
R11186 VDD.n8725 VDD.n8724 0.166
R11187 VDD.n8857 VDD.n8856 0.166
R11188 VDD.n9087 VDD.n9086 0.166
R11189 VDD.n9219 VDD.n9218 0.166
R11190 VDD.n9449 VDD.n9448 0.166
R11191 VDD.n9581 VDD.n9580 0.166
R11192 VDD.n9811 VDD.n9810 0.166
R11193 VDD.n9943 VDD.n9942 0.166
R11194 VDD.n1854 VDD.n1853 0.164
R11195 VDD.n1866 VDD.n1857 0.164
R11196 VDD.n1866 VDD.n1859 0.164
R11197 VDD.n1873 VDD.n1871 0.164
R11198 VDD.n1922 VDD.n1912 0.164
R11199 VDD.n1922 VDD.n1915 0.164
R11200 VDD.n10297 VDD.n10289 0.162
R11201 VDD.n10289 VDD.n10285 0.162
R11202 VDD.n10179 VDD.n10171 0.162
R11203 VDD.n10171 VDD.n10167 0.162
R11204 VDD.n10097 VDD.n10088 0.162
R11205 VDD.n10088 VDD.n10084 0.162
R11206 VDD.n10052 VDD.n10044 0.159
R11207 VDD.n10044 VDD.n10040 0.159
R11208 VDD.n10644 VDD.n10636 0.159
R11209 VDD.n10636 VDD.n10632 0.159
R11210 VDD.n10525 VDD.n10517 0.159
R11211 VDD.n10517 VDD.n10513 0.159
R11212 VDD.n2839 VDD.n2832 0.146
R11213 VDD.n2844 VDD.n2843 0.146
R11214 VDD.n2858 VDD.n2854 0.146
R11215 VDD.n2895 VDD.n2888 0.146
R11216 VDD.n2888 VDD.n2887 0.146
R11217 VDD.n2929 VDD.n2928 0.146
R11218 VDD.n4458 VDD.n4457 0.145
R11219 VDD.n4471 VDD.n4464 0.145
R11220 VDD.n4501 VDD.n4500 0.145
R11221 VDD.n4511 VDD.n4501 0.145
R11222 VDD.n4521 VDD.n4518 0.145
R11223 VDD.n4531 VDD.n4524 0.145
R11224 VDD.n4559 VDD.n4540 0.145
R11225 VDD.n4551 VDD.n4550 0.145
R11226 VDD.n10340 VDD.n10339 0.14
R11227 VDD.n10220 VDD.n10219 0.14
R11228 VDD.n10687 VDD.n10686 0.137
R11229 VDD.n10566 VDD.n10565 0.137
R11230 VDD.n260 VDD.n259 0.136
R11231 VDD.n271 VDD.n269 0.136
R11232 VDD.n268 VDD.n267 0.136
R11233 VDD.n267 VDD.n266 0.136
R11234 VDD.n309 VDD.n296 0.136
R11235 VDD.n302 VDD.n301 0.136
R11236 VDD.n10102 VDD.n10101 0.136
R11237 VDD.n10057 VDD.n10056 0.134
R11238 VDD.n421 VDD.n411 0.133
R11239 VDD.n421 VDD.n413 0.133
R11240 VDD.n433 VDD.n424 0.133
R11241 VDD.n433 VDD.n426 0.133
R11242 VDD.n654 VDD.n645 0.133
R11243 VDD.n654 VDD.n647 0.133
R11244 VDD.n666 VDD.n657 0.133
R11245 VDD.n666 VDD.n659 0.133
R11246 VDD.n888 VDD.n878 0.133
R11247 VDD.n888 VDD.n880 0.133
R11248 VDD.n900 VDD.n891 0.133
R11249 VDD.n900 VDD.n893 0.133
R11250 VDD.n1121 VDD.n1112 0.133
R11251 VDD.n1121 VDD.n1114 0.133
R11252 VDD.n1133 VDD.n1124 0.133
R11253 VDD.n1133 VDD.n1126 0.133
R11254 VDD.n1355 VDD.n1345 0.133
R11255 VDD.n1355 VDD.n1347 0.133
R11256 VDD.n1367 VDD.n1358 0.133
R11257 VDD.n1367 VDD.n1360 0.133
R11258 VDD.n1588 VDD.n1579 0.133
R11259 VDD.n1588 VDD.n1581 0.133
R11260 VDD.n1600 VDD.n1591 0.133
R11261 VDD.n1600 VDD.n1593 0.133
R11262 VDD.n1822 VDD.n1812 0.133
R11263 VDD.n1822 VDD.n1814 0.133
R11264 VDD.n1834 VDD.n1825 0.133
R11265 VDD.n1834 VDD.n1827 0.133
R11266 VDD.n5324 VDD.n5323 0.132
R11267 VDD.n5636 VDD.n5635 0.132
R11268 VDD.n5685 VDD.n5684 0.132
R11269 VDD.n5997 VDD.n5996 0.132
R11270 VDD.n6047 VDD.n6046 0.132
R11271 VDD.n6359 VDD.n6358 0.132
R11272 VDD.n6409 VDD.n6408 0.132
R11273 VDD.n6721 VDD.n6720 0.132
R11274 VDD.n6771 VDD.n6770 0.132
R11275 VDD.n7083 VDD.n7082 0.132
R11276 VDD.n7133 VDD.n7132 0.132
R11277 VDD.n7445 VDD.n7444 0.132
R11278 VDD.n7495 VDD.n7494 0.132
R11279 VDD.n7807 VDD.n7806 0.132
R11280 VDD.n7857 VDD.n7856 0.132
R11281 VDD.n8169 VDD.n8168 0.132
R11282 VDD.n8219 VDD.n8218 0.132
R11283 VDD.n8531 VDD.n8530 0.132
R11284 VDD.n8581 VDD.n8580 0.132
R11285 VDD.n8893 VDD.n8892 0.132
R11286 VDD.n8943 VDD.n8942 0.132
R11287 VDD.n9255 VDD.n9254 0.132
R11288 VDD.n9305 VDD.n9304 0.132
R11289 VDD.n9617 VDD.n9616 0.132
R11290 VDD.n9667 VDD.n9666 0.132
R11291 VDD.n9979 VDD.n9978 0.132
R11292 VDD.n1877 VDD.n1876 0.131
R11293 VDD.n1893 VDD.n1892 0.131
R11294 VDD.n1912 VDD.n1910 0.131
R11295 VDD.n1936 VDD.n1935 0.131
R11296 VDD.n200 VDD.n199 0.131
R11297 VDD.n12 VDD.n11 0.127
R11298 VDD.n5071 VDD.n5069 0.127
R11299 VDD.n5057 VDD.n5055 0.127
R11300 VDD.n5043 VDD.n5041 0.127
R11301 VDD.n5029 VDD.n5027 0.127
R11302 VDD.n5015 VDD.n5013 0.127
R11303 VDD.n4992 VDD.n4982 0.127
R11304 VDD.n4978 VDD.n4968 0.127
R11305 VDD.n4964 VDD.n4954 0.127
R11306 VDD.n4950 VDD.n4940 0.127
R11307 VDD.n4936 VDD.n4926 0.127
R11308 VDD.n4922 VDD.n4912 0.127
R11309 VDD.n4908 VDD.n4898 0.127
R11310 VDD.n4868 VDD.n4866 0.127
R11311 VDD.n4854 VDD.n4852 0.127
R11312 VDD.n4840 VDD.n4838 0.127
R11313 VDD.n4826 VDD.n4824 0.127
R11314 VDD.n4812 VDD.n4810 0.127
R11315 VDD.n4798 VDD.n4796 0.127
R11316 VDD.n4784 VDD.n4782 0.127
R11317 VDD.n4761 VDD.n4751 0.127
R11318 VDD.n4747 VDD.n4737 0.127
R11319 VDD.n4733 VDD.n4723 0.127
R11320 VDD.n4719 VDD.n4709 0.127
R11321 VDD.n4705 VDD.n4695 0.127
R11322 VDD.n4691 VDD.n4681 0.127
R11323 VDD.n4677 VDD.n4667 0.127
R11324 VDD.n2809 VDD.n2808 0.127
R11325 VDD.n2841 VDD.n2840 0.127
R11326 VDD.n2867 VDD.n2866 0.127
R11327 VDD.n2897 VDD.n2896 0.127
R11328 VDD.n2916 VDD.n2915 0.127
R11329 VDD.n2963 VDD.n2962 0.127
R11330 VDD.n2977 VDD.n2976 0.127
R11331 VDD.n2991 VDD.n2990 0.127
R11332 VDD.n3028 VDD.n3016 0.127
R11333 VDD.n3042 VDD.n3030 0.127
R11334 VDD.n3056 VDD.n3044 0.127
R11335 VDD.n3070 VDD.n3058 0.127
R11336 VDD.n3084 VDD.n3072 0.127
R11337 VDD.n3098 VDD.n3086 0.127
R11338 VDD.n3112 VDD.n3100 0.127
R11339 VDD.n3130 VDD.n3129 0.127
R11340 VDD.n3144 VDD.n3143 0.127
R11341 VDD.n3159 VDD.n3158 0.127
R11342 VDD.n3173 VDD.n3172 0.127
R11343 VDD.n3187 VDD.n3186 0.127
R11344 VDD.n3201 VDD.n3200 0.127
R11345 VDD.n3215 VDD.n3214 0.127
R11346 VDD.n3229 VDD.n3228 0.127
R11347 VDD.n3265 VDD.n3253 0.127
R11348 VDD.n3279 VDD.n3267 0.127
R11349 VDD.n3293 VDD.n3281 0.127
R11350 VDD.n3307 VDD.n3295 0.127
R11351 VDD.n3322 VDD.n3309 0.127
R11352 VDD.n3336 VDD.n3324 0.127
R11353 VDD.n3350 VDD.n3338 0.127
R11354 VDD.n3368 VDD.n3367 0.127
R11355 VDD.n3382 VDD.n3381 0.127
R11356 VDD.n3396 VDD.n3395 0.127
R11357 VDD.n3410 VDD.n3409 0.127
R11358 VDD.n3424 VDD.n3423 0.127
R11359 VDD.n3438 VDD.n3437 0.127
R11360 VDD.n3452 VDD.n3451 0.127
R11361 VDD.n3466 VDD.n3465 0.127
R11362 VDD.n3503 VDD.n3491 0.127
R11363 VDD.n3517 VDD.n3505 0.127
R11364 VDD.n3531 VDD.n3519 0.127
R11365 VDD.n3545 VDD.n3533 0.127
R11366 VDD.n3559 VDD.n3547 0.127
R11367 VDD.n3573 VDD.n3561 0.127
R11368 VDD.n3587 VDD.n3575 0.127
R11369 VDD.n3605 VDD.n3604 0.127
R11370 VDD.n3619 VDD.n3618 0.127
R11371 VDD.n3634 VDD.n3633 0.127
R11372 VDD.n3648 VDD.n3647 0.127
R11373 VDD.n3662 VDD.n3661 0.127
R11374 VDD.n3676 VDD.n3675 0.127
R11375 VDD.n3690 VDD.n3689 0.127
R11376 VDD.n3704 VDD.n3703 0.127
R11377 VDD.n3740 VDD.n3728 0.127
R11378 VDD.n3754 VDD.n3742 0.127
R11379 VDD.n3768 VDD.n3756 0.127
R11380 VDD.n3782 VDD.n3770 0.127
R11381 VDD.n3797 VDD.n3784 0.127
R11382 VDD.n3811 VDD.n3799 0.127
R11383 VDD.n3825 VDD.n3813 0.127
R11384 VDD.n3843 VDD.n3842 0.127
R11385 VDD.n3857 VDD.n3856 0.127
R11386 VDD.n3871 VDD.n3870 0.127
R11387 VDD.n3885 VDD.n3884 0.127
R11388 VDD.n3899 VDD.n3898 0.127
R11389 VDD.n3913 VDD.n3912 0.127
R11390 VDD.n3927 VDD.n3926 0.127
R11391 VDD.n3941 VDD.n3940 0.127
R11392 VDD.n3978 VDD.n3966 0.127
R11393 VDD.n3992 VDD.n3980 0.127
R11394 VDD.n4006 VDD.n3994 0.127
R11395 VDD.n4020 VDD.n4008 0.127
R11396 VDD.n4034 VDD.n4022 0.127
R11397 VDD.n4048 VDD.n4036 0.127
R11398 VDD.n4062 VDD.n4050 0.127
R11399 VDD.n4080 VDD.n4079 0.127
R11400 VDD.n4094 VDD.n4093 0.127
R11401 VDD.n4109 VDD.n4108 0.127
R11402 VDD.n4123 VDD.n4122 0.127
R11403 VDD.n4137 VDD.n4136 0.127
R11404 VDD.n4151 VDD.n4150 0.127
R11405 VDD.n4165 VDD.n4164 0.127
R11406 VDD.n4179 VDD.n4178 0.127
R11407 VDD.n4215 VDD.n4203 0.127
R11408 VDD.n4229 VDD.n4217 0.127
R11409 VDD.n4243 VDD.n4231 0.127
R11410 VDD.n4257 VDD.n4245 0.127
R11411 VDD.n4272 VDD.n4259 0.127
R11412 VDD.n4286 VDD.n4274 0.127
R11413 VDD.n4300 VDD.n4288 0.127
R11414 VDD.n4318 VDD.n4317 0.127
R11415 VDD.n4332 VDD.n4331 0.127
R11416 VDD.n4346 VDD.n4345 0.127
R11417 VDD.n4360 VDD.n4359 0.127
R11418 VDD.n4374 VDD.n4373 0.127
R11419 VDD.n4388 VDD.n4387 0.127
R11420 VDD.n4402 VDD.n4401 0.127
R11421 VDD.n4416 VDD.n4415 0.127
R11422 VDD.n4453 VDD.n4441 0.127
R11423 VDD.n4472 VDD.n4455 0.127
R11424 VDD.n4492 VDD.n4474 0.127
R11425 VDD.n4512 VDD.n4494 0.127
R11426 VDD.n4532 VDD.n4514 0.127
R11427 VDD.n4560 VDD.n4534 0.127
R11428 VDD.n4623 VDD.n4562 0.127
R11429 VDD.n257 VDD.n256 0.127
R11430 VDD.n280 VDD.n279 0.127
R11431 VDD.n311 VDD.n310 0.127
R11432 VDD.n329 VDD.n328 0.127
R11433 VDD.n380 VDD.n379 0.127
R11434 VDD.n394 VDD.n393 0.127
R11435 VDD.n408 VDD.n407 0.127
R11436 VDD.n448 VDD.n436 0.127
R11437 VDD.n462 VDD.n450 0.127
R11438 VDD.n476 VDD.n464 0.127
R11439 VDD.n490 VDD.n478 0.127
R11440 VDD.n504 VDD.n492 0.127
R11441 VDD.n518 VDD.n506 0.127
R11442 VDD.n532 VDD.n520 0.127
R11443 VDD.n557 VDD.n556 0.127
R11444 VDD.n572 VDD.n571 0.127
R11445 VDD.n586 VDD.n585 0.127
R11446 VDD.n600 VDD.n599 0.127
R11447 VDD.n614 VDD.n613 0.127
R11448 VDD.n628 VDD.n627 0.127
R11449 VDD.n642 VDD.n641 0.127
R11450 VDD.n681 VDD.n669 0.127
R11451 VDD.n695 VDD.n683 0.127
R11452 VDD.n709 VDD.n697 0.127
R11453 VDD.n723 VDD.n711 0.127
R11454 VDD.n738 VDD.n725 0.127
R11455 VDD.n752 VDD.n740 0.127
R11456 VDD.n766 VDD.n754 0.127
R11457 VDD.n791 VDD.n790 0.127
R11458 VDD.n805 VDD.n804 0.127
R11459 VDD.n819 VDD.n818 0.127
R11460 VDD.n833 VDD.n832 0.127
R11461 VDD.n847 VDD.n846 0.127
R11462 VDD.n861 VDD.n860 0.127
R11463 VDD.n875 VDD.n874 0.127
R11464 VDD.n915 VDD.n903 0.127
R11465 VDD.n929 VDD.n917 0.127
R11466 VDD.n943 VDD.n931 0.127
R11467 VDD.n957 VDD.n945 0.127
R11468 VDD.n971 VDD.n959 0.127
R11469 VDD.n985 VDD.n973 0.127
R11470 VDD.n999 VDD.n987 0.127
R11471 VDD.n1024 VDD.n1023 0.127
R11472 VDD.n1039 VDD.n1038 0.127
R11473 VDD.n1053 VDD.n1052 0.127
R11474 VDD.n1067 VDD.n1066 0.127
R11475 VDD.n1081 VDD.n1080 0.127
R11476 VDD.n1095 VDD.n1094 0.127
R11477 VDD.n1109 VDD.n1108 0.127
R11478 VDD.n1148 VDD.n1136 0.127
R11479 VDD.n1162 VDD.n1150 0.127
R11480 VDD.n1176 VDD.n1164 0.127
R11481 VDD.n1190 VDD.n1178 0.127
R11482 VDD.n1205 VDD.n1192 0.127
R11483 VDD.n1219 VDD.n1207 0.127
R11484 VDD.n1233 VDD.n1221 0.127
R11485 VDD.n1258 VDD.n1257 0.127
R11486 VDD.n1272 VDD.n1271 0.127
R11487 VDD.n1286 VDD.n1285 0.127
R11488 VDD.n1300 VDD.n1299 0.127
R11489 VDD.n1314 VDD.n1313 0.127
R11490 VDD.n1328 VDD.n1327 0.127
R11491 VDD.n1342 VDD.n1341 0.127
R11492 VDD.n1382 VDD.n1370 0.127
R11493 VDD.n1396 VDD.n1384 0.127
R11494 VDD.n1410 VDD.n1398 0.127
R11495 VDD.n1424 VDD.n1412 0.127
R11496 VDD.n1438 VDD.n1426 0.127
R11497 VDD.n1452 VDD.n1440 0.127
R11498 VDD.n1466 VDD.n1454 0.127
R11499 VDD.n1491 VDD.n1490 0.127
R11500 VDD.n1506 VDD.n1505 0.127
R11501 VDD.n1520 VDD.n1519 0.127
R11502 VDD.n1534 VDD.n1533 0.127
R11503 VDD.n1548 VDD.n1547 0.127
R11504 VDD.n1562 VDD.n1561 0.127
R11505 VDD.n1576 VDD.n1575 0.127
R11506 VDD.n1615 VDD.n1603 0.127
R11507 VDD.n1629 VDD.n1617 0.127
R11508 VDD.n1643 VDD.n1631 0.127
R11509 VDD.n1657 VDD.n1645 0.127
R11510 VDD.n1672 VDD.n1659 0.127
R11511 VDD.n1686 VDD.n1674 0.127
R11512 VDD.n1700 VDD.n1688 0.127
R11513 VDD.n1725 VDD.n1724 0.127
R11514 VDD.n1739 VDD.n1738 0.127
R11515 VDD.n1753 VDD.n1752 0.127
R11516 VDD.n1767 VDD.n1766 0.127
R11517 VDD.n1781 VDD.n1780 0.127
R11518 VDD.n1795 VDD.n1794 0.127
R11519 VDD.n1809 VDD.n1808 0.127
R11520 VDD.n1849 VDD.n1837 0.127
R11521 VDD.n1867 VDD.n1851 0.127
R11522 VDD.n1885 VDD.n1869 0.127
R11523 VDD.n1904 VDD.n1887 0.127
R11524 VDD.n1923 VDD.n1906 0.127
R11525 VDD.n1945 VDD.n1925 0.127
R11526 VDD.n2018 VDD.n1947 0.127
R11527 VDD.n2073 VDD.n2063 0.127
R11528 VDD.n2087 VDD.n2077 0.127
R11529 VDD.n2101 VDD.n2091 0.127
R11530 VDD.n2115 VDD.n2105 0.127
R11531 VDD.n2129 VDD.n2119 0.127
R11532 VDD.n2143 VDD.n2133 0.127
R11533 VDD.n2157 VDD.n2147 0.127
R11534 VDD.n2180 VDD.n2178 0.127
R11535 VDD.n2194 VDD.n2192 0.127
R11536 VDD.n2208 VDD.n2206 0.127
R11537 VDD.n2222 VDD.n2220 0.127
R11538 VDD.n2236 VDD.n2234 0.127
R11539 VDD.n2250 VDD.n2248 0.127
R11540 VDD.n2264 VDD.n2262 0.127
R11541 VDD.n2304 VDD.n2294 0.127
R11542 VDD.n2318 VDD.n2308 0.127
R11543 VDD.n2332 VDD.n2322 0.127
R11544 VDD.n2346 VDD.n2336 0.127
R11545 VDD.n2360 VDD.n2350 0.127
R11546 VDD.n2374 VDD.n2364 0.127
R11547 VDD.n2388 VDD.n2378 0.127
R11548 VDD.n2411 VDD.n2409 0.127
R11549 VDD.n2425 VDD.n2423 0.127
R11550 VDD.n2439 VDD.n2437 0.127
R11551 VDD.n2453 VDD.n2451 0.127
R11552 VDD.n2467 VDD.n2465 0.127
R11553 VDD.n12243 VDD.n12242 0.127
R11554 VDD.n10335 VDD.n10326 0.122
R11555 VDD.n10322 VDD.n10314 0.122
R11556 VDD.n10310 VDD.n10301 0.122
R11557 VDD.n10274 VDD.n10272 0.122
R11558 VDD.n10262 VDD.n10260 0.122
R11559 VDD.n10249 VDD.n10247 0.122
R11560 VDD.n10215 VDD.n10207 0.122
R11561 VDD.n10203 VDD.n10195 0.122
R11562 VDD.n10191 VDD.n10183 0.122
R11563 VDD.n10157 VDD.n10155 0.122
R11564 VDD.n10145 VDD.n10143 0.122
R11565 VDD.n10133 VDD.n10131 0.122
R11566 VDD.n5321 VDD.n5320 0.121
R11567 VDD.n5646 VDD.n5645 0.121
R11568 VDD.n5682 VDD.n5681 0.121
R11569 VDD.n6007 VDD.n6006 0.121
R11570 VDD.n6044 VDD.n6043 0.121
R11571 VDD.n6369 VDD.n6368 0.121
R11572 VDD.n6406 VDD.n6405 0.121
R11573 VDD.n6731 VDD.n6730 0.121
R11574 VDD.n6768 VDD.n6767 0.121
R11575 VDD.n7093 VDD.n7092 0.121
R11576 VDD.n7130 VDD.n7129 0.121
R11577 VDD.n7455 VDD.n7454 0.121
R11578 VDD.n7492 VDD.n7491 0.121
R11579 VDD.n7817 VDD.n7816 0.121
R11580 VDD.n7854 VDD.n7853 0.121
R11581 VDD.n8179 VDD.n8178 0.121
R11582 VDD.n8216 VDD.n8215 0.121
R11583 VDD.n8541 VDD.n8540 0.121
R11584 VDD.n8578 VDD.n8577 0.121
R11585 VDD.n8903 VDD.n8902 0.121
R11586 VDD.n8940 VDD.n8939 0.121
R11587 VDD.n9265 VDD.n9264 0.121
R11588 VDD.n9302 VDD.n9301 0.121
R11589 VDD.n9627 VDD.n9626 0.121
R11590 VDD.n9664 VDD.n9663 0.121
R11591 VDD.n9989 VDD.n9988 0.121
R11592 VDD.n10682 VDD.n10673 0.12
R11593 VDD.n10669 VDD.n10661 0.12
R11594 VDD.n10657 VDD.n10648 0.12
R11595 VDD.n10621 VDD.n10619 0.12
R11596 VDD.n10609 VDD.n10607 0.12
R11597 VDD.n10596 VDD.n10594 0.12
R11598 VDD.n10561 VDD.n10553 0.12
R11599 VDD.n10549 VDD.n10541 0.12
R11600 VDD.n10537 VDD.n10529 0.12
R11601 VDD.n10503 VDD.n10501 0.12
R11602 VDD.n10491 VDD.n10489 0.12
R11603 VDD.n10479 VDD.n10477 0.12
R11604 VDD.n2865 VDD.n2850 0.11
R11605 VDD.n2852 VDD.n2851 0.11
R11606 VDD.n2961 VDD.n2929 0.11
R11607 VDD.n2951 VDD.n2931 0.11
R11608 VDD.n4504 VDD.n4503 0.109
R11609 VDD.n69 VDD.n60 0.108
R11610 VDD.n12300 VDD.n12291 0.105
R11611 VDD.n4602 VDD.n4601 0.1
R11612 VDD.n4611 VDD.n4610 0.1
R11613 VDD.n2814 VDD.n2813 0.1
R11614 VDD.n2946 VDD.n2945 0.1
R11615 VDD.n238 VDD.n237 0.1
R11616 VDD.n363 VDD.n362 0.1
R11617 VDD.n1996 VDD.n1995 0.1
R11618 VDD.n2005 VDD.n2004 0.1
R11619 VDD.n10895 VDD.n10894 0.1
R11620 VDD.n10721 VDD.n10720 0.1
R11621 VDD.n11664 VDD.n11663 0.1
R11622 VDD.n11491 VDD.n11490 0.1
R11623 VDD.n1871 VDD.n1870 0.098
R11624 VDD.n1884 VDD.n1877 0.098
R11625 VDD.n1903 VDD.n1893 0.098
R11626 VDD.n1927 VDD.n1926 0.098
R11627 VDD.n1944 VDD.n1934 0.098
R11628 VDD.n1944 VDD.n1937 0.098
R11629 VDD.n87 VDD.n86 0.091
R11630 VDD.n10012 VDD.n9650 0.09
R11631 VDD.n9650 VDD.n9288 0.09
R11632 VDD.n9288 VDD.n8926 0.09
R11633 VDD.n8926 VDD.n8564 0.09
R11634 VDD.n8564 VDD.n8202 0.09
R11635 VDD.n8202 VDD.n7840 0.09
R11636 VDD.n7840 VDD.n7478 0.09
R11637 VDD.n7478 VDD.n7116 0.09
R11638 VDD.n7116 VDD.n6754 0.09
R11639 VDD.n6754 VDD.n6392 0.09
R11640 VDD.n6392 VDD.n6030 0.09
R11641 VDD.n10422 VDD.n10421 0.09
R11642 VDD.n12318 VDD.n12317 0.089
R11643 VDD.n12229 VDD.n11462 0.087
R11644 VDD.n67 VDD.n66 0.087
R11645 VDD.n58 VDD.n57 0.087
R11646 VDD.n11934 VDD.n11933 0.087
R11647 VDD.n11423 VDD.n11422 0.087
R11648 VDD.n11225 VDD.n11224 0.087
R11649 VDD.n12298 VDD.n12297 0.087
R11650 VDD.n12289 VDD.n12288 0.087
R11651 VDD.n10430 VDD.n10429 0.085
R11652 VDD.n10404 VDD.n10403 0.085
R11653 VDD.n10377 VDD.n10376 0.085
R11654 VDD.n10348 VDD.n10347 0.085
R11655 VDD.n82 VDD.n73 0.081
R11656 VDD.n50 VDD.n48 0.081
R11657 VDD.n10368 VDD.n10367 0.079
R11658 VDD.n10395 VDD.n10394 0.079
R11659 VDD.n11576 VDD.n11575 0.079
R11660 VDD.n11573 VDD.n11572 0.079
R11661 VDD.n11559 VDD.n11558 0.079
R11662 VDD.n11556 VDD.n11555 0.079
R11663 VDD.n11730 VDD.n11729 0.079
R11664 VDD.n11733 VDD.n11732 0.079
R11665 VDD.n11747 VDD.n11746 0.079
R11666 VDD.n10806 VDD.n10805 0.079
R11667 VDD.n10803 VDD.n10802 0.079
R11668 VDD.n10789 VDD.n10788 0.079
R11669 VDD.n10786 VDD.n10785 0.079
R11670 VDD.n10961 VDD.n10960 0.079
R11671 VDD.n10964 VDD.n10963 0.079
R11672 VDD.n10978 VDD.n10977 0.079
R11673 VDD.n12313 VDD.n12304 0.079
R11674 VDD.n12281 VDD.n12279 0.079
R11675 VDD VDD.n12230 0.078
R11676 VDD.n2480 VDD.n2479 0.077
R11677 VDD.n5084 VDD.n5083 0.076
R11678 VDD.n2812 VDD.n2811 0.073
R11679 VDD.n2828 VDD.n2827 0.073
R11680 VDD.n2854 VDD.n2853 0.073
R11681 VDD.n2887 VDD.n2884 0.073
R11682 VDD.n2907 VDD.n2906 0.073
R11683 VDD.n4476 VDD.n4475 0.072
R11684 VDD.n4481 VDD.n4480 0.072
R11685 VDD.n4491 VDD.n4484 0.072
R11686 VDD.n4500 VDD.n4496 0.072
R11687 VDD.n4516 VDD.n4515 0.072
R11688 VDD.n4518 VDD.n4517 0.072
R11689 VDD.n4536 VDD.n4535 0.072
R11690 VDD.n4559 VDD.n4552 0.072
R11691 VDD.n4568 VDD.n4567 0.072
R11692 VDD.n12197 VDD.n12188 0.072
R11693 VDD.n12090 VDD.n12088 0.072
R11694 VDD.n12088 VDD.n12084 0.072
R11695 VDD.n11993 VDD.n11984 0.072
R11696 VDD.n11425 VDD.n11417 0.072
R11697 VDD.n11321 VDD.n11319 0.072
R11698 VDD.n11319 VDD.n11315 0.072
R11699 VDD.n11227 VDD.n11219 0.072
R11700 VDD.n5307 VDD.n5306 0.071
R11701 VDD.n11136 VDD.n11135 0.071
R11702 VDD.n11885 VDD.n11884 0.071
R11703 VDD.n10689 VDD.n10688 0.069
R11704 VDD.n11072 VDD.n11071 0.068
R11705 VDD.n11838 VDD.n11837 0.068
R11706 VDD.n334 VDD.n333 0.068
R11707 VDD.n229 VDD.n228 0.068
R11708 VDD.n231 VDD.n230 0.068
R11709 VDD.n278 VDD.n265 0.068
R11710 VDD.n269 VDD.n268 0.068
R11711 VDD.n301 VDD.n299 0.068
R11712 VDD.n298 VDD.n297 0.068
R11713 VDD.n320 VDD.n319 0.068
R11714 VDD.n378 VDD.n348 0.068
R11715 VDD.n368 VDD.n350 0.068
R11716 VDD.n11769 VDD.n11768 0.067
R11717 VDD.n11001 VDD.n11000 0.067
R11718 VDD.n11939 VDD.n11938 0.066
R11719 VDD.n11182 VDD.n11181 0.065
R11720 VDD.n1874 VDD.n1873 0.065
R11721 VDD.n1892 VDD.n1890 0.065
R11722 VDD.n1896 VDD.n1895 0.065
R11723 VDD.n1910 VDD.n1909 0.065
R11724 VDD.n201 VDD.n200 0.065
R11725 VDD.n11182 VDD.n11153 0.065
R11726 VDD.n11939 VDD.n11911 0.064
R11727 VDD.n12226 VDD.n12225 0.063
R11728 VDD.n11459 VDD.n11453 0.063
R11729 VDD.n12320 VDD.n12319 0.056
R11730 VDD.n4605 VDD.n4604 0.055
R11731 VDD.n4607 VDD.n4606 0.055
R11732 VDD.n4608 VDD.n4607 0.055
R11733 VDD.n2940 VDD.n2939 0.055
R11734 VDD.n2942 VDD.n2941 0.055
R11735 VDD.n2943 VDD.n2942 0.055
R11736 VDD.n357 VDD.n356 0.055
R11737 VDD.n359 VDD.n358 0.055
R11738 VDD.n360 VDD.n359 0.055
R11739 VDD.n1999 VDD.n1998 0.055
R11740 VDD.n2001 VDD.n2000 0.055
R11741 VDD.n2002 VDD.n2001 0.055
R11742 VDD.n12221 VDD.n12213 0.055
R11743 VDD.n12209 VDD.n12201 0.055
R11744 VDD.n12177 VDD.n12175 0.055
R11745 VDD.n12165 VDD.n12163 0.055
R11746 VDD.n12152 VDD.n12150 0.055
R11747 VDD.n12140 VDD.n12138 0.055
R11748 VDD.n12127 VDD.n12125 0.055
R11749 VDD.n12115 VDD.n12113 0.055
R11750 VDD.n12102 VDD.n12100 0.055
R11751 VDD.n12080 VDD.n12072 0.055
R11752 VDD.n12068 VDD.n12059 0.055
R11753 VDD.n12055 VDD.n12047 0.055
R11754 VDD.n12043 VDD.n12034 0.055
R11755 VDD.n12030 VDD.n12022 0.055
R11756 VDD.n12018 VDD.n12009 0.055
R11757 VDD.n12005 VDD.n11997 0.055
R11758 VDD.n11973 VDD.n11971 0.055
R11759 VDD.n11449 VDD.n11441 0.055
R11760 VDD.n11437 VDD.n11429 0.055
R11761 VDD.n11407 VDD.n11405 0.055
R11762 VDD.n11395 VDD.n11393 0.055
R11763 VDD.n11383 VDD.n11381 0.055
R11764 VDD.n11371 VDD.n11369 0.055
R11765 VDD.n11359 VDD.n11357 0.055
R11766 VDD.n11347 VDD.n11345 0.055
R11767 VDD.n11335 VDD.n11333 0.055
R11768 VDD.n11311 VDD.n11303 0.055
R11769 VDD.n11299 VDD.n11291 0.055
R11770 VDD.n11287 VDD.n11279 0.055
R11771 VDD.n11275 VDD.n11267 0.055
R11772 VDD.n11263 VDD.n11255 0.055
R11773 VDD.n11251 VDD.n11243 0.055
R11774 VDD.n11239 VDD.n11231 0.055
R11775 VDD.n11209 VDD.n11207 0.055
R11776 VDD.n11882 VDD.n11880 0.054
R11777 VDD.n11926 VDD.n11925 0.054
R11778 VDD.n11168 VDD.n11167 0.053
R11779 VDD.n4606 VDD.n4605 0.052
R11780 VDD.n2941 VDD.n2940 0.052
R11781 VDD.n358 VDD.n357 0.052
R11782 VDD.n2000 VDD.n1999 0.052
R11783 VDD.n89 VDD.n88 0.052
R11784 VDD.n11140 VDD.n11139 0.052
R11785 VDD.n11899 VDD.n11898 0.052
R11786 VDD.n5529 VDD.n5464 0.049
R11787 VDD.n5415 VDD.n5406 0.049
R11788 VDD.n5460 VDD.n5451 0.049
R11789 VDD.n5564 VDD.n5558 0.049
R11790 VDD.n5890 VDD.n5825 0.049
R11791 VDD.n5776 VDD.n5767 0.049
R11792 VDD.n5821 VDD.n5812 0.049
R11793 VDD.n5925 VDD.n5919 0.049
R11794 VDD.n6252 VDD.n6187 0.049
R11795 VDD.n6138 VDD.n6129 0.049
R11796 VDD.n6183 VDD.n6174 0.049
R11797 VDD.n6287 VDD.n6281 0.049
R11798 VDD.n6614 VDD.n6549 0.049
R11799 VDD.n6500 VDD.n6491 0.049
R11800 VDD.n6545 VDD.n6536 0.049
R11801 VDD.n6649 VDD.n6643 0.049
R11802 VDD.n6976 VDD.n6911 0.049
R11803 VDD.n6862 VDD.n6853 0.049
R11804 VDD.n6907 VDD.n6898 0.049
R11805 VDD.n7011 VDD.n7005 0.049
R11806 VDD.n7338 VDD.n7273 0.049
R11807 VDD.n7224 VDD.n7215 0.049
R11808 VDD.n7269 VDD.n7260 0.049
R11809 VDD.n7373 VDD.n7367 0.049
R11810 VDD.n7700 VDD.n7635 0.049
R11811 VDD.n7586 VDD.n7577 0.049
R11812 VDD.n7631 VDD.n7622 0.049
R11813 VDD.n7735 VDD.n7729 0.049
R11814 VDD.n8062 VDD.n7997 0.049
R11815 VDD.n7948 VDD.n7939 0.049
R11816 VDD.n7993 VDD.n7984 0.049
R11817 VDD.n8097 VDD.n8091 0.049
R11818 VDD.n8424 VDD.n8359 0.049
R11819 VDD.n8310 VDD.n8301 0.049
R11820 VDD.n8355 VDD.n8346 0.049
R11821 VDD.n8459 VDD.n8453 0.049
R11822 VDD.n8786 VDD.n8721 0.049
R11823 VDD.n8672 VDD.n8663 0.049
R11824 VDD.n8717 VDD.n8708 0.049
R11825 VDD.n8821 VDD.n8815 0.049
R11826 VDD.n9148 VDD.n9083 0.049
R11827 VDD.n9034 VDD.n9025 0.049
R11828 VDD.n9079 VDD.n9070 0.049
R11829 VDD.n9183 VDD.n9177 0.049
R11830 VDD.n9510 VDD.n9445 0.049
R11831 VDD.n9396 VDD.n9387 0.049
R11832 VDD.n9441 VDD.n9432 0.049
R11833 VDD.n9545 VDD.n9539 0.049
R11834 VDD.n9872 VDD.n9807 0.049
R11835 VDD.n9758 VDD.n9749 0.049
R11836 VDD.n9803 VDD.n9794 0.049
R11837 VDD.n9907 VDD.n9901 0.049
R11838 VDD.n11141 VDD.n11140 0.048
R11839 VDD.n11900 VDD.n11899 0.048
R11840 VDD.n4574 VDD.n4573 0.048
R11841 VDD.n4579 VDD.n4578 0.048
R11842 VDD.n4592 VDD.n4591 0.048
R11843 VDD.n4597 VDD.n4596 0.048
R11844 VDD.n2821 VDD.n2820 0.048
R11845 VDD.n2846 VDD.n2845 0.048
R11846 VDD.n2875 VDD.n2874 0.048
R11847 VDD.n2936 VDD.n2935 0.048
R11848 VDD.n245 VDD.n244 0.048
R11849 VDD.n262 VDD.n261 0.048
R11850 VDD.n290 VDD.n289 0.048
R11851 VDD.n354 VDD.n353 0.048
R11852 VDD.n1968 VDD.n1967 0.048
R11853 VDD.n1973 VDD.n1972 0.048
R11854 VDD.n1986 VDD.n1985 0.048
R11855 VDD.n1991 VDD.n1990 0.048
R11856 VDD.n11169 VDD.n11168 0.047
R11857 VDD.n2547 VDD.n2546 0.047
R11858 VDD.n135 VDD.n134 0.047
R11859 VDD.n152 VDD.n151 0.047
R11860 VDD.n5169 VDD.n5168 0.047
R11861 VDD.n2650 VDD.n2649 0.047
R11862 VDD.n2674 VDD.n2673 0.047
R11863 VDD.n2654 VDD.n2653 0.047
R11864 VDD.n5380 VDD.n5379 0.047
R11865 VDD.n5363 VDD.n5361 0.047
R11866 VDD.n5361 VDD.n5360 0.047
R11867 VDD.n5356 VDD.n5354 0.047
R11868 VDD.n5492 VDD.n5491 0.047
R11869 VDD.n5513 VDD.n5512 0.047
R11870 VDD.n5633 VDD.n5631 0.047
R11871 VDD.n5638 VDD.n5637 0.047
R11872 VDD.n5641 VDD.n5639 0.047
R11873 VDD.n5663 VDD.n5662 0.047
R11874 VDD.n5571 VDD.n5569 0.047
R11875 VDD.n5741 VDD.n5740 0.047
R11876 VDD.n5724 VDD.n5722 0.047
R11877 VDD.n5722 VDD.n5721 0.047
R11878 VDD.n5717 VDD.n5715 0.047
R11879 VDD.n5853 VDD.n5852 0.047
R11880 VDD.n5874 VDD.n5873 0.047
R11881 VDD.n5994 VDD.n5992 0.047
R11882 VDD.n5999 VDD.n5998 0.047
R11883 VDD.n6002 VDD.n6000 0.047
R11884 VDD.n6024 VDD.n6023 0.047
R11885 VDD.n5932 VDD.n5930 0.047
R11886 VDD.n6103 VDD.n6102 0.047
R11887 VDD.n6086 VDD.n6084 0.047
R11888 VDD.n6084 VDD.n6083 0.047
R11889 VDD.n6079 VDD.n6077 0.047
R11890 VDD.n6215 VDD.n6214 0.047
R11891 VDD.n6236 VDD.n6235 0.047
R11892 VDD.n6356 VDD.n6354 0.047
R11893 VDD.n6361 VDD.n6360 0.047
R11894 VDD.n6364 VDD.n6362 0.047
R11895 VDD.n6386 VDD.n6385 0.047
R11896 VDD.n6294 VDD.n6292 0.047
R11897 VDD.n6465 VDD.n6464 0.047
R11898 VDD.n6448 VDD.n6446 0.047
R11899 VDD.n6446 VDD.n6445 0.047
R11900 VDD.n6441 VDD.n6439 0.047
R11901 VDD.n6577 VDD.n6576 0.047
R11902 VDD.n6598 VDD.n6597 0.047
R11903 VDD.n6718 VDD.n6716 0.047
R11904 VDD.n6723 VDD.n6722 0.047
R11905 VDD.n6726 VDD.n6724 0.047
R11906 VDD.n6748 VDD.n6747 0.047
R11907 VDD.n6656 VDD.n6654 0.047
R11908 VDD.n6827 VDD.n6826 0.047
R11909 VDD.n6810 VDD.n6808 0.047
R11910 VDD.n6808 VDD.n6807 0.047
R11911 VDD.n6803 VDD.n6801 0.047
R11912 VDD.n6939 VDD.n6938 0.047
R11913 VDD.n6960 VDD.n6959 0.047
R11914 VDD.n7080 VDD.n7078 0.047
R11915 VDD.n7085 VDD.n7084 0.047
R11916 VDD.n7088 VDD.n7086 0.047
R11917 VDD.n7110 VDD.n7109 0.047
R11918 VDD.n7018 VDD.n7016 0.047
R11919 VDD.n7189 VDD.n7188 0.047
R11920 VDD.n7172 VDD.n7170 0.047
R11921 VDD.n7170 VDD.n7169 0.047
R11922 VDD.n7165 VDD.n7163 0.047
R11923 VDD.n7301 VDD.n7300 0.047
R11924 VDD.n7322 VDD.n7321 0.047
R11925 VDD.n7442 VDD.n7440 0.047
R11926 VDD.n7447 VDD.n7446 0.047
R11927 VDD.n7450 VDD.n7448 0.047
R11928 VDD.n7472 VDD.n7471 0.047
R11929 VDD.n7380 VDD.n7378 0.047
R11930 VDD.n7551 VDD.n7550 0.047
R11931 VDD.n7534 VDD.n7532 0.047
R11932 VDD.n7532 VDD.n7531 0.047
R11933 VDD.n7527 VDD.n7525 0.047
R11934 VDD.n7663 VDD.n7662 0.047
R11935 VDD.n7684 VDD.n7683 0.047
R11936 VDD.n7804 VDD.n7802 0.047
R11937 VDD.n7809 VDD.n7808 0.047
R11938 VDD.n7812 VDD.n7810 0.047
R11939 VDD.n7834 VDD.n7833 0.047
R11940 VDD.n7742 VDD.n7740 0.047
R11941 VDD.n7913 VDD.n7912 0.047
R11942 VDD.n7896 VDD.n7894 0.047
R11943 VDD.n7894 VDD.n7893 0.047
R11944 VDD.n7889 VDD.n7887 0.047
R11945 VDD.n8025 VDD.n8024 0.047
R11946 VDD.n8046 VDD.n8045 0.047
R11947 VDD.n8166 VDD.n8164 0.047
R11948 VDD.n8171 VDD.n8170 0.047
R11949 VDD.n8174 VDD.n8172 0.047
R11950 VDD.n8196 VDD.n8195 0.047
R11951 VDD.n8104 VDD.n8102 0.047
R11952 VDD.n8275 VDD.n8274 0.047
R11953 VDD.n8258 VDD.n8256 0.047
R11954 VDD.n8256 VDD.n8255 0.047
R11955 VDD.n8251 VDD.n8249 0.047
R11956 VDD.n8387 VDD.n8386 0.047
R11957 VDD.n8408 VDD.n8407 0.047
R11958 VDD.n8528 VDD.n8526 0.047
R11959 VDD.n8533 VDD.n8532 0.047
R11960 VDD.n8536 VDD.n8534 0.047
R11961 VDD.n8558 VDD.n8557 0.047
R11962 VDD.n8466 VDD.n8464 0.047
R11963 VDD.n8637 VDD.n8636 0.047
R11964 VDD.n8620 VDD.n8618 0.047
R11965 VDD.n8618 VDD.n8617 0.047
R11966 VDD.n8613 VDD.n8611 0.047
R11967 VDD.n8749 VDD.n8748 0.047
R11968 VDD.n8770 VDD.n8769 0.047
R11969 VDD.n8890 VDD.n8888 0.047
R11970 VDD.n8895 VDD.n8894 0.047
R11971 VDD.n8898 VDD.n8896 0.047
R11972 VDD.n8920 VDD.n8919 0.047
R11973 VDD.n8828 VDD.n8826 0.047
R11974 VDD.n8999 VDD.n8998 0.047
R11975 VDD.n8982 VDD.n8980 0.047
R11976 VDD.n8980 VDD.n8979 0.047
R11977 VDD.n8975 VDD.n8973 0.047
R11978 VDD.n9111 VDD.n9110 0.047
R11979 VDD.n9132 VDD.n9131 0.047
R11980 VDD.n9252 VDD.n9250 0.047
R11981 VDD.n9257 VDD.n9256 0.047
R11982 VDD.n9260 VDD.n9258 0.047
R11983 VDD.n9282 VDD.n9281 0.047
R11984 VDD.n9190 VDD.n9188 0.047
R11985 VDD.n9361 VDD.n9360 0.047
R11986 VDD.n9344 VDD.n9342 0.047
R11987 VDD.n9342 VDD.n9341 0.047
R11988 VDD.n9337 VDD.n9335 0.047
R11989 VDD.n9473 VDD.n9472 0.047
R11990 VDD.n9494 VDD.n9493 0.047
R11991 VDD.n9614 VDD.n9612 0.047
R11992 VDD.n9619 VDD.n9618 0.047
R11993 VDD.n9622 VDD.n9620 0.047
R11994 VDD.n9644 VDD.n9643 0.047
R11995 VDD.n9552 VDD.n9550 0.047
R11996 VDD.n9723 VDD.n9722 0.047
R11997 VDD.n9706 VDD.n9704 0.047
R11998 VDD.n9704 VDD.n9703 0.047
R11999 VDD.n9699 VDD.n9697 0.047
R12000 VDD.n9835 VDD.n9834 0.047
R12001 VDD.n9856 VDD.n9855 0.047
R12002 VDD.n9976 VDD.n9974 0.047
R12003 VDD.n9981 VDD.n9980 0.047
R12004 VDD.n9984 VDD.n9982 0.047
R12005 VDD.n10006 VDD.n10005 0.047
R12006 VDD.n9914 VDD.n9912 0.047
R12007 VDD.n11570 VDD.n11569 0.047
R12008 VDD.n11566 VDD.n11565 0.047
R12009 VDD.n11562 VDD.n11561 0.047
R12010 VDD.n11736 VDD.n11735 0.047
R12011 VDD.n11740 VDD.n11739 0.047
R12012 VDD.n11744 VDD.n11743 0.047
R12013 VDD.n10800 VDD.n10799 0.047
R12014 VDD.n10796 VDD.n10795 0.047
R12015 VDD.n10792 VDD.n10791 0.047
R12016 VDD.n10967 VDD.n10966 0.047
R12017 VDD.n10971 VDD.n10970 0.047
R12018 VDD.n10975 VDD.n10974 0.047
R12019 VDD.n10944 VDD.n10943 0.047
R12020 VDD.n11024 VDD.n11023 0.047
R12021 VDD.n11039 VDD.n11038 0.047
R12022 VDD.n11056 VDD.n11055 0.047
R12023 VDD.n10854 VDD.n10853 0.047
R12024 VDD.n10843 VDD.n10842 0.047
R12025 VDD.n10827 VDD.n10826 0.047
R12026 VDD.n10821 VDD.n10820 0.047
R12027 VDD.n10731 VDD.n10730 0.047
R12028 VDD.n10747 VDD.n10746 0.047
R12029 VDD.n11701 VDD.n11700 0.047
R12030 VDD.n11791 VDD.n11790 0.047
R12031 VDD.n11806 VDD.n11805 0.047
R12032 VDD.n11822 VDD.n11821 0.047
R12033 VDD.n11635 VDD.n11634 0.047
R12034 VDD.n11622 VDD.n11621 0.047
R12035 VDD.n11607 VDD.n11606 0.047
R12036 VDD.n11590 VDD.n11589 0.047
R12037 VDD.n11502 VDD.n11501 0.047
R12038 VDD.n11518 VDD.n11517 0.047
R12039 VDD.n11927 VDD.n11926 0.047
R12040 VDD.n4604 VDD.n4603 0.045
R12041 VDD.n2939 VDD.n2938 0.045
R12042 VDD.n1998 VDD.n1997 0.045
R12043 VDD.n5490 VDD.n5489 0.045
R12044 VDD.n5514 VDD.n5513 0.045
R12045 VDD.n5851 VDD.n5850 0.045
R12046 VDD.n5875 VDD.n5874 0.045
R12047 VDD.n6213 VDD.n6212 0.045
R12048 VDD.n6237 VDD.n6236 0.045
R12049 VDD.n6575 VDD.n6574 0.045
R12050 VDD.n6599 VDD.n6598 0.045
R12051 VDD.n6937 VDD.n6936 0.045
R12052 VDD.n6961 VDD.n6960 0.045
R12053 VDD.n7299 VDD.n7298 0.045
R12054 VDD.n7323 VDD.n7322 0.045
R12055 VDD.n7661 VDD.n7660 0.045
R12056 VDD.n7685 VDD.n7684 0.045
R12057 VDD.n8023 VDD.n8022 0.045
R12058 VDD.n8047 VDD.n8046 0.045
R12059 VDD.n8385 VDD.n8384 0.045
R12060 VDD.n8409 VDD.n8408 0.045
R12061 VDD.n8747 VDD.n8746 0.045
R12062 VDD.n8771 VDD.n8770 0.045
R12063 VDD.n9109 VDD.n9108 0.045
R12064 VDD.n9133 VDD.n9132 0.045
R12065 VDD.n9471 VDD.n9470 0.045
R12066 VDD.n9495 VDD.n9494 0.045
R12067 VDD.n9833 VDD.n9832 0.045
R12068 VDD.n9857 VDD.n9856 0.045
R12069 VDD.n10763 VDD.n10762 0.045
R12070 VDD.n11533 VDD.n11532 0.045
R12071 VDD.n10782 VDD.n10724 0.044
R12072 VDD.n11552 VDD.n11494 0.044
R12073 VDD.n4586 VDD.n4585 0.044
R12074 VDD.n2880 VDD.n2873 0.044
R12075 VDD.n295 VDD.n287 0.044
R12076 VDD.n1980 VDD.n1979 0.044
R12077 VDD.n10957 VDD.n10909 0.044
R12078 VDD.n11726 VDD.n11677 0.044
R12079 VDD.n11855 VDD.n11782 0.044
R12080 VDD.n11088 VDD.n11014 0.043
R12081 VDD.n4609 VDD.n4608 0.043
R12082 VDD.n2944 VDD.n2943 0.043
R12083 VDD.n361 VDD.n360 0.043
R12084 VDD.n2003 VDD.n2002 0.043
R12085 VDD.n5500 VDD.n5499 0.043
R12086 VDD.n5621 VDD.n5617 0.043
R12087 VDD.n5403 VDD.n5402 0.043
R12088 VDD.n5421 VDD.n5420 0.043
R12089 VDD.n5861 VDD.n5860 0.043
R12090 VDD.n5982 VDD.n5978 0.043
R12091 VDD.n5764 VDD.n5763 0.043
R12092 VDD.n5782 VDD.n5781 0.043
R12093 VDD.n6223 VDD.n6222 0.043
R12094 VDD.n6344 VDD.n6340 0.043
R12095 VDD.n6126 VDD.n6125 0.043
R12096 VDD.n6144 VDD.n6143 0.043
R12097 VDD.n6585 VDD.n6584 0.043
R12098 VDD.n6706 VDD.n6702 0.043
R12099 VDD.n6488 VDD.n6487 0.043
R12100 VDD.n6506 VDD.n6505 0.043
R12101 VDD.n6947 VDD.n6946 0.043
R12102 VDD.n7068 VDD.n7064 0.043
R12103 VDD.n6850 VDD.n6849 0.043
R12104 VDD.n6868 VDD.n6867 0.043
R12105 VDD.n7309 VDD.n7308 0.043
R12106 VDD.n7430 VDD.n7426 0.043
R12107 VDD.n7212 VDD.n7211 0.043
R12108 VDD.n7230 VDD.n7229 0.043
R12109 VDD.n7671 VDD.n7670 0.043
R12110 VDD.n7792 VDD.n7788 0.043
R12111 VDD.n7574 VDD.n7573 0.043
R12112 VDD.n7592 VDD.n7591 0.043
R12113 VDD.n8033 VDD.n8032 0.043
R12114 VDD.n8154 VDD.n8150 0.043
R12115 VDD.n7936 VDD.n7935 0.043
R12116 VDD.n7954 VDD.n7953 0.043
R12117 VDD.n8395 VDD.n8394 0.043
R12118 VDD.n8516 VDD.n8512 0.043
R12119 VDD.n8298 VDD.n8297 0.043
R12120 VDD.n8316 VDD.n8315 0.043
R12121 VDD.n8757 VDD.n8756 0.043
R12122 VDD.n8878 VDD.n8874 0.043
R12123 VDD.n8660 VDD.n8659 0.043
R12124 VDD.n8678 VDD.n8677 0.043
R12125 VDD.n9119 VDD.n9118 0.043
R12126 VDD.n9240 VDD.n9236 0.043
R12127 VDD.n9022 VDD.n9021 0.043
R12128 VDD.n9040 VDD.n9039 0.043
R12129 VDD.n9481 VDD.n9480 0.043
R12130 VDD.n9602 VDD.n9598 0.043
R12131 VDD.n9384 VDD.n9383 0.043
R12132 VDD.n9402 VDD.n9401 0.043
R12133 VDD.n9843 VDD.n9842 0.043
R12134 VDD.n9964 VDD.n9960 0.043
R12135 VDD.n9746 VDD.n9745 0.043
R12136 VDD.n9764 VDD.n9763 0.043
R12137 VDD.n11645 VDD.n11644 0.043
R12138 VDD.n11644 VDD.n11578 0.043
R12139 VDD.n10874 VDD.n10873 0.043
R12140 VDD.n10873 VDD.n10808 0.043
R12141 VDD.n10950 VDD.n10949 0.043
R12142 VDD.n11716 VDD.n11715 0.043
R12143 VDD.n11643 VDD.n11579 0.043
R12144 VDD.n5382 VDD.n5380 0.043
R12145 VDD.n5743 VDD.n5741 0.043
R12146 VDD.n6105 VDD.n6103 0.043
R12147 VDD.n6467 VDD.n6465 0.043
R12148 VDD.n6829 VDD.n6827 0.043
R12149 VDD.n7191 VDD.n7189 0.043
R12150 VDD.n7553 VDD.n7551 0.043
R12151 VDD.n7915 VDD.n7913 0.043
R12152 VDD.n8277 VDD.n8275 0.043
R12153 VDD.n8639 VDD.n8637 0.043
R12154 VDD.n9001 VDD.n8999 0.043
R12155 VDD.n9363 VDD.n9361 0.043
R12156 VDD.n9725 VDD.n9723 0.043
R12157 VDD.n11855 VDD.n11854 0.043
R12158 VDD.n4585 VDD.n4584 0.042
R12159 VDD.n2873 VDD.n2872 0.042
R12160 VDD.n287 VDD.n286 0.042
R12161 VDD.n1979 VDD.n1978 0.042
R12162 VDD.n11880 VDD.n11879 0.042
R12163 VDD.n11088 VDD.n11087 0.042
R12164 VDD.n10957 VDD.n10956 0.041
R12165 VDD.n11726 VDD.n11725 0.041
R12166 VDD.n1 VDD.n0 0.041
R12167 VDD.n5103 VDD.n5102 0.041
R12168 VDD.n5353 VDD.n5352 0.041
R12169 VDD.n5346 VDD.n5345 0.041
R12170 VDD.n5504 VDD.n5503 0.041
R12171 VDD.n5604 VDD.n5603 0.041
R12172 VDD.n5653 VDD.n5652 0.041
R12173 VDD.n5411 VDD.n5410 0.041
R12174 VDD.n5459 VDD.n5455 0.041
R12175 VDD.n5714 VDD.n5713 0.041
R12176 VDD.n5707 VDD.n5706 0.041
R12177 VDD.n5865 VDD.n5864 0.041
R12178 VDD.n5965 VDD.n5964 0.041
R12179 VDD.n6014 VDD.n6013 0.041
R12180 VDD.n5772 VDD.n5771 0.041
R12181 VDD.n5820 VDD.n5816 0.041
R12182 VDD.n6076 VDD.n6075 0.041
R12183 VDD.n6069 VDD.n6068 0.041
R12184 VDD.n6227 VDD.n6226 0.041
R12185 VDD.n6327 VDD.n6326 0.041
R12186 VDD.n6376 VDD.n6375 0.041
R12187 VDD.n6134 VDD.n6133 0.041
R12188 VDD.n6182 VDD.n6178 0.041
R12189 VDD.n6438 VDD.n6437 0.041
R12190 VDD.n6431 VDD.n6430 0.041
R12191 VDD.n6589 VDD.n6588 0.041
R12192 VDD.n6689 VDD.n6688 0.041
R12193 VDD.n6738 VDD.n6737 0.041
R12194 VDD.n6496 VDD.n6495 0.041
R12195 VDD.n6544 VDD.n6540 0.041
R12196 VDD.n6800 VDD.n6799 0.041
R12197 VDD.n6793 VDD.n6792 0.041
R12198 VDD.n6951 VDD.n6950 0.041
R12199 VDD.n7051 VDD.n7050 0.041
R12200 VDD.n7100 VDD.n7099 0.041
R12201 VDD.n6858 VDD.n6857 0.041
R12202 VDD.n6906 VDD.n6902 0.041
R12203 VDD.n7162 VDD.n7161 0.041
R12204 VDD.n7155 VDD.n7154 0.041
R12205 VDD.n7313 VDD.n7312 0.041
R12206 VDD.n7413 VDD.n7412 0.041
R12207 VDD.n7462 VDD.n7461 0.041
R12208 VDD.n7220 VDD.n7219 0.041
R12209 VDD.n7268 VDD.n7264 0.041
R12210 VDD.n7524 VDD.n7523 0.041
R12211 VDD.n7517 VDD.n7516 0.041
R12212 VDD.n7675 VDD.n7674 0.041
R12213 VDD.n7775 VDD.n7774 0.041
R12214 VDD.n7824 VDD.n7823 0.041
R12215 VDD.n7582 VDD.n7581 0.041
R12216 VDD.n7630 VDD.n7626 0.041
R12217 VDD.n7886 VDD.n7885 0.041
R12218 VDD.n7879 VDD.n7878 0.041
R12219 VDD.n8037 VDD.n8036 0.041
R12220 VDD.n8137 VDD.n8136 0.041
R12221 VDD.n8186 VDD.n8185 0.041
R12222 VDD.n7944 VDD.n7943 0.041
R12223 VDD.n7992 VDD.n7988 0.041
R12224 VDD.n8248 VDD.n8247 0.041
R12225 VDD.n8241 VDD.n8240 0.041
R12226 VDD.n8399 VDD.n8398 0.041
R12227 VDD.n8499 VDD.n8498 0.041
R12228 VDD.n8548 VDD.n8547 0.041
R12229 VDD.n8306 VDD.n8305 0.041
R12230 VDD.n8354 VDD.n8350 0.041
R12231 VDD.n8610 VDD.n8609 0.041
R12232 VDD.n8603 VDD.n8602 0.041
R12233 VDD.n8761 VDD.n8760 0.041
R12234 VDD.n8861 VDD.n8860 0.041
R12235 VDD.n8910 VDD.n8909 0.041
R12236 VDD.n8668 VDD.n8667 0.041
R12237 VDD.n8716 VDD.n8712 0.041
R12238 VDD.n8972 VDD.n8971 0.041
R12239 VDD.n8965 VDD.n8964 0.041
R12240 VDD.n9123 VDD.n9122 0.041
R12241 VDD.n9223 VDD.n9222 0.041
R12242 VDD.n9272 VDD.n9271 0.041
R12243 VDD.n9030 VDD.n9029 0.041
R12244 VDD.n9078 VDD.n9074 0.041
R12245 VDD.n9334 VDD.n9333 0.041
R12246 VDD.n9327 VDD.n9326 0.041
R12247 VDD.n9485 VDD.n9484 0.041
R12248 VDD.n9585 VDD.n9584 0.041
R12249 VDD.n9634 VDD.n9633 0.041
R12250 VDD.n9392 VDD.n9391 0.041
R12251 VDD.n9440 VDD.n9436 0.041
R12252 VDD.n9696 VDD.n9695 0.041
R12253 VDD.n9689 VDD.n9688 0.041
R12254 VDD.n9847 VDD.n9846 0.041
R12255 VDD.n9947 VDD.n9946 0.041
R12256 VDD.n9996 VDD.n9995 0.041
R12257 VDD.n9754 VDD.n9753 0.041
R12258 VDD.n9802 VDD.n9798 0.041
R12259 VDD.n11101 VDD.n11100 0.041
R12260 VDD.n12232 VDD.n12231 0.041
R12261 VDD.n5666 VDD.n5663 0.041
R12262 VDD.n6027 VDD.n6024 0.041
R12263 VDD.n6389 VDD.n6386 0.041
R12264 VDD.n6751 VDD.n6748 0.041
R12265 VDD.n7113 VDD.n7110 0.041
R12266 VDD.n7475 VDD.n7472 0.041
R12267 VDD.n7837 VDD.n7834 0.041
R12268 VDD.n8199 VDD.n8196 0.041
R12269 VDD.n8561 VDD.n8558 0.041
R12270 VDD.n8923 VDD.n8920 0.041
R12271 VDD.n9285 VDD.n9282 0.041
R12272 VDD.n9647 VDD.n9644 0.041
R12273 VDD.n10009 VDD.n10006 0.041
R12274 VDD.n10782 VDD.n10781 0.041
R12275 VDD.n11552 VDD.n11551 0.041
R12276 VDD.n11 VDD.n7 0.04
R12277 VDD.n2808 VDD.n2794 0.04
R12278 VDD.n3129 VDD.n3118 0.04
R12279 VDD.n3367 VDD.n3356 0.04
R12280 VDD.n3604 VDD.n3593 0.04
R12281 VDD.n3842 VDD.n3831 0.04
R12282 VDD.n4079 VDD.n4068 0.04
R12283 VDD.n4317 VDD.n4306 0.04
R12284 VDD.n12242 VDD.n12238 0.04
R12285 VDD.n2499 VDD.n2498 0.039
R12286 VDD.n5137 VDD.n5136 0.039
R12287 VDD.n5372 VDD.n5371 0.039
R12288 VDD.n5469 VDD.n5466 0.039
R12289 VDD.n5602 VDD.n5601 0.039
R12290 VDD.n5630 VDD.n5629 0.039
R12291 VDD.n5563 VDD.n5561 0.039
R12292 VDD.n5733 VDD.n5732 0.039
R12293 VDD.n5830 VDD.n5827 0.039
R12294 VDD.n5963 VDD.n5962 0.039
R12295 VDD.n5991 VDD.n5990 0.039
R12296 VDD.n5924 VDD.n5922 0.039
R12297 VDD.n6095 VDD.n6094 0.039
R12298 VDD.n6192 VDD.n6189 0.039
R12299 VDD.n6325 VDD.n6324 0.039
R12300 VDD.n6353 VDD.n6352 0.039
R12301 VDD.n6286 VDD.n6284 0.039
R12302 VDD.n6457 VDD.n6456 0.039
R12303 VDD.n6554 VDD.n6551 0.039
R12304 VDD.n6687 VDD.n6686 0.039
R12305 VDD.n6715 VDD.n6714 0.039
R12306 VDD.n6648 VDD.n6646 0.039
R12307 VDD.n6819 VDD.n6818 0.039
R12308 VDD.n6916 VDD.n6913 0.039
R12309 VDD.n7049 VDD.n7048 0.039
R12310 VDD.n7077 VDD.n7076 0.039
R12311 VDD.n7010 VDD.n7008 0.039
R12312 VDD.n7181 VDD.n7180 0.039
R12313 VDD.n7278 VDD.n7275 0.039
R12314 VDD.n7411 VDD.n7410 0.039
R12315 VDD.n7439 VDD.n7438 0.039
R12316 VDD.n7372 VDD.n7370 0.039
R12317 VDD.n7543 VDD.n7542 0.039
R12318 VDD.n7640 VDD.n7637 0.039
R12319 VDD.n7773 VDD.n7772 0.039
R12320 VDD.n7801 VDD.n7800 0.039
R12321 VDD.n7734 VDD.n7732 0.039
R12322 VDD.n7905 VDD.n7904 0.039
R12323 VDD.n8002 VDD.n7999 0.039
R12324 VDD.n8135 VDD.n8134 0.039
R12325 VDD.n8163 VDD.n8162 0.039
R12326 VDD.n8096 VDD.n8094 0.039
R12327 VDD.n8267 VDD.n8266 0.039
R12328 VDD.n8364 VDD.n8361 0.039
R12329 VDD.n8497 VDD.n8496 0.039
R12330 VDD.n8525 VDD.n8524 0.039
R12331 VDD.n8458 VDD.n8456 0.039
R12332 VDD.n8629 VDD.n8628 0.039
R12333 VDD.n8726 VDD.n8723 0.039
R12334 VDD.n8859 VDD.n8858 0.039
R12335 VDD.n8887 VDD.n8886 0.039
R12336 VDD.n8820 VDD.n8818 0.039
R12337 VDD.n8991 VDD.n8990 0.039
R12338 VDD.n9088 VDD.n9085 0.039
R12339 VDD.n9221 VDD.n9220 0.039
R12340 VDD.n9249 VDD.n9248 0.039
R12341 VDD.n9182 VDD.n9180 0.039
R12342 VDD.n9353 VDD.n9352 0.039
R12343 VDD.n9450 VDD.n9447 0.039
R12344 VDD.n9583 VDD.n9582 0.039
R12345 VDD.n9611 VDD.n9610 0.039
R12346 VDD.n9544 VDD.n9542 0.039
R12347 VDD.n9715 VDD.n9714 0.039
R12348 VDD.n9812 VDD.n9809 0.039
R12349 VDD.n9945 VDD.n9944 0.039
R12350 VDD.n9973 VDD.n9972 0.039
R12351 VDD.n9906 VDD.n9904 0.039
R12352 VDD.n5013 VDD.n5002 0.038
R12353 VDD.n4994 VDD.n4992 0.038
R12354 VDD.n4782 VDD.n4771 0.038
R12355 VDD.n4763 VDD.n4761 0.038
R12356 VDD.n2992 VDD.n2991 0.038
R12357 VDD.n3016 VDD.n3015 0.038
R12358 VDD.n3230 VDD.n3229 0.038
R12359 VDD.n3253 VDD.n3252 0.038
R12360 VDD.n3467 VDD.n3466 0.038
R12361 VDD.n3491 VDD.n3490 0.038
R12362 VDD.n3705 VDD.n3704 0.038
R12363 VDD.n3728 VDD.n3727 0.038
R12364 VDD.n3942 VDD.n3941 0.038
R12365 VDD.n3966 VDD.n3965 0.038
R12366 VDD.n4180 VDD.n4179 0.038
R12367 VDD.n4203 VDD.n4202 0.038
R12368 VDD.n4417 VDD.n4416 0.038
R12369 VDD.n4441 VDD.n4440 0.038
R12370 VDD.n409 VDD.n408 0.038
R12371 VDD.n436 VDD.n435 0.038
R12372 VDD.n643 VDD.n642 0.038
R12373 VDD.n669 VDD.n668 0.038
R12374 VDD.n876 VDD.n875 0.038
R12375 VDD.n903 VDD.n902 0.038
R12376 VDD.n1110 VDD.n1109 0.038
R12377 VDD.n1136 VDD.n1135 0.038
R12378 VDD.n1343 VDD.n1342 0.038
R12379 VDD.n1370 VDD.n1369 0.038
R12380 VDD.n1577 VDD.n1576 0.038
R12381 VDD.n1603 VDD.n1602 0.038
R12382 VDD.n1810 VDD.n1809 0.038
R12383 VDD.n1837 VDD.n1836 0.038
R12384 VDD.n2159 VDD.n2157 0.038
R12385 VDD.n2178 VDD.n2167 0.038
R12386 VDD.n2390 VDD.n2388 0.038
R12387 VDD.n2409 VDD.n2398 0.038
R12388 VDD.n185 VDD.n184 0.037
R12389 VDD.n2698 VDD.n2697 0.037
R12390 VDD.n5344 VDD.n5343 0.037
R12391 VDD.n5705 VDD.n5704 0.037
R12392 VDD.n6067 VDD.n6066 0.037
R12393 VDD.n6429 VDD.n6428 0.037
R12394 VDD.n6791 VDD.n6790 0.037
R12395 VDD.n7153 VDD.n7152 0.037
R12396 VDD.n7515 VDD.n7514 0.037
R12397 VDD.n7877 VDD.n7876 0.037
R12398 VDD.n8239 VDD.n8238 0.037
R12399 VDD.n8601 VDD.n8600 0.037
R12400 VDD.n8963 VDD.n8962 0.037
R12401 VDD.n9325 VDD.n9324 0.037
R12402 VDD.n9687 VDD.n9686 0.037
R12403 VDD.n11567 VDD.n11566 0.037
R12404 VDD.n11563 VDD.n11562 0.037
R12405 VDD.n11739 VDD.n11738 0.037
R12406 VDD.n11743 VDD.n11742 0.037
R12407 VDD.n10797 VDD.n10796 0.037
R12408 VDD.n10793 VDD.n10792 0.037
R12409 VDD.n10970 VDD.n10969 0.037
R12410 VDD.n10974 VDD.n10973 0.037
R12411 VDD.n11023 VDD.n11022 0.037
R12412 VDD.n10822 VDD.n10821 0.037
R12413 VDD.n10730 VDD.n10729 0.037
R12414 VDD.n11790 VDD.n11789 0.037
R12415 VDD.n11591 VDD.n11590 0.037
R12416 VDD.n11501 VDD.n11500 0.037
R12417 VDD.n4898 VDD.n4896 0.036
R12418 VDD.n4870 VDD.n4868 0.036
R12419 VDD.n4667 VDD.n4665 0.036
R12420 VDD.n4639 VDD.n4637 0.036
R12421 VDD.n4601 VDD.n4600 0.036
R12422 VDD.n4581 VDD.n4580 0.036
R12423 VDD.n2815 VDD.n2814 0.036
R12424 VDD.n2849 VDD.n2847 0.036
R12425 VDD.n2788 VDD.n2787 0.036
R12426 VDD.n2840 VDD.n2810 0.036
R12427 VDD.n3113 VDD.n3112 0.036
R12428 VDD.n3143 VDD.n3131 0.036
R12429 VDD.n3351 VDD.n3350 0.036
R12430 VDD.n3381 VDD.n3369 0.036
R12431 VDD.n3588 VDD.n3587 0.036
R12432 VDD.n3618 VDD.n3606 0.036
R12433 VDD.n3826 VDD.n3825 0.036
R12434 VDD.n3856 VDD.n3844 0.036
R12435 VDD.n4063 VDD.n4062 0.036
R12436 VDD.n4093 VDD.n4081 0.036
R12437 VDD.n4301 VDD.n4300 0.036
R12438 VDD.n4331 VDD.n4319 0.036
R12439 VDD.n4624 VDD.n4623 0.036
R12440 VDD.n2807 VDD.n2800 0.036
R12441 VDD.n2797 VDD.n2796 0.036
R12442 VDD.n2796 VDD.n2795 0.036
R12443 VDD.n2839 VDD.n2825 0.036
R12444 VDD.n2827 VDD.n2826 0.036
R12445 VDD.n2883 VDD.n2882 0.036
R12446 VDD.n2914 VDD.n2901 0.036
R12447 VDD.n2903 VDD.n2902 0.036
R12448 VDD.n2954 VDD.n2953 0.036
R12449 VDD.n4461 VDD.n4460 0.036
R12450 VDD.n4464 VDD.n4463 0.036
R12451 VDD.n4537 VDD.n4536 0.036
R12452 VDD.n4564 VDD.n4563 0.036
R12453 VDD.n239 VDD.n238 0.036
R12454 VDD.n264 VDD.n263 0.036
R12455 VDD.n1995 VDD.n1994 0.036
R12456 VDD.n1975 VDD.n1974 0.036
R12457 VDD.n216 VDD.n215 0.036
R12458 VDD.n256 VDD.n227 0.036
R12459 VDD.n533 VDD.n532 0.036
R12460 VDD.n556 VDD.n544 0.036
R12461 VDD.n767 VDD.n766 0.036
R12462 VDD.n790 VDD.n778 0.036
R12463 VDD.n1000 VDD.n999 0.036
R12464 VDD.n1023 VDD.n1011 0.036
R12465 VDD.n1234 VDD.n1233 0.036
R12466 VDD.n1257 VDD.n1245 0.036
R12467 VDD.n1467 VDD.n1466 0.036
R12468 VDD.n1490 VDD.n1478 0.036
R12469 VDD.n1701 VDD.n1700 0.036
R12470 VDD.n1724 VDD.n1712 0.036
R12471 VDD.n2019 VDD.n2018 0.036
R12472 VDD.n2035 VDD.n2033 0.036
R12473 VDD.n2063 VDD.n2061 0.036
R12474 VDD.n2266 VDD.n2264 0.036
R12475 VDD.n2294 VDD.n2292 0.036
R12476 VDD.n2527 VDD.n2526 0.035
R12477 VDD.n5296 VDD.n5233 0.035
R12478 VDD.n5296 VDD.n5295 0.035
R12479 VDD.n2529 VDD.n2528 0.035
R12480 VDD.n179 VDD.n178 0.035
R12481 VDD.n157 VDD.n156 0.035
R12482 VDD.n5298 VDD.n5297 0.035
R12483 VDD.n2691 VDD.n2690 0.035
R12484 VDD.n5616 VDD.n5615 0.035
R12485 VDD.n5314 VDD.n5313 0.035
R12486 VDD.n5977 VDD.n5976 0.035
R12487 VDD.n5675 VDD.n5674 0.035
R12488 VDD.n6339 VDD.n6338 0.035
R12489 VDD.n6037 VDD.n6036 0.035
R12490 VDD.n6701 VDD.n6700 0.035
R12491 VDD.n6399 VDD.n6398 0.035
R12492 VDD.n7063 VDD.n7062 0.035
R12493 VDD.n6761 VDD.n6760 0.035
R12494 VDD.n7425 VDD.n7424 0.035
R12495 VDD.n7123 VDD.n7122 0.035
R12496 VDD.n7787 VDD.n7786 0.035
R12497 VDD.n7485 VDD.n7484 0.035
R12498 VDD.n8149 VDD.n8148 0.035
R12499 VDD.n7847 VDD.n7846 0.035
R12500 VDD.n8511 VDD.n8510 0.035
R12501 VDD.n8209 VDD.n8208 0.035
R12502 VDD.n8873 VDD.n8872 0.035
R12503 VDD.n8571 VDD.n8570 0.035
R12504 VDD.n9235 VDD.n9234 0.035
R12505 VDD.n8933 VDD.n8932 0.035
R12506 VDD.n9597 VDD.n9596 0.035
R12507 VDD.n9295 VDD.n9294 0.035
R12508 VDD.n9959 VDD.n9958 0.035
R12509 VDD.n9657 VDD.n9656 0.035
R12510 VDD.n10436 VDD.n10435 0.035
R12511 VDD.n10442 VDD.n10441 0.035
R12512 VDD.n10399 VDD.n10398 0.035
R12513 VDD.n10416 VDD.n10415 0.035
R12514 VDD.n10372 VDD.n10371 0.035
R12515 VDD.n10389 VDD.n10388 0.035
R12516 VDD.n10355 VDD.n10354 0.035
R12517 VDD.n10362 VDD.n10361 0.035
R12518 VDD.n11940 VDD.n11645 0.035
R12519 VDD.n11569 VDD.n11568 0.035
R12520 VDD.n11565 VDD.n11564 0.035
R12521 VDD.n11554 VDD.n11553 0.035
R12522 VDD.n11737 VDD.n11736 0.035
R12523 VDD.n11741 VDD.n11740 0.035
R12524 VDD.n11183 VDD.n10874 0.035
R12525 VDD.n10799 VDD.n10798 0.035
R12526 VDD.n10795 VDD.n10794 0.035
R12527 VDD.n10784 VDD.n10783 0.035
R12528 VDD.n10968 VDD.n10967 0.035
R12529 VDD.n10972 VDD.n10971 0.035
R12530 VDD.n11021 VDD.n11017 0.035
R12531 VDD.n11025 VDD.n11024 0.035
R12532 VDD.n10768 VDD.n10764 0.035
R12533 VDD.n11788 VDD.n11783 0.035
R12534 VDD.n11792 VDD.n11791 0.035
R12535 VDD.n11538 VDD.n11534 0.035
R12536 VDD.n5085 VDD.n5084 0.035
R12537 VDD.n164 VDD.n158 0.034
R12538 VDD.n4590 VDD.n4589 0.034
R12539 VDD.n2877 VDD.n2876 0.034
R12540 VDD.n292 VDD.n291 0.034
R12541 VDD.n1984 VDD.n1983 0.034
R12542 VDD.n371 VDD.n370 0.034
R12543 VDD.n5273 VDD.n5272 0.034
R12544 VDD.n5125 VDD.n2764 0.034
R12545 VDD.n186 VDD.n185 0.034
R12546 VDD.n5127 VDD.n5126 0.034
R12547 VDD.n5138 VDD.n5137 0.034
R12548 VDD.n5482 VDD.n5479 0.034
R12549 VDD.n5502 VDD.n5501 0.034
R12550 VDD.n5402 VDD.n5401 0.034
R12551 VDD.n5409 VDD.n5408 0.034
R12552 VDD.n5454 VDD.n5453 0.034
R12553 VDD.n5464 VDD.n5463 0.034
R12554 VDD.n5560 VDD.n5559 0.034
R12555 VDD.n5568 VDD.n5567 0.034
R12556 VDD.n5843 VDD.n5840 0.034
R12557 VDD.n5863 VDD.n5862 0.034
R12558 VDD.n5763 VDD.n5762 0.034
R12559 VDD.n5770 VDD.n5769 0.034
R12560 VDD.n5815 VDD.n5814 0.034
R12561 VDD.n5825 VDD.n5824 0.034
R12562 VDD.n5921 VDD.n5920 0.034
R12563 VDD.n5929 VDD.n5928 0.034
R12564 VDD.n6205 VDD.n6202 0.034
R12565 VDD.n6225 VDD.n6224 0.034
R12566 VDD.n6125 VDD.n6124 0.034
R12567 VDD.n6132 VDD.n6131 0.034
R12568 VDD.n6177 VDD.n6176 0.034
R12569 VDD.n6187 VDD.n6186 0.034
R12570 VDD.n6283 VDD.n6282 0.034
R12571 VDD.n6291 VDD.n6290 0.034
R12572 VDD.n6567 VDD.n6564 0.034
R12573 VDD.n6587 VDD.n6586 0.034
R12574 VDD.n6487 VDD.n6486 0.034
R12575 VDD.n6494 VDD.n6493 0.034
R12576 VDD.n6539 VDD.n6538 0.034
R12577 VDD.n6549 VDD.n6548 0.034
R12578 VDD.n6645 VDD.n6644 0.034
R12579 VDD.n6653 VDD.n6652 0.034
R12580 VDD.n6929 VDD.n6926 0.034
R12581 VDD.n6949 VDD.n6948 0.034
R12582 VDD.n6849 VDD.n6848 0.034
R12583 VDD.n6856 VDD.n6855 0.034
R12584 VDD.n6901 VDD.n6900 0.034
R12585 VDD.n6911 VDD.n6910 0.034
R12586 VDD.n7007 VDD.n7006 0.034
R12587 VDD.n7015 VDD.n7014 0.034
R12588 VDD.n7291 VDD.n7288 0.034
R12589 VDD.n7311 VDD.n7310 0.034
R12590 VDD.n7211 VDD.n7210 0.034
R12591 VDD.n7218 VDD.n7217 0.034
R12592 VDD.n7263 VDD.n7262 0.034
R12593 VDD.n7273 VDD.n7272 0.034
R12594 VDD.n7369 VDD.n7368 0.034
R12595 VDD.n7377 VDD.n7376 0.034
R12596 VDD.n7653 VDD.n7650 0.034
R12597 VDD.n7673 VDD.n7672 0.034
R12598 VDD.n7573 VDD.n7572 0.034
R12599 VDD.n7580 VDD.n7579 0.034
R12600 VDD.n7625 VDD.n7624 0.034
R12601 VDD.n7635 VDD.n7634 0.034
R12602 VDD.n7731 VDD.n7730 0.034
R12603 VDD.n7739 VDD.n7738 0.034
R12604 VDD.n8015 VDD.n8012 0.034
R12605 VDD.n8035 VDD.n8034 0.034
R12606 VDD.n7935 VDD.n7934 0.034
R12607 VDD.n7942 VDD.n7941 0.034
R12608 VDD.n7987 VDD.n7986 0.034
R12609 VDD.n7997 VDD.n7996 0.034
R12610 VDD.n8093 VDD.n8092 0.034
R12611 VDD.n8101 VDD.n8100 0.034
R12612 VDD.n8377 VDD.n8374 0.034
R12613 VDD.n8397 VDD.n8396 0.034
R12614 VDD.n8297 VDD.n8296 0.034
R12615 VDD.n8304 VDD.n8303 0.034
R12616 VDD.n8349 VDD.n8348 0.034
R12617 VDD.n8359 VDD.n8358 0.034
R12618 VDD.n8455 VDD.n8454 0.034
R12619 VDD.n8463 VDD.n8462 0.034
R12620 VDD.n8739 VDD.n8736 0.034
R12621 VDD.n8759 VDD.n8758 0.034
R12622 VDD.n8659 VDD.n8658 0.034
R12623 VDD.n8666 VDD.n8665 0.034
R12624 VDD.n8711 VDD.n8710 0.034
R12625 VDD.n8721 VDD.n8720 0.034
R12626 VDD.n8817 VDD.n8816 0.034
R12627 VDD.n8825 VDD.n8824 0.034
R12628 VDD.n9101 VDD.n9098 0.034
R12629 VDD.n9121 VDD.n9120 0.034
R12630 VDD.n9021 VDD.n9020 0.034
R12631 VDD.n9028 VDD.n9027 0.034
R12632 VDD.n9073 VDD.n9072 0.034
R12633 VDD.n9083 VDD.n9082 0.034
R12634 VDD.n9179 VDD.n9178 0.034
R12635 VDD.n9187 VDD.n9186 0.034
R12636 VDD.n9463 VDD.n9460 0.034
R12637 VDD.n9483 VDD.n9482 0.034
R12638 VDD.n9383 VDD.n9382 0.034
R12639 VDD.n9390 VDD.n9389 0.034
R12640 VDD.n9435 VDD.n9434 0.034
R12641 VDD.n9445 VDD.n9444 0.034
R12642 VDD.n9541 VDD.n9540 0.034
R12643 VDD.n9549 VDD.n9548 0.034
R12644 VDD.n9825 VDD.n9822 0.034
R12645 VDD.n9845 VDD.n9844 0.034
R12646 VDD.n9745 VDD.n9744 0.034
R12647 VDD.n9752 VDD.n9751 0.034
R12648 VDD.n9797 VDD.n9796 0.034
R12649 VDD.n9807 VDD.n9806 0.034
R12650 VDD.n9903 VDD.n9902 0.034
R12651 VDD.n9911 VDD.n9910 0.034
R12652 VDD.n10301 VDD.n10299 0.034
R12653 VDD.n10276 VDD.n10274 0.034
R12654 VDD.n10183 VDD.n10181 0.034
R12655 VDD.n10159 VDD.n10157 0.034
R12656 VDD.n10101 VDD.n10099 0.034
R12657 VDD.n10076 VDD.n10074 0.034
R12658 VDD.n10056 VDD.n10054 0.034
R12659 VDD.n10031 VDD.n10029 0.034
R12660 VDD.n10648 VDD.n10646 0.034
R12661 VDD.n10623 VDD.n10621 0.034
R12662 VDD.n10529 VDD.n10527 0.034
R12663 VDD.n10505 VDD.n10503 0.034
R12664 VDD.n11578 VDD.n11577 0.034
R12665 VDD.n11728 VDD.n11727 0.034
R12666 VDD.n10808 VDD.n10807 0.034
R12667 VDD.n10959 VDD.n10958 0.034
R12668 VDD.n10952 VDD.n10951 0.034
R12669 VDD.n10858 VDD.n10855 0.034
R12670 VDD.n11721 VDD.n11717 0.034
R12671 VDD.n11639 VDD.n11636 0.034
R12672 VDD.n2481 VDD.n2480 0.034
R12673 VDD.n5027 VDD.n5017 0.033
R12674 VDD.n4980 VDD.n4978 0.033
R12675 VDD.n4796 VDD.n4786 0.033
R12676 VDD.n4749 VDD.n4747 0.033
R12677 VDD.n4612 VDD.n4611 0.033
R12678 VDD.n2947 VDD.n2946 0.033
R12679 VDD.n2978 VDD.n2977 0.033
R12680 VDD.n3030 VDD.n3029 0.033
R12681 VDD.n3216 VDD.n3215 0.033
R12682 VDD.n3267 VDD.n3266 0.033
R12683 VDD.n3453 VDD.n3452 0.033
R12684 VDD.n3505 VDD.n3504 0.033
R12685 VDD.n3691 VDD.n3690 0.033
R12686 VDD.n3742 VDD.n3741 0.033
R12687 VDD.n3928 VDD.n3927 0.033
R12688 VDD.n3980 VDD.n3979 0.033
R12689 VDD.n4166 VDD.n4165 0.033
R12690 VDD.n4217 VDD.n4216 0.033
R12691 VDD.n4403 VDD.n4402 0.033
R12692 VDD.n4455 VDD.n4454 0.033
R12693 VDD.n364 VDD.n363 0.033
R12694 VDD.n2006 VDD.n2005 0.033
R12695 VDD.n395 VDD.n394 0.033
R12696 VDD.n450 VDD.n449 0.033
R12697 VDD.n629 VDD.n628 0.033
R12698 VDD.n683 VDD.n682 0.033
R12699 VDD.n862 VDD.n861 0.033
R12700 VDD.n917 VDD.n916 0.033
R12701 VDD.n1096 VDD.n1095 0.033
R12702 VDD.n1150 VDD.n1149 0.033
R12703 VDD.n1329 VDD.n1328 0.033
R12704 VDD.n1384 VDD.n1383 0.033
R12705 VDD.n1563 VDD.n1562 0.033
R12706 VDD.n1617 VDD.n1616 0.033
R12707 VDD.n1796 VDD.n1795 0.033
R12708 VDD.n1851 VDD.n1850 0.033
R12709 VDD.n2145 VDD.n2143 0.033
R12710 VDD.n2192 VDD.n2182 0.033
R12711 VDD.n2376 VDD.n2374 0.033
R12712 VDD.n2423 VDD.n2413 0.033
R12713 VDD.n1857 VDD.n1856 0.032
R12714 VDD.n1889 VDD.n1888 0.032
R12715 VDD.n1908 VDD.n1907 0.032
R12716 VDD.n1928 VDD.n1927 0.032
R12717 VDD.n1960 VDD.n1959 0.032
R12718 VDD.n1961 VDD.n1960 0.032
R12719 VDD.n2017 VDD.n2010 0.032
R12720 VDD.n5208 VDD.n5207 0.032
R12721 VDD.n2607 VDD.n2606 0.032
R12722 VDD.n5378 VDD.n5377 0.032
R12723 VDD.n5525 VDD.n5522 0.032
R12724 VDD.n5661 VDD.n5660 0.032
R12725 VDD.n5446 VDD.n5445 0.032
R12726 VDD.n5739 VDD.n5738 0.032
R12727 VDD.n5886 VDD.n5883 0.032
R12728 VDD.n6022 VDD.n6021 0.032
R12729 VDD.n5807 VDD.n5806 0.032
R12730 VDD.n6101 VDD.n6100 0.032
R12731 VDD.n6248 VDD.n6245 0.032
R12732 VDD.n6384 VDD.n6383 0.032
R12733 VDD.n6169 VDD.n6168 0.032
R12734 VDD.n6463 VDD.n6462 0.032
R12735 VDD.n6610 VDD.n6607 0.032
R12736 VDD.n6746 VDD.n6745 0.032
R12737 VDD.n6531 VDD.n6530 0.032
R12738 VDD.n6825 VDD.n6824 0.032
R12739 VDD.n6972 VDD.n6969 0.032
R12740 VDD.n7108 VDD.n7107 0.032
R12741 VDD.n6893 VDD.n6892 0.032
R12742 VDD.n7187 VDD.n7186 0.032
R12743 VDD.n7334 VDD.n7331 0.032
R12744 VDD.n7470 VDD.n7469 0.032
R12745 VDD.n7255 VDD.n7254 0.032
R12746 VDD.n7549 VDD.n7548 0.032
R12747 VDD.n7696 VDD.n7693 0.032
R12748 VDD.n7832 VDD.n7831 0.032
R12749 VDD.n7617 VDD.n7616 0.032
R12750 VDD.n7911 VDD.n7910 0.032
R12751 VDD.n8058 VDD.n8055 0.032
R12752 VDD.n8194 VDD.n8193 0.032
R12753 VDD.n7979 VDD.n7978 0.032
R12754 VDD.n8273 VDD.n8272 0.032
R12755 VDD.n8420 VDD.n8417 0.032
R12756 VDD.n8556 VDD.n8555 0.032
R12757 VDD.n8341 VDD.n8340 0.032
R12758 VDD.n8635 VDD.n8634 0.032
R12759 VDD.n8782 VDD.n8779 0.032
R12760 VDD.n8918 VDD.n8917 0.032
R12761 VDD.n8703 VDD.n8702 0.032
R12762 VDD.n8997 VDD.n8996 0.032
R12763 VDD.n9144 VDD.n9141 0.032
R12764 VDD.n9280 VDD.n9279 0.032
R12765 VDD.n9065 VDD.n9064 0.032
R12766 VDD.n9359 VDD.n9358 0.032
R12767 VDD.n9506 VDD.n9503 0.032
R12768 VDD.n9642 VDD.n9641 0.032
R12769 VDD.n9427 VDD.n9426 0.032
R12770 VDD.n9721 VDD.n9720 0.032
R12771 VDD.n9868 VDD.n9865 0.032
R12772 VDD.n10004 VDD.n10003 0.032
R12773 VDD.n9789 VDD.n9788 0.032
R12774 VDD.n10943 VDD.n10935 0.032
R12775 VDD.n11134 VDD.n11118 0.032
R12776 VDD.n10853 VDD.n10845 0.032
R12777 VDD.n11700 VDD.n11690 0.032
R12778 VDD.n11883 VDD.n11882 0.032
R12779 VDD.n11634 VDD.n11626 0.032
R12780 VDD.n102 VDD.n101 0.031
R12781 VDD.n4912 VDD.n4910 0.031
R12782 VDD.n4856 VDD.n4854 0.031
R12783 VDD.n4681 VDD.n4679 0.031
R12784 VDD.n2866 VDD.n2842 0.031
R12785 VDD.n3099 VDD.n3098 0.031
R12786 VDD.n3158 VDD.n3145 0.031
R12787 VDD.n3337 VDD.n3336 0.031
R12788 VDD.n3395 VDD.n3383 0.031
R12789 VDD.n3574 VDD.n3573 0.031
R12790 VDD.n3633 VDD.n3620 0.031
R12791 VDD.n3812 VDD.n3811 0.031
R12792 VDD.n3870 VDD.n3858 0.031
R12793 VDD.n4049 VDD.n4048 0.031
R12794 VDD.n4108 VDD.n4095 0.031
R12795 VDD.n4287 VDD.n4286 0.031
R12796 VDD.n4345 VDD.n4333 0.031
R12797 VDD.n4561 VDD.n4560 0.031
R12798 VDD.n279 VDD.n258 0.031
R12799 VDD.n519 VDD.n518 0.031
R12800 VDD.n571 VDD.n558 0.031
R12801 VDD.n753 VDD.n752 0.031
R12802 VDD.n804 VDD.n792 0.031
R12803 VDD.n986 VDD.n985 0.031
R12804 VDD.n1038 VDD.n1025 0.031
R12805 VDD.n1220 VDD.n1219 0.031
R12806 VDD.n1271 VDD.n1259 0.031
R12807 VDD.n1453 VDD.n1452 0.031
R12808 VDD.n1505 VDD.n1492 0.031
R12809 VDD.n1687 VDD.n1686 0.031
R12810 VDD.n1738 VDD.n1726 0.031
R12811 VDD.n1946 VDD.n1945 0.031
R12812 VDD.n2077 VDD.n2075 0.031
R12813 VDD.n2252 VDD.n2250 0.031
R12814 VDD.n2308 VDD.n2306 0.031
R12815 VDD.n5385 VDD.n5384 0.031
R12816 VDD.n5399 VDD.n5398 0.031
R12817 VDD.n5423 VDD.n5417 0.031
R12818 VDD.n5442 VDD.n5441 0.031
R12819 VDD.n5530 VDD.n5462 0.031
R12820 VDD.n5549 VDD.n5548 0.031
R12821 VDD.n5572 VDD.n5566 0.031
R12822 VDD.n5592 VDD.n5591 0.031
R12823 VDD.n5746 VDD.n5745 0.031
R12824 VDD.n5760 VDD.n5759 0.031
R12825 VDD.n5784 VDD.n5778 0.031
R12826 VDD.n5803 VDD.n5802 0.031
R12827 VDD.n5891 VDD.n5823 0.031
R12828 VDD.n5910 VDD.n5909 0.031
R12829 VDD.n5933 VDD.n5927 0.031
R12830 VDD.n5953 VDD.n5952 0.031
R12831 VDD.n6108 VDD.n6107 0.031
R12832 VDD.n6122 VDD.n6121 0.031
R12833 VDD.n6146 VDD.n6140 0.031
R12834 VDD.n6165 VDD.n6164 0.031
R12835 VDD.n6253 VDD.n6185 0.031
R12836 VDD.n6272 VDD.n6271 0.031
R12837 VDD.n6295 VDD.n6289 0.031
R12838 VDD.n6315 VDD.n6314 0.031
R12839 VDD.n6470 VDD.n6469 0.031
R12840 VDD.n6484 VDD.n6483 0.031
R12841 VDD.n6508 VDD.n6502 0.031
R12842 VDD.n6527 VDD.n6526 0.031
R12843 VDD.n6615 VDD.n6547 0.031
R12844 VDD.n6634 VDD.n6633 0.031
R12845 VDD.n6657 VDD.n6651 0.031
R12846 VDD.n6677 VDD.n6676 0.031
R12847 VDD.n6832 VDD.n6831 0.031
R12848 VDD.n6846 VDD.n6845 0.031
R12849 VDD.n6870 VDD.n6864 0.031
R12850 VDD.n6889 VDD.n6888 0.031
R12851 VDD.n6977 VDD.n6909 0.031
R12852 VDD.n6996 VDD.n6995 0.031
R12853 VDD.n7019 VDD.n7013 0.031
R12854 VDD.n7039 VDD.n7038 0.031
R12855 VDD.n7194 VDD.n7193 0.031
R12856 VDD.n7208 VDD.n7207 0.031
R12857 VDD.n7232 VDD.n7226 0.031
R12858 VDD.n7251 VDD.n7250 0.031
R12859 VDD.n7339 VDD.n7271 0.031
R12860 VDD.n7358 VDD.n7357 0.031
R12861 VDD.n7381 VDD.n7375 0.031
R12862 VDD.n7401 VDD.n7400 0.031
R12863 VDD.n7556 VDD.n7555 0.031
R12864 VDD.n7570 VDD.n7569 0.031
R12865 VDD.n7594 VDD.n7588 0.031
R12866 VDD.n7613 VDD.n7612 0.031
R12867 VDD.n7701 VDD.n7633 0.031
R12868 VDD.n7720 VDD.n7719 0.031
R12869 VDD.n7743 VDD.n7737 0.031
R12870 VDD.n7763 VDD.n7762 0.031
R12871 VDD.n7918 VDD.n7917 0.031
R12872 VDD.n7932 VDD.n7931 0.031
R12873 VDD.n7956 VDD.n7950 0.031
R12874 VDD.n7975 VDD.n7974 0.031
R12875 VDD.n8063 VDD.n7995 0.031
R12876 VDD.n8082 VDD.n8081 0.031
R12877 VDD.n8105 VDD.n8099 0.031
R12878 VDD.n8125 VDD.n8124 0.031
R12879 VDD.n8280 VDD.n8279 0.031
R12880 VDD.n8294 VDD.n8293 0.031
R12881 VDD.n8318 VDD.n8312 0.031
R12882 VDD.n8337 VDD.n8336 0.031
R12883 VDD.n8425 VDD.n8357 0.031
R12884 VDD.n8444 VDD.n8443 0.031
R12885 VDD.n8467 VDD.n8461 0.031
R12886 VDD.n8487 VDD.n8486 0.031
R12887 VDD.n8642 VDD.n8641 0.031
R12888 VDD.n8656 VDD.n8655 0.031
R12889 VDD.n8680 VDD.n8674 0.031
R12890 VDD.n8699 VDD.n8698 0.031
R12891 VDD.n8787 VDD.n8719 0.031
R12892 VDD.n8806 VDD.n8805 0.031
R12893 VDD.n8829 VDD.n8823 0.031
R12894 VDD.n8849 VDD.n8848 0.031
R12895 VDD.n9004 VDD.n9003 0.031
R12896 VDD.n9018 VDD.n9017 0.031
R12897 VDD.n9042 VDD.n9036 0.031
R12898 VDD.n9061 VDD.n9060 0.031
R12899 VDD.n9149 VDD.n9081 0.031
R12900 VDD.n9168 VDD.n9167 0.031
R12901 VDD.n9191 VDD.n9185 0.031
R12902 VDD.n9211 VDD.n9210 0.031
R12903 VDD.n9366 VDD.n9365 0.031
R12904 VDD.n9380 VDD.n9379 0.031
R12905 VDD.n9404 VDD.n9398 0.031
R12906 VDD.n9423 VDD.n9422 0.031
R12907 VDD.n9511 VDD.n9443 0.031
R12908 VDD.n9530 VDD.n9529 0.031
R12909 VDD.n9553 VDD.n9547 0.031
R12910 VDD.n9573 VDD.n9572 0.031
R12911 VDD.n9728 VDD.n9727 0.031
R12912 VDD.n9742 VDD.n9741 0.031
R12913 VDD.n9766 VDD.n9760 0.031
R12914 VDD.n9785 VDD.n9784 0.031
R12915 VDD.n9873 VDD.n9805 0.031
R12916 VDD.n9892 VDD.n9891 0.031
R12917 VDD.n9915 VDD.n9909 0.031
R12918 VDD.n9935 VDD.n9934 0.031
R12919 VDD.n173 VDD.n172 0.03
R12920 VDD.n2728 VDD.n2727 0.03
R12921 VDD.n116 VDD.n115 0.03
R12922 VDD.n108 VDD.n107 0.03
R12923 VDD.n2701 VDD.n2700 0.03
R12924 VDD.n5359 VDD.n5358 0.03
R12925 VDD.n5498 VDD.n5495 0.03
R12926 VDD.n5511 VDD.n5508 0.03
R12927 VDD.n5634 VDD.n5633 0.03
R12928 VDD.n5651 VDD.n5650 0.03
R12929 VDD.n5457 VDD.n5456 0.03
R12930 VDD.n5581 VDD.n5580 0.03
R12931 VDD.n5720 VDD.n5719 0.03
R12932 VDD.n5859 VDD.n5856 0.03
R12933 VDD.n5872 VDD.n5869 0.03
R12934 VDD.n5995 VDD.n5994 0.03
R12935 VDD.n6012 VDD.n6011 0.03
R12936 VDD.n5818 VDD.n5817 0.03
R12937 VDD.n5942 VDD.n5941 0.03
R12938 VDD.n6082 VDD.n6081 0.03
R12939 VDD.n6221 VDD.n6218 0.03
R12940 VDD.n6234 VDD.n6231 0.03
R12941 VDD.n6357 VDD.n6356 0.03
R12942 VDD.n6374 VDD.n6373 0.03
R12943 VDD.n6180 VDD.n6179 0.03
R12944 VDD.n6304 VDD.n6303 0.03
R12945 VDD.n6444 VDD.n6443 0.03
R12946 VDD.n6583 VDD.n6580 0.03
R12947 VDD.n6596 VDD.n6593 0.03
R12948 VDD.n6719 VDD.n6718 0.03
R12949 VDD.n6736 VDD.n6735 0.03
R12950 VDD.n6542 VDD.n6541 0.03
R12951 VDD.n6666 VDD.n6665 0.03
R12952 VDD.n6806 VDD.n6805 0.03
R12953 VDD.n6945 VDD.n6942 0.03
R12954 VDD.n6958 VDD.n6955 0.03
R12955 VDD.n7081 VDD.n7080 0.03
R12956 VDD.n7098 VDD.n7097 0.03
R12957 VDD.n6904 VDD.n6903 0.03
R12958 VDD.n7028 VDD.n7027 0.03
R12959 VDD.n7168 VDD.n7167 0.03
R12960 VDD.n7307 VDD.n7304 0.03
R12961 VDD.n7320 VDD.n7317 0.03
R12962 VDD.n7443 VDD.n7442 0.03
R12963 VDD.n7460 VDD.n7459 0.03
R12964 VDD.n7266 VDD.n7265 0.03
R12965 VDD.n7390 VDD.n7389 0.03
R12966 VDD.n7530 VDD.n7529 0.03
R12967 VDD.n7669 VDD.n7666 0.03
R12968 VDD.n7682 VDD.n7679 0.03
R12969 VDD.n7805 VDD.n7804 0.03
R12970 VDD.n7822 VDD.n7821 0.03
R12971 VDD.n7628 VDD.n7627 0.03
R12972 VDD.n7752 VDD.n7751 0.03
R12973 VDD.n7892 VDD.n7891 0.03
R12974 VDD.n8031 VDD.n8028 0.03
R12975 VDD.n8044 VDD.n8041 0.03
R12976 VDD.n8167 VDD.n8166 0.03
R12977 VDD.n8184 VDD.n8183 0.03
R12978 VDD.n7990 VDD.n7989 0.03
R12979 VDD.n8114 VDD.n8113 0.03
R12980 VDD.n8254 VDD.n8253 0.03
R12981 VDD.n8393 VDD.n8390 0.03
R12982 VDD.n8406 VDD.n8403 0.03
R12983 VDD.n8529 VDD.n8528 0.03
R12984 VDD.n8546 VDD.n8545 0.03
R12985 VDD.n8352 VDD.n8351 0.03
R12986 VDD.n8476 VDD.n8475 0.03
R12987 VDD.n8616 VDD.n8615 0.03
R12988 VDD.n8755 VDD.n8752 0.03
R12989 VDD.n8768 VDD.n8765 0.03
R12990 VDD.n8891 VDD.n8890 0.03
R12991 VDD.n8908 VDD.n8907 0.03
R12992 VDD.n8714 VDD.n8713 0.03
R12993 VDD.n8838 VDD.n8837 0.03
R12994 VDD.n8978 VDD.n8977 0.03
R12995 VDD.n9117 VDD.n9114 0.03
R12996 VDD.n9130 VDD.n9127 0.03
R12997 VDD.n9253 VDD.n9252 0.03
R12998 VDD.n9270 VDD.n9269 0.03
R12999 VDD.n9076 VDD.n9075 0.03
R13000 VDD.n9200 VDD.n9199 0.03
R13001 VDD.n9340 VDD.n9339 0.03
R13002 VDD.n9479 VDD.n9476 0.03
R13003 VDD.n9492 VDD.n9489 0.03
R13004 VDD.n9615 VDD.n9614 0.03
R13005 VDD.n9632 VDD.n9631 0.03
R13006 VDD.n9438 VDD.n9437 0.03
R13007 VDD.n9562 VDD.n9561 0.03
R13008 VDD.n9702 VDD.n9701 0.03
R13009 VDD.n9841 VDD.n9838 0.03
R13010 VDD.n9854 VDD.n9851 0.03
R13011 VDD.n9977 VDD.n9976 0.03
R13012 VDD.n9994 VDD.n9993 0.03
R13013 VDD.n9800 VDD.n9799 0.03
R13014 VDD.n9924 VDD.n9923 0.03
R13015 VDD.n10314 VDD.n10312 0.03
R13016 VDD.n10264 VDD.n10262 0.03
R13017 VDD.n10195 VDD.n10193 0.03
R13018 VDD.n10147 VDD.n10145 0.03
R13019 VDD.n11571 VDD.n11570 0.03
R13020 VDD.n11735 VDD.n11734 0.03
R13021 VDD.n10801 VDD.n10800 0.03
R13022 VDD.n10966 VDD.n10965 0.03
R13023 VDD.n10934 VDD.n10933 0.03
R13024 VDD.n11070 VDD.n11069 0.03
R13025 VDD.n10999 VDD.n10998 0.03
R13026 VDD.n11166 VDD.n11155 0.03
R13027 VDD.n11180 VDD.n11169 0.03
R13028 VDD.n11152 VDD.n11141 0.03
R13029 VDD.n10828 VDD.n10827 0.03
R13030 VDD.n10745 VDD.n10744 0.03
R13031 VDD.n10761 VDD.n10760 0.03
R13032 VDD.n11688 VDD.n11687 0.03
R13033 VDD.n11836 VDD.n11835 0.03
R13034 VDD.n11767 VDD.n11766 0.03
R13035 VDD.n11924 VDD.n11913 0.03
R13036 VDD.n11937 VDD.n11927 0.03
R13037 VDD.n11910 VDD.n11900 0.03
R13038 VDD.n11608 VDD.n11607 0.03
R13039 VDD.n11516 VDD.n11515 0.03
R13040 VDD.n11531 VDD.n11530 0.03
R13041 VDD.n193 VDD.n192 0.03
R13042 VDD.n2692 VDD.n2691 0.03
R13043 VDD.n5129 VDD.n5128 0.03
R13044 VDD.n193 VDD.n190 0.03
R13045 VDD.n5143 VDD.n5142 0.029
R13046 VDD.n2593 VDD.n2529 0.029
R13047 VDD.n5143 VDD.n5132 0.029
R13048 VDD.n5383 VDD.n5317 0.029
R13049 VDD.n5744 VDD.n5678 0.029
R13050 VDD.n6106 VDD.n6040 0.029
R13051 VDD.n6468 VDD.n6402 0.029
R13052 VDD.n6830 VDD.n6764 0.029
R13053 VDD.n7192 VDD.n7126 0.029
R13054 VDD.n7554 VDD.n7488 0.029
R13055 VDD.n7916 VDD.n7850 0.029
R13056 VDD.n8278 VDD.n8212 0.029
R13057 VDD.n8640 VDD.n8574 0.029
R13058 VDD.n9002 VDD.n8936 0.029
R13059 VDD.n9364 VDD.n9298 0.029
R13060 VDD.n9726 VDD.n9660 0.029
R13061 VDD.n10661 VDD.n10659 0.029
R13062 VDD.n10611 VDD.n10609 0.029
R13063 VDD.n10541 VDD.n10539 0.029
R13064 VDD.n10493 VDD.n10491 0.029
R13065 VDD.n5305 VDD.n5299 0.029
R13066 VDD.n11010 VDD.n11001 0.029
R13067 VDD.n11106 VDD.n11105 0.028
R13068 VDD.n11073 VDD.n11072 0.028
R13069 VDD.n11841 VDD.n11838 0.028
R13070 VDD.n11778 VDD.n11769 0.028
R13071 VDD.n5041 VDD.n5031 0.028
R13072 VDD.n4966 VDD.n4964 0.028
R13073 VDD.n4810 VDD.n4800 0.028
R13074 VDD.n4735 VDD.n4733 0.028
R13075 VDD.n4613 VDD.n4612 0.028
R13076 VDD.n4576 VDD.n4575 0.028
R13077 VDD.n2948 VDD.n2947 0.028
R13078 VDD.n2824 VDD.n2822 0.028
R13079 VDD.n2964 VDD.n2963 0.028
R13080 VDD.n3044 VDD.n3043 0.028
R13081 VDD.n3202 VDD.n3201 0.028
R13082 VDD.n3281 VDD.n3280 0.028
R13083 VDD.n3439 VDD.n3438 0.028
R13084 VDD.n3519 VDD.n3518 0.028
R13085 VDD.n3677 VDD.n3676 0.028
R13086 VDD.n3756 VDD.n3755 0.028
R13087 VDD.n3914 VDD.n3913 0.028
R13088 VDD.n3994 VDD.n3993 0.028
R13089 VDD.n4152 VDD.n4151 0.028
R13090 VDD.n4231 VDD.n4230 0.028
R13091 VDD.n4389 VDD.n4388 0.028
R13092 VDD.n4474 VDD.n4473 0.028
R13093 VDD.n365 VDD.n364 0.028
R13094 VDD.n248 VDD.n246 0.028
R13095 VDD.n2007 VDD.n2006 0.028
R13096 VDD.n1970 VDD.n1969 0.028
R13097 VDD.n381 VDD.n380 0.028
R13098 VDD.n464 VDD.n463 0.028
R13099 VDD.n615 VDD.n614 0.028
R13100 VDD.n697 VDD.n696 0.028
R13101 VDD.n848 VDD.n847 0.028
R13102 VDD.n931 VDD.n930 0.028
R13103 VDD.n1082 VDD.n1081 0.028
R13104 VDD.n1164 VDD.n1163 0.028
R13105 VDD.n1315 VDD.n1314 0.028
R13106 VDD.n1398 VDD.n1397 0.028
R13107 VDD.n1549 VDD.n1548 0.028
R13108 VDD.n1631 VDD.n1630 0.028
R13109 VDD.n1782 VDD.n1781 0.028
R13110 VDD.n1869 VDD.n1868 0.028
R13111 VDD.n2131 VDD.n2129 0.028
R13112 VDD.n2206 VDD.n2196 0.028
R13113 VDD.n2362 VDD.n2360 0.028
R13114 VDD.n2437 VDD.n2427 0.028
R13115 VDD.n2589 VDD.n2588 0.028
R13116 VDD.n2568 VDD.n2567 0.028
R13117 VDD.n2754 VDD.n2748 0.028
R13118 VDD.n2590 VDD.n2538 0.028
R13119 VDD.n2531 VDD.n2530 0.028
R13120 VDD.n171 VDD.n170 0.028
R13121 VDD.n2615 VDD.n2614 0.028
R13122 VDD.n2630 VDD.n2629 0.028
R13123 VDD.n2695 VDD.n2694 0.028
R13124 VDD.n2755 VDD.n2708 0.028
R13125 VDD.n5370 VDD.n5369 0.028
R13126 VDD.n5485 VDD.n5484 0.028
R13127 VDD.n5528 VDD.n5527 0.028
R13128 VDD.n5520 VDD.n5519 0.028
R13129 VDD.n5413 VDD.n5412 0.028
R13130 VDD.n5419 VDD.n5418 0.028
R13131 VDD.n5448 VDD.n5447 0.028
R13132 VDD.n5539 VDD.n5538 0.028
R13133 VDD.n5731 VDD.n5730 0.028
R13134 VDD.n5846 VDD.n5845 0.028
R13135 VDD.n5889 VDD.n5888 0.028
R13136 VDD.n5881 VDD.n5880 0.028
R13137 VDD.n5774 VDD.n5773 0.028
R13138 VDD.n5780 VDD.n5779 0.028
R13139 VDD.n5809 VDD.n5808 0.028
R13140 VDD.n5900 VDD.n5899 0.028
R13141 VDD.n6093 VDD.n6092 0.028
R13142 VDD.n6208 VDD.n6207 0.028
R13143 VDD.n6251 VDD.n6250 0.028
R13144 VDD.n6243 VDD.n6242 0.028
R13145 VDD.n6136 VDD.n6135 0.028
R13146 VDD.n6142 VDD.n6141 0.028
R13147 VDD.n6171 VDD.n6170 0.028
R13148 VDD.n6262 VDD.n6261 0.028
R13149 VDD.n6455 VDD.n6454 0.028
R13150 VDD.n6570 VDD.n6569 0.028
R13151 VDD.n6613 VDD.n6612 0.028
R13152 VDD.n6605 VDD.n6604 0.028
R13153 VDD.n6498 VDD.n6497 0.028
R13154 VDD.n6504 VDD.n6503 0.028
R13155 VDD.n6533 VDD.n6532 0.028
R13156 VDD.n6624 VDD.n6623 0.028
R13157 VDD.n6817 VDD.n6816 0.028
R13158 VDD.n6932 VDD.n6931 0.028
R13159 VDD.n6975 VDD.n6974 0.028
R13160 VDD.n6967 VDD.n6966 0.028
R13161 VDD.n6860 VDD.n6859 0.028
R13162 VDD.n6866 VDD.n6865 0.028
R13163 VDD.n6895 VDD.n6894 0.028
R13164 VDD.n6986 VDD.n6985 0.028
R13165 VDD.n7179 VDD.n7178 0.028
R13166 VDD.n7294 VDD.n7293 0.028
R13167 VDD.n7337 VDD.n7336 0.028
R13168 VDD.n7329 VDD.n7328 0.028
R13169 VDD.n7222 VDD.n7221 0.028
R13170 VDD.n7228 VDD.n7227 0.028
R13171 VDD.n7257 VDD.n7256 0.028
R13172 VDD.n7348 VDD.n7347 0.028
R13173 VDD.n7541 VDD.n7540 0.028
R13174 VDD.n7656 VDD.n7655 0.028
R13175 VDD.n7699 VDD.n7698 0.028
R13176 VDD.n7691 VDD.n7690 0.028
R13177 VDD.n7584 VDD.n7583 0.028
R13178 VDD.n7590 VDD.n7589 0.028
R13179 VDD.n7619 VDD.n7618 0.028
R13180 VDD.n7710 VDD.n7709 0.028
R13181 VDD.n7903 VDD.n7902 0.028
R13182 VDD.n8018 VDD.n8017 0.028
R13183 VDD.n8061 VDD.n8060 0.028
R13184 VDD.n8053 VDD.n8052 0.028
R13185 VDD.n7946 VDD.n7945 0.028
R13186 VDD.n7952 VDD.n7951 0.028
R13187 VDD.n7981 VDD.n7980 0.028
R13188 VDD.n8072 VDD.n8071 0.028
R13189 VDD.n8265 VDD.n8264 0.028
R13190 VDD.n8380 VDD.n8379 0.028
R13191 VDD.n8423 VDD.n8422 0.028
R13192 VDD.n8415 VDD.n8414 0.028
R13193 VDD.n8308 VDD.n8307 0.028
R13194 VDD.n8314 VDD.n8313 0.028
R13195 VDD.n8343 VDD.n8342 0.028
R13196 VDD.n8434 VDD.n8433 0.028
R13197 VDD.n8627 VDD.n8626 0.028
R13198 VDD.n8742 VDD.n8741 0.028
R13199 VDD.n8785 VDD.n8784 0.028
R13200 VDD.n8777 VDD.n8776 0.028
R13201 VDD.n8670 VDD.n8669 0.028
R13202 VDD.n8676 VDD.n8675 0.028
R13203 VDD.n8705 VDD.n8704 0.028
R13204 VDD.n8796 VDD.n8795 0.028
R13205 VDD.n8989 VDD.n8988 0.028
R13206 VDD.n9104 VDD.n9103 0.028
R13207 VDD.n9147 VDD.n9146 0.028
R13208 VDD.n9139 VDD.n9138 0.028
R13209 VDD.n9032 VDD.n9031 0.028
R13210 VDD.n9038 VDD.n9037 0.028
R13211 VDD.n9067 VDD.n9066 0.028
R13212 VDD.n9158 VDD.n9157 0.028
R13213 VDD.n9351 VDD.n9350 0.028
R13214 VDD.n9466 VDD.n9465 0.028
R13215 VDD.n9509 VDD.n9508 0.028
R13216 VDD.n9501 VDD.n9500 0.028
R13217 VDD.n9394 VDD.n9393 0.028
R13218 VDD.n9400 VDD.n9399 0.028
R13219 VDD.n9429 VDD.n9428 0.028
R13220 VDD.n9520 VDD.n9519 0.028
R13221 VDD.n9713 VDD.n9712 0.028
R13222 VDD.n9828 VDD.n9827 0.028
R13223 VDD.n9871 VDD.n9870 0.028
R13224 VDD.n9863 VDD.n9862 0.028
R13225 VDD.n9756 VDD.n9755 0.028
R13226 VDD.n9762 VDD.n9761 0.028
R13227 VDD.n9791 VDD.n9790 0.028
R13228 VDD.n9882 VDD.n9881 0.028
R13229 VDD.n11561 VDD.n11560 0.028
R13230 VDD.n11557 VDD.n11556 0.028
R13231 VDD.n11745 VDD.n11744 0.028
R13232 VDD.n10791 VDD.n10790 0.028
R13233 VDD.n10787 VDD.n10786 0.028
R13234 VDD.n10976 VDD.n10975 0.028
R13235 VDD.n10948 VDD.n10947 0.028
R13236 VDD.n11037 VDD.n11036 0.028
R13237 VDD.n11040 VDD.n11039 0.028
R13238 VDD.n11138 VDD.n11137 0.028
R13239 VDD.n10841 VDD.n10840 0.028
R13240 VDD.n10825 VDD.n10824 0.028
R13241 VDD.n10732 VDD.n10731 0.028
R13242 VDD.n10759 VDD.n10748 0.028
R13243 VDD.n11714 VDD.n11713 0.028
R13244 VDD.n11804 VDD.n11803 0.028
R13245 VDD.n11807 VDD.n11806 0.028
R13246 VDD.n11897 VDD.n11886 0.028
R13247 VDD.n11620 VDD.n11619 0.028
R13248 VDD.n11605 VDD.n11604 0.028
R13249 VDD.n11503 VDD.n11502 0.028
R13250 VDD.n11529 VDD.n11519 0.028
R13251 VDD.n2628 VDD.n2627 0.027
R13252 VDD.n5392 VDD.n5388 0.027
R13253 VDD.n5434 VDD.n5430 0.027
R13254 VDD.n5541 VDD.n5537 0.027
R13255 VDD.n5583 VDD.n5579 0.027
R13256 VDD.n5753 VDD.n5749 0.027
R13257 VDD.n5795 VDD.n5791 0.027
R13258 VDD.n5902 VDD.n5898 0.027
R13259 VDD.n5944 VDD.n5940 0.027
R13260 VDD.n6115 VDD.n6111 0.027
R13261 VDD.n6157 VDD.n6153 0.027
R13262 VDD.n6264 VDD.n6260 0.027
R13263 VDD.n6306 VDD.n6302 0.027
R13264 VDD.n6477 VDD.n6473 0.027
R13265 VDD.n6519 VDD.n6515 0.027
R13266 VDD.n6626 VDD.n6622 0.027
R13267 VDD.n6668 VDD.n6664 0.027
R13268 VDD.n6839 VDD.n6835 0.027
R13269 VDD.n6881 VDD.n6877 0.027
R13270 VDD.n6988 VDD.n6984 0.027
R13271 VDD.n7030 VDD.n7026 0.027
R13272 VDD.n7201 VDD.n7197 0.027
R13273 VDD.n7243 VDD.n7239 0.027
R13274 VDD.n7350 VDD.n7346 0.027
R13275 VDD.n7392 VDD.n7388 0.027
R13276 VDD.n7563 VDD.n7559 0.027
R13277 VDD.n7605 VDD.n7601 0.027
R13278 VDD.n7712 VDD.n7708 0.027
R13279 VDD.n7754 VDD.n7750 0.027
R13280 VDD.n7925 VDD.n7921 0.027
R13281 VDD.n7967 VDD.n7963 0.027
R13282 VDD.n8074 VDD.n8070 0.027
R13283 VDD.n8116 VDD.n8112 0.027
R13284 VDD.n8287 VDD.n8283 0.027
R13285 VDD.n8329 VDD.n8325 0.027
R13286 VDD.n8436 VDD.n8432 0.027
R13287 VDD.n8478 VDD.n8474 0.027
R13288 VDD.n8649 VDD.n8645 0.027
R13289 VDD.n8691 VDD.n8687 0.027
R13290 VDD.n8798 VDD.n8794 0.027
R13291 VDD.n8840 VDD.n8836 0.027
R13292 VDD.n9011 VDD.n9007 0.027
R13293 VDD.n9053 VDD.n9049 0.027
R13294 VDD.n9160 VDD.n9156 0.027
R13295 VDD.n9202 VDD.n9198 0.027
R13296 VDD.n9373 VDD.n9369 0.027
R13297 VDD.n9415 VDD.n9411 0.027
R13298 VDD.n9522 VDD.n9518 0.027
R13299 VDD.n9564 VDD.n9560 0.027
R13300 VDD.n9735 VDD.n9731 0.027
R13301 VDD.n9777 VDD.n9773 0.027
R13302 VDD.n9884 VDD.n9880 0.027
R13303 VDD.n9926 VDD.n9922 0.027
R13304 VDD.n11135 VDD.n11134 0.026
R13305 VDD.n11884 VDD.n11883 0.026
R13306 VDD.n5073 VDD.n5071 0.026
R13307 VDD.n4926 VDD.n4924 0.026
R13308 VDD.n4842 VDD.n4840 0.026
R13309 VDD.n4695 VDD.n4693 0.026
R13310 VDD.n4600 VDD.n4599 0.026
R13311 VDD.n4595 VDD.n4594 0.026
R13312 VDD.n2816 VDD.n2815 0.026
R13313 VDD.n2934 VDD.n2933 0.026
R13314 VDD.n2896 VDD.n2868 0.026
R13315 VDD.n3085 VDD.n3084 0.026
R13316 VDD.n3172 VDD.n3160 0.026
R13317 VDD.n3323 VDD.n3322 0.026
R13318 VDD.n3409 VDD.n3397 0.026
R13319 VDD.n3560 VDD.n3559 0.026
R13320 VDD.n3647 VDD.n3635 0.026
R13321 VDD.n3798 VDD.n3797 0.026
R13322 VDD.n3884 VDD.n3872 0.026
R13323 VDD.n4035 VDD.n4034 0.026
R13324 VDD.n4122 VDD.n4110 0.026
R13325 VDD.n4273 VDD.n4272 0.026
R13326 VDD.n4359 VDD.n4347 0.026
R13327 VDD.n4533 VDD.n4532 0.026
R13328 VDD.n240 VDD.n239 0.026
R13329 VDD.n352 VDD.n351 0.026
R13330 VDD.n1994 VDD.n1993 0.026
R13331 VDD.n1989 VDD.n1988 0.026
R13332 VDD.n310 VDD.n281 0.026
R13333 VDD.n505 VDD.n504 0.026
R13334 VDD.n585 VDD.n573 0.026
R13335 VDD.n739 VDD.n738 0.026
R13336 VDD.n818 VDD.n806 0.026
R13337 VDD.n972 VDD.n971 0.026
R13338 VDD.n1052 VDD.n1040 0.026
R13339 VDD.n1206 VDD.n1205 0.026
R13340 VDD.n1285 VDD.n1273 0.026
R13341 VDD.n1439 VDD.n1438 0.026
R13342 VDD.n1519 VDD.n1507 0.026
R13343 VDD.n1673 VDD.n1672 0.026
R13344 VDD.n1752 VDD.n1740 0.026
R13345 VDD.n1924 VDD.n1923 0.026
R13346 VDD.n2091 VDD.n2089 0.026
R13347 VDD.n2238 VDD.n2236 0.026
R13348 VDD.n2322 VDD.n2320 0.026
R13349 VDD.n2469 VDD.n2467 0.026
R13350 VDD.n154 VDD.n153 0.026
R13351 VDD.n5253 VDD.n5252 0.026
R13352 VDD.n2651 VDD.n2650 0.026
R13353 VDD.n5123 VDD.n5122 0.026
R13354 VDD.n176 VDD.n175 0.026
R13355 VDD.n5477 VDD.n5476 0.026
R13356 VDD.n5316 VDD.n5315 0.026
R13357 VDD.n5553 VDD.n5552 0.026
R13358 VDD.n5555 VDD.n5554 0.026
R13359 VDD.n5838 VDD.n5837 0.026
R13360 VDD.n5677 VDD.n5676 0.026
R13361 VDD.n5914 VDD.n5913 0.026
R13362 VDD.n5916 VDD.n5915 0.026
R13363 VDD.n6200 VDD.n6199 0.026
R13364 VDD.n6039 VDD.n6038 0.026
R13365 VDD.n6276 VDD.n6275 0.026
R13366 VDD.n6278 VDD.n6277 0.026
R13367 VDD.n6562 VDD.n6561 0.026
R13368 VDD.n6401 VDD.n6400 0.026
R13369 VDD.n6638 VDD.n6637 0.026
R13370 VDD.n6640 VDD.n6639 0.026
R13371 VDD.n6924 VDD.n6923 0.026
R13372 VDD.n6763 VDD.n6762 0.026
R13373 VDD.n7000 VDD.n6999 0.026
R13374 VDD.n7002 VDD.n7001 0.026
R13375 VDD.n7286 VDD.n7285 0.026
R13376 VDD.n7125 VDD.n7124 0.026
R13377 VDD.n7362 VDD.n7361 0.026
R13378 VDD.n7364 VDD.n7363 0.026
R13379 VDD.n7648 VDD.n7647 0.026
R13380 VDD.n7487 VDD.n7486 0.026
R13381 VDD.n7724 VDD.n7723 0.026
R13382 VDD.n7726 VDD.n7725 0.026
R13383 VDD.n8010 VDD.n8009 0.026
R13384 VDD.n7849 VDD.n7848 0.026
R13385 VDD.n8086 VDD.n8085 0.026
R13386 VDD.n8088 VDD.n8087 0.026
R13387 VDD.n8372 VDD.n8371 0.026
R13388 VDD.n8211 VDD.n8210 0.026
R13389 VDD.n8448 VDD.n8447 0.026
R13390 VDD.n8450 VDD.n8449 0.026
R13391 VDD.n8734 VDD.n8733 0.026
R13392 VDD.n8573 VDD.n8572 0.026
R13393 VDD.n8810 VDD.n8809 0.026
R13394 VDD.n8812 VDD.n8811 0.026
R13395 VDD.n9096 VDD.n9095 0.026
R13396 VDD.n8935 VDD.n8934 0.026
R13397 VDD.n9172 VDD.n9171 0.026
R13398 VDD.n9174 VDD.n9173 0.026
R13399 VDD.n9458 VDD.n9457 0.026
R13400 VDD.n9297 VDD.n9296 0.026
R13401 VDD.n9534 VDD.n9533 0.026
R13402 VDD.n9536 VDD.n9535 0.026
R13403 VDD.n9820 VDD.n9819 0.026
R13404 VDD.n9659 VDD.n9658 0.026
R13405 VDD.n9896 VDD.n9895 0.026
R13406 VDD.n9898 VDD.n9897 0.026
R13407 VDD.n11575 VDD.n11574 0.026
R13408 VDD.n11731 VDD.n11730 0.026
R13409 VDD.n10805 VDD.n10804 0.026
R13410 VDD.n10962 VDD.n10961 0.026
R13411 VDD.n10946 VDD.n10945 0.026
R13412 VDD.n11054 VDD.n11053 0.026
R13413 VDD.n11058 VDD.n11057 0.026
R13414 VDD.n10845 VDD.n10844 0.026
R13415 VDD.n11712 VDD.n11702 0.026
R13416 VDD.n11820 VDD.n11819 0.026
R13417 VDD.n11824 VDD.n11823 0.026
R13418 VDD.n11626 VDD.n11623 0.026
R13419 VDD.n10997 VDD.n10996 0.026
R13420 VDD.n11765 VDD.n11754 0.025
R13421 VDD.n10326 VDD.n10324 0.025
R13422 VDD.n10251 VDD.n10249 0.025
R13423 VDD.n10207 VDD.n10205 0.025
R13424 VDD.n10135 VDD.n10133 0.025
R13425 VDD.n10673 VDD.n10671 0.025
R13426 VDD.n10598 VDD.n10596 0.025
R13427 VDD.n10553 VDD.n10551 0.025
R13428 VDD.n10481 VDD.n10479 0.025
R13429 VDD.n73 VDD.n71 0.024
R13430 VDD.n52 VDD.n50 0.024
R13431 VDD.n5055 VDD.n5045 0.024
R13432 VDD.n4952 VDD.n4950 0.024
R13433 VDD.n4824 VDD.n4814 0.024
R13434 VDD.n4721 VDD.n4719 0.024
R13435 VDD.n2917 VDD.n2916 0.024
R13436 VDD.n3058 VDD.n3057 0.024
R13437 VDD.n3188 VDD.n3187 0.024
R13438 VDD.n3295 VDD.n3294 0.024
R13439 VDD.n3425 VDD.n3424 0.024
R13440 VDD.n3533 VDD.n3532 0.024
R13441 VDD.n3663 VDD.n3662 0.024
R13442 VDD.n3770 VDD.n3769 0.024
R13443 VDD.n3900 VDD.n3899 0.024
R13444 VDD.n4008 VDD.n4007 0.024
R13445 VDD.n4138 VDD.n4137 0.024
R13446 VDD.n4245 VDD.n4244 0.024
R13447 VDD.n4375 VDD.n4374 0.024
R13448 VDD.n4494 VDD.n4493 0.024
R13449 VDD.n330 VDD.n329 0.024
R13450 VDD.n478 VDD.n477 0.024
R13451 VDD.n601 VDD.n600 0.024
R13452 VDD.n711 VDD.n710 0.024
R13453 VDD.n834 VDD.n833 0.024
R13454 VDD.n945 VDD.n944 0.024
R13455 VDD.n1068 VDD.n1067 0.024
R13456 VDD.n1178 VDD.n1177 0.024
R13457 VDD.n1301 VDD.n1300 0.024
R13458 VDD.n1412 VDD.n1411 0.024
R13459 VDD.n1535 VDD.n1534 0.024
R13460 VDD.n1645 VDD.n1644 0.024
R13461 VDD.n1768 VDD.n1767 0.024
R13462 VDD.n1887 VDD.n1886 0.024
R13463 VDD.n2117 VDD.n2115 0.024
R13464 VDD.n2220 VDD.n2210 0.024
R13465 VDD.n2348 VDD.n2346 0.024
R13466 VDD.n2451 VDD.n2441 0.024
R13467 VDD.n2519 VDD.n2518 0.024
R13468 VDD.n5188 VDD.n5187 0.024
R13469 VDD.n5235 VDD.n5234 0.024
R13470 VDD.n2536 VDD.n2535 0.024
R13471 VDD.n2610 VDD.n2609 0.024
R13472 VDD.n5312 VDD.n5311 0.024
R13473 VDD.n5310 VDD.n5309 0.024
R13474 VDD.n5397 VDD.n5396 0.024
R13475 VDD.n5429 VDD.n5427 0.024
R13476 VDD.n5440 VDD.n5438 0.024
R13477 VDD.n5536 VDD.n5534 0.024
R13478 VDD.n5547 VDD.n5545 0.024
R13479 VDD.n5578 VDD.n5576 0.024
R13480 VDD.n5596 VDD.n5595 0.024
R13481 VDD.n5673 VDD.n5672 0.024
R13482 VDD.n5671 VDD.n5670 0.024
R13483 VDD.n5758 VDD.n5757 0.024
R13484 VDD.n5790 VDD.n5788 0.024
R13485 VDD.n5801 VDD.n5799 0.024
R13486 VDD.n5897 VDD.n5895 0.024
R13487 VDD.n5908 VDD.n5906 0.024
R13488 VDD.n5939 VDD.n5937 0.024
R13489 VDD.n5957 VDD.n5956 0.024
R13490 VDD.n6035 VDD.n6034 0.024
R13491 VDD.n6033 VDD.n6032 0.024
R13492 VDD.n6120 VDD.n6119 0.024
R13493 VDD.n6152 VDD.n6150 0.024
R13494 VDD.n6163 VDD.n6161 0.024
R13495 VDD.n6259 VDD.n6257 0.024
R13496 VDD.n6270 VDD.n6268 0.024
R13497 VDD.n6301 VDD.n6299 0.024
R13498 VDD.n6319 VDD.n6318 0.024
R13499 VDD.n6397 VDD.n6396 0.024
R13500 VDD.n6395 VDD.n6394 0.024
R13501 VDD.n6482 VDD.n6481 0.024
R13502 VDD.n6514 VDD.n6512 0.024
R13503 VDD.n6525 VDD.n6523 0.024
R13504 VDD.n6621 VDD.n6619 0.024
R13505 VDD.n6632 VDD.n6630 0.024
R13506 VDD.n6663 VDD.n6661 0.024
R13507 VDD.n6681 VDD.n6680 0.024
R13508 VDD.n6759 VDD.n6758 0.024
R13509 VDD.n6757 VDD.n6756 0.024
R13510 VDD.n6844 VDD.n6843 0.024
R13511 VDD.n6876 VDD.n6874 0.024
R13512 VDD.n6887 VDD.n6885 0.024
R13513 VDD.n6983 VDD.n6981 0.024
R13514 VDD.n6994 VDD.n6992 0.024
R13515 VDD.n7025 VDD.n7023 0.024
R13516 VDD.n7043 VDD.n7042 0.024
R13517 VDD.n7121 VDD.n7120 0.024
R13518 VDD.n7119 VDD.n7118 0.024
R13519 VDD.n7206 VDD.n7205 0.024
R13520 VDD.n7238 VDD.n7236 0.024
R13521 VDD.n7249 VDD.n7247 0.024
R13522 VDD.n7345 VDD.n7343 0.024
R13523 VDD.n7356 VDD.n7354 0.024
R13524 VDD.n7387 VDD.n7385 0.024
R13525 VDD.n7405 VDD.n7404 0.024
R13526 VDD.n7483 VDD.n7482 0.024
R13527 VDD.n7481 VDD.n7480 0.024
R13528 VDD.n7568 VDD.n7567 0.024
R13529 VDD.n7600 VDD.n7598 0.024
R13530 VDD.n7611 VDD.n7609 0.024
R13531 VDD.n7707 VDD.n7705 0.024
R13532 VDD.n7718 VDD.n7716 0.024
R13533 VDD.n7749 VDD.n7747 0.024
R13534 VDD.n7767 VDD.n7766 0.024
R13535 VDD.n7845 VDD.n7844 0.024
R13536 VDD.n7843 VDD.n7842 0.024
R13537 VDD.n7930 VDD.n7929 0.024
R13538 VDD.n7962 VDD.n7960 0.024
R13539 VDD.n7973 VDD.n7971 0.024
R13540 VDD.n8069 VDD.n8067 0.024
R13541 VDD.n8080 VDD.n8078 0.024
R13542 VDD.n8111 VDD.n8109 0.024
R13543 VDD.n8129 VDD.n8128 0.024
R13544 VDD.n8207 VDD.n8206 0.024
R13545 VDD.n8205 VDD.n8204 0.024
R13546 VDD.n8292 VDD.n8291 0.024
R13547 VDD.n8324 VDD.n8322 0.024
R13548 VDD.n8335 VDD.n8333 0.024
R13549 VDD.n8431 VDD.n8429 0.024
R13550 VDD.n8442 VDD.n8440 0.024
R13551 VDD.n8473 VDD.n8471 0.024
R13552 VDD.n8491 VDD.n8490 0.024
R13553 VDD.n8569 VDD.n8568 0.024
R13554 VDD.n8567 VDD.n8566 0.024
R13555 VDD.n8654 VDD.n8653 0.024
R13556 VDD.n8686 VDD.n8684 0.024
R13557 VDD.n8697 VDD.n8695 0.024
R13558 VDD.n8793 VDD.n8791 0.024
R13559 VDD.n8804 VDD.n8802 0.024
R13560 VDD.n8835 VDD.n8833 0.024
R13561 VDD.n8853 VDD.n8852 0.024
R13562 VDD.n8931 VDD.n8930 0.024
R13563 VDD.n8929 VDD.n8928 0.024
R13564 VDD.n9016 VDD.n9015 0.024
R13565 VDD.n9048 VDD.n9046 0.024
R13566 VDD.n9059 VDD.n9057 0.024
R13567 VDD.n9155 VDD.n9153 0.024
R13568 VDD.n9166 VDD.n9164 0.024
R13569 VDD.n9197 VDD.n9195 0.024
R13570 VDD.n9215 VDD.n9214 0.024
R13571 VDD.n9293 VDD.n9292 0.024
R13572 VDD.n9291 VDD.n9290 0.024
R13573 VDD.n9378 VDD.n9377 0.024
R13574 VDD.n9410 VDD.n9408 0.024
R13575 VDD.n9421 VDD.n9419 0.024
R13576 VDD.n9517 VDD.n9515 0.024
R13577 VDD.n9528 VDD.n9526 0.024
R13578 VDD.n9559 VDD.n9557 0.024
R13579 VDD.n9577 VDD.n9576 0.024
R13580 VDD.n9655 VDD.n9654 0.024
R13581 VDD.n9653 VDD.n9652 0.024
R13582 VDD.n9740 VDD.n9739 0.024
R13583 VDD.n9772 VDD.n9770 0.024
R13584 VDD.n9783 VDD.n9781 0.024
R13585 VDD.n9879 VDD.n9877 0.024
R13586 VDD.n9890 VDD.n9888 0.024
R13587 VDD.n9921 VDD.n9919 0.024
R13588 VDD.n9939 VDD.n9938 0.024
R13589 VDD.n10437 VDD.n10434 0.024
R13590 VDD.n10442 VDD.n10440 0.024
R13591 VDD.n10424 VDD.n10423 0.024
R13592 VDD.n10431 VDD.n10428 0.024
R13593 VDD.n10401 VDD.n10400 0.024
R13594 VDD.n10416 VDD.n10414 0.024
R13595 VDD.n10411 VDD.n10410 0.024
R13596 VDD.n10374 VDD.n10373 0.024
R13597 VDD.n10389 VDD.n10387 0.024
R13598 VDD.n10384 VDD.n10383 0.024
R13599 VDD.n10357 VDD.n10356 0.024
R13600 VDD.n10362 VDD.n10360 0.024
R13601 VDD.n10343 VDD.n10342 0.024
R13602 VDD.n10349 VDD.n10346 0.024
R13603 VDD.n12304 VDD.n12302 0.024
R13604 VDD.n12283 VDD.n12281 0.024
R13605 VDD.n4578 VDD.n4577 0.023
R13606 VDD.n4596 VDD.n4595 0.023
R13607 VDD.n2935 VDD.n2934 0.023
R13608 VDD.n353 VDD.n352 0.023
R13609 VDD.n1972 VDD.n1971 0.023
R13610 VDD.n1990 VDD.n1989 0.023
R13611 VDD.n2705 VDD.n2704 0.023
R13612 VDD.n2498 VDD.n2497 0.022
R13613 VDD.n2520 VDD.n2519 0.022
R13614 VDD.n2575 VDD.n2574 0.022
R13615 VDD.n5170 VDD.n5169 0.022
R13616 VDD.n5189 VDD.n5188 0.022
R13617 VDD.n5255 VDD.n5254 0.022
R13618 VDD.n2753 VDD.n2752 0.022
R13619 VDD.n5105 VDD.n5104 0.022
R13620 VDD.n192 VDD.n191 0.022
R13621 VDD.n111 VDD.n110 0.022
R13622 VDD.n104 VDD.n103 0.022
R13623 VDD.n2604 VDD.n2603 0.022
R13624 VDD.n2706 VDD.n2705 0.022
R13625 VDD.n2757 VDD.n2756 0.022
R13626 VDD.n5140 VDD.n5139 0.022
R13627 VDD.n5472 VDD.n5471 0.022
R13628 VDD.n5478 VDD.n5477 0.022
R13629 VDD.n5432 VDD.n5431 0.022
R13630 VDD.n5590 VDD.n5588 0.022
R13631 VDD.n5597 VDD.n5596 0.022
R13632 VDD.n5833 VDD.n5832 0.022
R13633 VDD.n5839 VDD.n5838 0.022
R13634 VDD.n5793 VDD.n5792 0.022
R13635 VDD.n5951 VDD.n5949 0.022
R13636 VDD.n5958 VDD.n5957 0.022
R13637 VDD.n6195 VDD.n6194 0.022
R13638 VDD.n6201 VDD.n6200 0.022
R13639 VDD.n6155 VDD.n6154 0.022
R13640 VDD.n6313 VDD.n6311 0.022
R13641 VDD.n6320 VDD.n6319 0.022
R13642 VDD.n6557 VDD.n6556 0.022
R13643 VDD.n6563 VDD.n6562 0.022
R13644 VDD.n6517 VDD.n6516 0.022
R13645 VDD.n6675 VDD.n6673 0.022
R13646 VDD.n6682 VDD.n6681 0.022
R13647 VDD.n6919 VDD.n6918 0.022
R13648 VDD.n6925 VDD.n6924 0.022
R13649 VDD.n6879 VDD.n6878 0.022
R13650 VDD.n7037 VDD.n7035 0.022
R13651 VDD.n7044 VDD.n7043 0.022
R13652 VDD.n7281 VDD.n7280 0.022
R13653 VDD.n7287 VDD.n7286 0.022
R13654 VDD.n7241 VDD.n7240 0.022
R13655 VDD.n7399 VDD.n7397 0.022
R13656 VDD.n7406 VDD.n7405 0.022
R13657 VDD.n7643 VDD.n7642 0.022
R13658 VDD.n7649 VDD.n7648 0.022
R13659 VDD.n7603 VDD.n7602 0.022
R13660 VDD.n7761 VDD.n7759 0.022
R13661 VDD.n7768 VDD.n7767 0.022
R13662 VDD.n8005 VDD.n8004 0.022
R13663 VDD.n8011 VDD.n8010 0.022
R13664 VDD.n7965 VDD.n7964 0.022
R13665 VDD.n8123 VDD.n8121 0.022
R13666 VDD.n8130 VDD.n8129 0.022
R13667 VDD.n8367 VDD.n8366 0.022
R13668 VDD.n8373 VDD.n8372 0.022
R13669 VDD.n8327 VDD.n8326 0.022
R13670 VDD.n8485 VDD.n8483 0.022
R13671 VDD.n8492 VDD.n8491 0.022
R13672 VDD.n8729 VDD.n8728 0.022
R13673 VDD.n8735 VDD.n8734 0.022
R13674 VDD.n8689 VDD.n8688 0.022
R13675 VDD.n8847 VDD.n8845 0.022
R13676 VDD.n8854 VDD.n8853 0.022
R13677 VDD.n9091 VDD.n9090 0.022
R13678 VDD.n9097 VDD.n9096 0.022
R13679 VDD.n9051 VDD.n9050 0.022
R13680 VDD.n9209 VDD.n9207 0.022
R13681 VDD.n9216 VDD.n9215 0.022
R13682 VDD.n9453 VDD.n9452 0.022
R13683 VDD.n9459 VDD.n9458 0.022
R13684 VDD.n9413 VDD.n9412 0.022
R13685 VDD.n9571 VDD.n9569 0.022
R13686 VDD.n9578 VDD.n9577 0.022
R13687 VDD.n9815 VDD.n9814 0.022
R13688 VDD.n9821 VDD.n9820 0.022
R13689 VDD.n9775 VDD.n9774 0.022
R13690 VDD.n9933 VDD.n9931 0.022
R13691 VDD.n9940 VDD.n9939 0.022
R13692 VDD.n11574 VDD.n11573 0.022
R13693 VDD.n11732 VDD.n11731 0.022
R13694 VDD.n10804 VDD.n10803 0.022
R13695 VDD.n10963 VDD.n10962 0.022
R13696 VDD.n10945 VDD.n10944 0.022
R13697 VDD.n11075 VDD.n11074 0.022
R13698 VDD.n10860 VDD.n10859 0.022
R13699 VDD.n10844 VDD.n10843 0.022
R13700 VDD.n10723 VDD.n10722 0.022
R13701 VDD.n11702 VDD.n11701 0.022
R13702 VDD.n11843 VDD.n11842 0.022
R13703 VDD.n11641 VDD.n11640 0.022
R13704 VDD.n11623 VDD.n11622 0.022
R13705 VDD.n11493 VDD.n11492 0.022
R13706 VDD.n2627 VDD.n2626 0.021
R13707 VDD.n86 VDD.n84 0.021
R13708 VDD.n39 VDD.n37 0.021
R13709 VDD.n5059 VDD.n5057 0.021
R13710 VDD.n4940 VDD.n4938 0.021
R13711 VDD.n4828 VDD.n4826 0.021
R13712 VDD.n4709 VDD.n4707 0.021
R13713 VDD.n4573 VDD.n4572 0.021
R13714 VDD.n4575 VDD.n4574 0.021
R13715 VDD.n4593 VDD.n4592 0.021
R13716 VDD.n2820 VDD.n2819 0.021
R13717 VDD.n2822 VDD.n2821 0.021
R13718 VDD.n2915 VDD.n2898 0.021
R13719 VDD.n3071 VDD.n3070 0.021
R13720 VDD.n3186 VDD.n3174 0.021
R13721 VDD.n3308 VDD.n3307 0.021
R13722 VDD.n3423 VDD.n3411 0.021
R13723 VDD.n3546 VDD.n3545 0.021
R13724 VDD.n3661 VDD.n3649 0.021
R13725 VDD.n3783 VDD.n3782 0.021
R13726 VDD.n3898 VDD.n3886 0.021
R13727 VDD.n4021 VDD.n4020 0.021
R13728 VDD.n4136 VDD.n4124 0.021
R13729 VDD.n4258 VDD.n4257 0.021
R13730 VDD.n4373 VDD.n4361 0.021
R13731 VDD.n4513 VDD.n4512 0.021
R13732 VDD.n244 VDD.n243 0.021
R13733 VDD.n246 VDD.n245 0.021
R13734 VDD.n289 VDD.n288 0.021
R13735 VDD.n1967 VDD.n1966 0.021
R13736 VDD.n1969 VDD.n1968 0.021
R13737 VDD.n1987 VDD.n1986 0.021
R13738 VDD.n328 VDD.n312 0.021
R13739 VDD.n491 VDD.n490 0.021
R13740 VDD.n599 VDD.n587 0.021
R13741 VDD.n724 VDD.n723 0.021
R13742 VDD.n832 VDD.n820 0.021
R13743 VDD.n958 VDD.n957 0.021
R13744 VDD.n1066 VDD.n1054 0.021
R13745 VDD.n1191 VDD.n1190 0.021
R13746 VDD.n1299 VDD.n1287 0.021
R13747 VDD.n1425 VDD.n1424 0.021
R13748 VDD.n1533 VDD.n1521 0.021
R13749 VDD.n1658 VDD.n1657 0.021
R13750 VDD.n1766 VDD.n1754 0.021
R13751 VDD.n1905 VDD.n1904 0.021
R13752 VDD.n2105 VDD.n2103 0.021
R13753 VDD.n2224 VDD.n2222 0.021
R13754 VDD.n2336 VDD.n2334 0.021
R13755 VDD.n2455 VDD.n2453 0.021
R13756 VDD.n12317 VDD.n12315 0.021
R13757 VDD.n12270 VDD.n12268 0.021
R13758 VDD.n2535 VDD.n2534 0.021
R13759 VDD.n2501 VDD.n2500 0.02
R13760 VDD.n2543 VDD.n2542 0.02
R13761 VDD.n2589 VDD.n2543 0.02
R13762 VDD.n133 VDD.n132 0.02
R13763 VDD.n5184 VDD.n5171 0.02
R13764 VDD.n5190 VDD.n5189 0.02
R13765 VDD.n5211 VDD.n5210 0.02
R13766 VDD.n5290 VDD.n5289 0.02
R13767 VDD.n5276 VDD.n5275 0.02
R13768 VDD.n5254 VDD.n5253 0.02
R13769 VDD.n2672 VDD.n2671 0.02
R13770 VDD.n2742 VDD.n2741 0.02
R13771 VDD.n2754 VDD.n2753 0.02
R13772 VDD.n5124 VDD.n5123 0.02
R13773 VDD.n5102 VDD.n5101 0.02
R13774 VDD.n188 VDD.n187 0.02
R13775 VDD.n189 VDD.n188 0.02
R13776 VDD.n2592 VDD.n2591 0.02
R13777 VDD.n2591 VDD.n2590 0.02
R13778 VDD.n168 VDD.n167 0.02
R13779 VDD.n162 VDD.n161 0.02
R13780 VDD.n160 VDD.n159 0.02
R13781 VDD.n112 VDD.n111 0.02
R13782 VDD.n105 VDD.n104 0.02
R13783 VDD.n98 VDD.n97 0.02
R13784 VDD.n5303 VDD.n5302 0.02
R13785 VDD.n2603 VDD.n2602 0.02
R13786 VDD.n2618 VDD.n2617 0.02
R13787 VDD.n2620 VDD.n2619 0.02
R13788 VDD.n2625 VDD.n2624 0.02
R13789 VDD.n2624 VDD.n2623 0.02
R13790 VDD.n2707 VDD.n2706 0.02
R13791 VDD.n2756 VDD.n2755 0.02
R13792 VDD.n5132 VDD.n5131 0.02
R13793 VDD.n5141 VDD.n5140 0.02
R13794 VDD.n5341 VDD.n5340 0.02
R13795 VDD.n5521 VDD.n5520 0.02
R13796 VDD.n5609 VDD.n5608 0.02
R13797 VDD.n5317 VDD.n5316 0.02
R13798 VDD.n5390 VDD.n5389 0.02
R13799 VDD.n5598 VDD.n5597 0.02
R13800 VDD.n5702 VDD.n5701 0.02
R13801 VDD.n5882 VDD.n5881 0.02
R13802 VDD.n5970 VDD.n5969 0.02
R13803 VDD.n5678 VDD.n5677 0.02
R13804 VDD.n5751 VDD.n5750 0.02
R13805 VDD.n5959 VDD.n5958 0.02
R13806 VDD.n6064 VDD.n6063 0.02
R13807 VDD.n6244 VDD.n6243 0.02
R13808 VDD.n6332 VDD.n6331 0.02
R13809 VDD.n6040 VDD.n6039 0.02
R13810 VDD.n6113 VDD.n6112 0.02
R13811 VDD.n6321 VDD.n6320 0.02
R13812 VDD.n6426 VDD.n6425 0.02
R13813 VDD.n6606 VDD.n6605 0.02
R13814 VDD.n6694 VDD.n6693 0.02
R13815 VDD.n6402 VDD.n6401 0.02
R13816 VDD.n6475 VDD.n6474 0.02
R13817 VDD.n6683 VDD.n6682 0.02
R13818 VDD.n6788 VDD.n6787 0.02
R13819 VDD.n6968 VDD.n6967 0.02
R13820 VDD.n7056 VDD.n7055 0.02
R13821 VDD.n6764 VDD.n6763 0.02
R13822 VDD.n6837 VDD.n6836 0.02
R13823 VDD.n7045 VDD.n7044 0.02
R13824 VDD.n7150 VDD.n7149 0.02
R13825 VDD.n7330 VDD.n7329 0.02
R13826 VDD.n7418 VDD.n7417 0.02
R13827 VDD.n7126 VDD.n7125 0.02
R13828 VDD.n7199 VDD.n7198 0.02
R13829 VDD.n7407 VDD.n7406 0.02
R13830 VDD.n7512 VDD.n7511 0.02
R13831 VDD.n7692 VDD.n7691 0.02
R13832 VDD.n7780 VDD.n7779 0.02
R13833 VDD.n7488 VDD.n7487 0.02
R13834 VDD.n7561 VDD.n7560 0.02
R13835 VDD.n7769 VDD.n7768 0.02
R13836 VDD.n7874 VDD.n7873 0.02
R13837 VDD.n8054 VDD.n8053 0.02
R13838 VDD.n8142 VDD.n8141 0.02
R13839 VDD.n7850 VDD.n7849 0.02
R13840 VDD.n7923 VDD.n7922 0.02
R13841 VDD.n8131 VDD.n8130 0.02
R13842 VDD.n8236 VDD.n8235 0.02
R13843 VDD.n8416 VDD.n8415 0.02
R13844 VDD.n8504 VDD.n8503 0.02
R13845 VDD.n8212 VDD.n8211 0.02
R13846 VDD.n8285 VDD.n8284 0.02
R13847 VDD.n8493 VDD.n8492 0.02
R13848 VDD.n8598 VDD.n8597 0.02
R13849 VDD.n8778 VDD.n8777 0.02
R13850 VDD.n8866 VDD.n8865 0.02
R13851 VDD.n8574 VDD.n8573 0.02
R13852 VDD.n8647 VDD.n8646 0.02
R13853 VDD.n8855 VDD.n8854 0.02
R13854 VDD.n8960 VDD.n8959 0.02
R13855 VDD.n9140 VDD.n9139 0.02
R13856 VDD.n9228 VDD.n9227 0.02
R13857 VDD.n8936 VDD.n8935 0.02
R13858 VDD.n9009 VDD.n9008 0.02
R13859 VDD.n9217 VDD.n9216 0.02
R13860 VDD.n9322 VDD.n9321 0.02
R13861 VDD.n9502 VDD.n9501 0.02
R13862 VDD.n9590 VDD.n9589 0.02
R13863 VDD.n9298 VDD.n9297 0.02
R13864 VDD.n9371 VDD.n9370 0.02
R13865 VDD.n9579 VDD.n9578 0.02
R13866 VDD.n9684 VDD.n9683 0.02
R13867 VDD.n9864 VDD.n9863 0.02
R13868 VDD.n9952 VDD.n9951 0.02
R13869 VDD.n9660 VDD.n9659 0.02
R13870 VDD.n9733 VDD.n9732 0.02
R13871 VDD.n9941 VDD.n9940 0.02
R13872 VDD.n10339 VDD.n10337 0.02
R13873 VDD.n10239 VDD.n10237 0.02
R13874 VDD.n10219 VDD.n10217 0.02
R13875 VDD.n10122 VDD.n10120 0.02
R13876 VDD.n10686 VDD.n10684 0.02
R13877 VDD.n10586 VDD.n10584 0.02
R13878 VDD.n10565 VDD.n10563 0.02
R13879 VDD.n10468 VDD.n10466 0.02
R13880 VDD.n11560 VDD.n11559 0.02
R13881 VDD.n11558 VDD.n11557 0.02
R13882 VDD.n11746 VDD.n11745 0.02
R13883 VDD.n11748 VDD.n11747 0.02
R13884 VDD.n10790 VDD.n10789 0.02
R13885 VDD.n10788 VDD.n10787 0.02
R13886 VDD.n10977 VDD.n10976 0.02
R13887 VDD.n10979 VDD.n10978 0.02
R13888 VDD.n10897 VDD.n10896 0.02
R13889 VDD.n11057 VDD.n11056 0.02
R13890 VDD.n11012 VDD.n11011 0.02
R13891 VDD.n11104 VDD.n11103 0.02
R13892 VDD.n10748 VDD.n10747 0.02
R13893 VDD.n11666 VDD.n11665 0.02
R13894 VDD.n11823 VDD.n11822 0.02
R13895 VDD.n11780 VDD.n11779 0.02
R13896 VDD.n11878 VDD.n11877 0.02
R13897 VDD.n11519 VDD.n11518 0.02
R13898 VDD.n90 VDD.n22 0.02
R13899 VDD.n12321 VDD.n12253 0.02
R13900 VDD.n12253 VDD.n12252 0.02
R13901 VDD.n173 VDD.n169 0.02
R13902 VDD.n2692 VDD.n2621 0.02
R13903 VDD.n5069 VDD.n5059 0.019
R13904 VDD.n4938 VDD.n4936 0.019
R13905 VDD.n4838 VDD.n4828 0.019
R13906 VDD.n4707 VDD.n4705 0.019
R13907 VDD.n4610 VDD.n4609 0.019
R13908 VDD.n4584 VDD.n4583 0.019
R13909 VDD.n4589 VDD.n4588 0.019
R13910 VDD.n4598 VDD.n4597 0.019
R13911 VDD.n2945 VDD.n2944 0.019
R13912 VDD.n2872 VDD.n2871 0.019
R13913 VDD.n2878 VDD.n2877 0.019
R13914 VDD.n2937 VDD.n2936 0.019
R13915 VDD.n2898 VDD.n2897 0.019
R13916 VDD.n3072 VDD.n3071 0.019
R13917 VDD.n3174 VDD.n3173 0.019
R13918 VDD.n3309 VDD.n3308 0.019
R13919 VDD.n3411 VDD.n3410 0.019
R13920 VDD.n3547 VDD.n3546 0.019
R13921 VDD.n3649 VDD.n3648 0.019
R13922 VDD.n3784 VDD.n3783 0.019
R13923 VDD.n3886 VDD.n3885 0.019
R13924 VDD.n4022 VDD.n4021 0.019
R13925 VDD.n4124 VDD.n4123 0.019
R13926 VDD.n4259 VDD.n4258 0.019
R13927 VDD.n4361 VDD.n4360 0.019
R13928 VDD.n4514 VDD.n4513 0.019
R13929 VDD.n362 VDD.n361 0.019
R13930 VDD.n286 VDD.n285 0.019
R13931 VDD.n293 VDD.n292 0.019
R13932 VDD.n355 VDD.n354 0.019
R13933 VDD.n2004 VDD.n2003 0.019
R13934 VDD.n1978 VDD.n1977 0.019
R13935 VDD.n1983 VDD.n1982 0.019
R13936 VDD.n1992 VDD.n1991 0.019
R13937 VDD.n312 VDD.n311 0.019
R13938 VDD.n492 VDD.n491 0.019
R13939 VDD.n587 VDD.n586 0.019
R13940 VDD.n725 VDD.n724 0.019
R13941 VDD.n820 VDD.n819 0.019
R13942 VDD.n959 VDD.n958 0.019
R13943 VDD.n1054 VDD.n1053 0.019
R13944 VDD.n1192 VDD.n1191 0.019
R13945 VDD.n1287 VDD.n1286 0.019
R13946 VDD.n1426 VDD.n1425 0.019
R13947 VDD.n1521 VDD.n1520 0.019
R13948 VDD.n1659 VDD.n1658 0.019
R13949 VDD.n1754 VDD.n1753 0.019
R13950 VDD.n1906 VDD.n1905 0.019
R13951 VDD.n2103 VDD.n2101 0.019
R13952 VDD.n2234 VDD.n2224 0.019
R13953 VDD.n2334 VDD.n2332 0.019
R13954 VDD.n2465 VDD.n2455 0.019
R13955 VDD.n2518 VDD.n2517 0.018
R13956 VDD.n2542 VDD.n2539 0.018
R13957 VDD.n2571 VDD.n2570 0.018
R13958 VDD.n2567 VDD.n2566 0.018
R13959 VDD.n5225 VDD.n5224 0.018
R13960 VDD.n5232 VDD.n5226 0.018
R13961 VDD.n5249 VDD.n5236 0.018
R13962 VDD.n2670 VDD.n2669 0.018
R13963 VDD.n2655 VDD.n2654 0.018
R13964 VDD.n2731 VDD.n2730 0.018
R13965 VDD.n2747 VDD.n2743 0.018
R13966 VDD.n2537 VDD.n2536 0.018
R13967 VDD.n167 VDD.n166 0.018
R13968 VDD.n2611 VDD.n2610 0.018
R13969 VDD.n2616 VDD.n2615 0.018
R13970 VDD.n10337 VDD.n10335 0.018
R13971 VDD.n10247 VDD.n10239 0.018
R13972 VDD.n10217 VDD.n10215 0.018
R13973 VDD.n10131 VDD.n10122 0.018
R13974 VDD.n10684 VDD.n10682 0.018
R13975 VDD.n10594 VDD.n10586 0.018
R13976 VDD.n10563 VDD.n10561 0.018
R13977 VDD.n10477 VDD.n10468 0.018
R13978 VDD.n11572 VDD.n11571 0.018
R13979 VDD.n11734 VDD.n11733 0.018
R13980 VDD.n10802 VDD.n10801 0.018
R13981 VDD.n10965 VDD.n10964 0.018
R13982 VDD.n10894 VDD.n10892 0.018
R13983 VDD.n10954 VDD.n10953 0.018
R13984 VDD.n10935 VDD.n10934 0.018
R13985 VDD.n10733 VDD.n10732 0.018
R13986 VDD.n10770 VDD.n10769 0.018
R13987 VDD.n10720 VDD.n10718 0.018
R13988 VDD.n11663 VDD.n11661 0.018
R13989 VDD.n11723 VDD.n11722 0.018
R13990 VDD.n11690 VDD.n11688 0.018
R13991 VDD.n11504 VDD.n11503 0.018
R13992 VDD.n11540 VDD.n11539 0.018
R13993 VDD.n11490 VDD.n11488 0.018
R13994 VDD.n2614 VDD.n2613 0.018
R13995 VDD.n4582 VDD.n4581 0.017
R13996 VDD.n4587 VDD.n4586 0.017
R13997 VDD.n2849 VDD.n2848 0.017
R13998 VDD.n2880 VDD.n2879 0.017
R13999 VDD.n295 VDD.n294 0.017
R14000 VDD.n1976 VDD.n1975 0.017
R14001 VDD.n1981 VDD.n1980 0.017
R14002 VDD.n2526 VDD.n2525 0.017
R14003 VDD.n2587 VDD.n2576 0.017
R14004 VDD.n2564 VDD.n2563 0.017
R14005 VDD.n2548 VDD.n2547 0.017
R14006 VDD.n2546 VDD.n2545 0.017
R14007 VDD.n131 VDD.n130 0.017
R14008 VDD.n5168 VDD.n5167 0.017
R14009 VDD.n5205 VDD.n5192 0.017
R14010 VDD.n5207 VDD.n5206 0.017
R14011 VDD.n5294 VDD.n5291 0.017
R14012 VDD.n5271 VDD.n5270 0.017
R14013 VDD.n2649 VDD.n2648 0.017
R14014 VDD.n2727 VDD.n2726 0.017
R14015 VDD.n2752 VDD.n2749 0.017
R14016 VDD.n2759 VDD.n2758 0.017
R14017 VDD.n5122 VDD.n5121 0.017
R14018 VDD.n175 VDD.n174 0.017
R14019 VDD.n115 VDD.n114 0.017
R14020 VDD.n2621 VDD.n2620 0.017
R14021 VDD.n5350 VDD.n5349 0.017
R14022 VDD.n5624 VDD.n5623 0.017
R14023 VDD.n5648 VDD.n5644 0.017
R14024 VDD.n5554 VDD.n5553 0.017
R14025 VDD.n5578 VDD.n5577 0.017
R14026 VDD.n5711 VDD.n5710 0.017
R14027 VDD.n5985 VDD.n5984 0.017
R14028 VDD.n6009 VDD.n6005 0.017
R14029 VDD.n5915 VDD.n5914 0.017
R14030 VDD.n5939 VDD.n5938 0.017
R14031 VDD.n6073 VDD.n6072 0.017
R14032 VDD.n6347 VDD.n6346 0.017
R14033 VDD.n6371 VDD.n6367 0.017
R14034 VDD.n6277 VDD.n6276 0.017
R14035 VDD.n6301 VDD.n6300 0.017
R14036 VDD.n6435 VDD.n6434 0.017
R14037 VDD.n6709 VDD.n6708 0.017
R14038 VDD.n6733 VDD.n6729 0.017
R14039 VDD.n6639 VDD.n6638 0.017
R14040 VDD.n6663 VDD.n6662 0.017
R14041 VDD.n6797 VDD.n6796 0.017
R14042 VDD.n7071 VDD.n7070 0.017
R14043 VDD.n7095 VDD.n7091 0.017
R14044 VDD.n7001 VDD.n7000 0.017
R14045 VDD.n7025 VDD.n7024 0.017
R14046 VDD.n7159 VDD.n7158 0.017
R14047 VDD.n7433 VDD.n7432 0.017
R14048 VDD.n7457 VDD.n7453 0.017
R14049 VDD.n7363 VDD.n7362 0.017
R14050 VDD.n7387 VDD.n7386 0.017
R14051 VDD.n7521 VDD.n7520 0.017
R14052 VDD.n7795 VDD.n7794 0.017
R14053 VDD.n7819 VDD.n7815 0.017
R14054 VDD.n7725 VDD.n7724 0.017
R14055 VDD.n7749 VDD.n7748 0.017
R14056 VDD.n7883 VDD.n7882 0.017
R14057 VDD.n8157 VDD.n8156 0.017
R14058 VDD.n8181 VDD.n8177 0.017
R14059 VDD.n8087 VDD.n8086 0.017
R14060 VDD.n8111 VDD.n8110 0.017
R14061 VDD.n8245 VDD.n8244 0.017
R14062 VDD.n8519 VDD.n8518 0.017
R14063 VDD.n8543 VDD.n8539 0.017
R14064 VDD.n8449 VDD.n8448 0.017
R14065 VDD.n8473 VDD.n8472 0.017
R14066 VDD.n8607 VDD.n8606 0.017
R14067 VDD.n8881 VDD.n8880 0.017
R14068 VDD.n8905 VDD.n8901 0.017
R14069 VDD.n8811 VDD.n8810 0.017
R14070 VDD.n8835 VDD.n8834 0.017
R14071 VDD.n8969 VDD.n8968 0.017
R14072 VDD.n9243 VDD.n9242 0.017
R14073 VDD.n9267 VDD.n9263 0.017
R14074 VDD.n9173 VDD.n9172 0.017
R14075 VDD.n9197 VDD.n9196 0.017
R14076 VDD.n9331 VDD.n9330 0.017
R14077 VDD.n9605 VDD.n9604 0.017
R14078 VDD.n9629 VDD.n9625 0.017
R14079 VDD.n9535 VDD.n9534 0.017
R14080 VDD.n9559 VDD.n9558 0.017
R14081 VDD.n9693 VDD.n9692 0.017
R14082 VDD.n9967 VDD.n9966 0.017
R14083 VDD.n9991 VDD.n9987 0.017
R14084 VDD.n9897 VDD.n9896 0.017
R14085 VDD.n9921 VDD.n9920 0.017
R14086 VDD.n10688 VDD.n10567 0.017
R14087 VDD.n5045 VDD.n5043 0.016
R14088 VDD.n4954 VDD.n4952 0.016
R14089 VDD.n4814 VDD.n4812 0.016
R14090 VDD.n4723 VDD.n4721 0.016
R14091 VDD.n4603 VDD.n4602 0.016
R14092 VDD.n2962 VDD.n2917 0.016
R14093 VDD.n3057 VDD.n3056 0.016
R14094 VDD.n3200 VDD.n3188 0.016
R14095 VDD.n3294 VDD.n3293 0.016
R14096 VDD.n3437 VDD.n3425 0.016
R14097 VDD.n3532 VDD.n3531 0.016
R14098 VDD.n3675 VDD.n3663 0.016
R14099 VDD.n3769 VDD.n3768 0.016
R14100 VDD.n3912 VDD.n3900 0.016
R14101 VDD.n4007 VDD.n4006 0.016
R14102 VDD.n4150 VDD.n4138 0.016
R14103 VDD.n4244 VDD.n4243 0.016
R14104 VDD.n4387 VDD.n4375 0.016
R14105 VDD.n4493 VDD.n4492 0.016
R14106 VDD.n237 VDD.n236 0.016
R14107 VDD.n1997 VDD.n1996 0.016
R14108 VDD.n379 VDD.n330 0.016
R14109 VDD.n477 VDD.n476 0.016
R14110 VDD.n613 VDD.n601 0.016
R14111 VDD.n710 VDD.n709 0.016
R14112 VDD.n846 VDD.n834 0.016
R14113 VDD.n944 VDD.n943 0.016
R14114 VDD.n1080 VDD.n1068 0.016
R14115 VDD.n1177 VDD.n1176 0.016
R14116 VDD.n1313 VDD.n1301 0.016
R14117 VDD.n1411 VDD.n1410 0.016
R14118 VDD.n1547 VDD.n1535 0.016
R14119 VDD.n1644 VDD.n1643 0.016
R14120 VDD.n1780 VDD.n1768 0.016
R14121 VDD.n1886 VDD.n1885 0.016
R14122 VDD.n2119 VDD.n2117 0.016
R14123 VDD.n2210 VDD.n2208 0.016
R14124 VDD.n2350 VDD.n2348 0.016
R14125 VDD.n2441 VDD.n2439 0.016
R14126 VDD.n5400 VDD.n5399 0.016
R14127 VDD.n5417 VDD.n5416 0.016
R14128 VDD.n5443 VDD.n5442 0.016
R14129 VDD.n5462 VDD.n5461 0.016
R14130 VDD.n5550 VDD.n5549 0.016
R14131 VDD.n5566 VDD.n5565 0.016
R14132 VDD.n5593 VDD.n5592 0.016
R14133 VDD.n5761 VDD.n5760 0.016
R14134 VDD.n5778 VDD.n5777 0.016
R14135 VDD.n5804 VDD.n5803 0.016
R14136 VDD.n5823 VDD.n5822 0.016
R14137 VDD.n5911 VDD.n5910 0.016
R14138 VDD.n5927 VDD.n5926 0.016
R14139 VDD.n5954 VDD.n5953 0.016
R14140 VDD.n6123 VDD.n6122 0.016
R14141 VDD.n6140 VDD.n6139 0.016
R14142 VDD.n6166 VDD.n6165 0.016
R14143 VDD.n6185 VDD.n6184 0.016
R14144 VDD.n6273 VDD.n6272 0.016
R14145 VDD.n6289 VDD.n6288 0.016
R14146 VDD.n6316 VDD.n6315 0.016
R14147 VDD.n6485 VDD.n6484 0.016
R14148 VDD.n6502 VDD.n6501 0.016
R14149 VDD.n6528 VDD.n6527 0.016
R14150 VDD.n6547 VDD.n6546 0.016
R14151 VDD.n6635 VDD.n6634 0.016
R14152 VDD.n6651 VDD.n6650 0.016
R14153 VDD.n6678 VDD.n6677 0.016
R14154 VDD.n6847 VDD.n6846 0.016
R14155 VDD.n6864 VDD.n6863 0.016
R14156 VDD.n6890 VDD.n6889 0.016
R14157 VDD.n6909 VDD.n6908 0.016
R14158 VDD.n6997 VDD.n6996 0.016
R14159 VDD.n7013 VDD.n7012 0.016
R14160 VDD.n7040 VDD.n7039 0.016
R14161 VDD.n7209 VDD.n7208 0.016
R14162 VDD.n7226 VDD.n7225 0.016
R14163 VDD.n7252 VDD.n7251 0.016
R14164 VDD.n7271 VDD.n7270 0.016
R14165 VDD.n7359 VDD.n7358 0.016
R14166 VDD.n7375 VDD.n7374 0.016
R14167 VDD.n7402 VDD.n7401 0.016
R14168 VDD.n7571 VDD.n7570 0.016
R14169 VDD.n7588 VDD.n7587 0.016
R14170 VDD.n7614 VDD.n7613 0.016
R14171 VDD.n7633 VDD.n7632 0.016
R14172 VDD.n7721 VDD.n7720 0.016
R14173 VDD.n7737 VDD.n7736 0.016
R14174 VDD.n7764 VDD.n7763 0.016
R14175 VDD.n7933 VDD.n7932 0.016
R14176 VDD.n7950 VDD.n7949 0.016
R14177 VDD.n7976 VDD.n7975 0.016
R14178 VDD.n7995 VDD.n7994 0.016
R14179 VDD.n8083 VDD.n8082 0.016
R14180 VDD.n8099 VDD.n8098 0.016
R14181 VDD.n8126 VDD.n8125 0.016
R14182 VDD.n8295 VDD.n8294 0.016
R14183 VDD.n8312 VDD.n8311 0.016
R14184 VDD.n8338 VDD.n8337 0.016
R14185 VDD.n8357 VDD.n8356 0.016
R14186 VDD.n8445 VDD.n8444 0.016
R14187 VDD.n8461 VDD.n8460 0.016
R14188 VDD.n8488 VDD.n8487 0.016
R14189 VDD.n8657 VDD.n8656 0.016
R14190 VDD.n8674 VDD.n8673 0.016
R14191 VDD.n8700 VDD.n8699 0.016
R14192 VDD.n8719 VDD.n8718 0.016
R14193 VDD.n8807 VDD.n8806 0.016
R14194 VDD.n8823 VDD.n8822 0.016
R14195 VDD.n8850 VDD.n8849 0.016
R14196 VDD.n9019 VDD.n9018 0.016
R14197 VDD.n9036 VDD.n9035 0.016
R14198 VDD.n9062 VDD.n9061 0.016
R14199 VDD.n9081 VDD.n9080 0.016
R14200 VDD.n9169 VDD.n9168 0.016
R14201 VDD.n9185 VDD.n9184 0.016
R14202 VDD.n9212 VDD.n9211 0.016
R14203 VDD.n9381 VDD.n9380 0.016
R14204 VDD.n9398 VDD.n9397 0.016
R14205 VDD.n9424 VDD.n9423 0.016
R14206 VDD.n9443 VDD.n9442 0.016
R14207 VDD.n9531 VDD.n9530 0.016
R14208 VDD.n9547 VDD.n9546 0.016
R14209 VDD.n9574 VDD.n9573 0.016
R14210 VDD.n9743 VDD.n9742 0.016
R14211 VDD.n9760 VDD.n9759 0.016
R14212 VDD.n9786 VDD.n9785 0.016
R14213 VDD.n9805 VDD.n9804 0.016
R14214 VDD.n9893 VDD.n9892 0.016
R14215 VDD.n9909 VDD.n9908 0.016
R14216 VDD.n9936 VDD.n9935 0.016
R14217 VDD.n12201 VDD.n12199 0.016
R14218 VDD.n12179 VDD.n12177 0.016
R14219 VDD.n11997 VDD.n11995 0.016
R14220 VDD.n11975 VDD.n11973 0.016
R14221 VDD.n11429 VDD.n11427 0.016
R14222 VDD.n11409 VDD.n11407 0.016
R14223 VDD.n11231 VDD.n11229 0.016
R14224 VDD.n11211 VDD.n11209 0.016
R14225 VDD.n117 VDD.n116 0.016
R14226 VDD.n109 VDD.n108 0.016
R14227 VDD.n5305 VDD.n5304 0.015
R14228 VDD.n4591 VDD.n4590 0.015
R14229 VDD.n2876 VDD.n2875 0.015
R14230 VDD.n291 VDD.n290 0.015
R14231 VDD.n1985 VDD.n1984 0.015
R14232 VDD.n2496 VDD.n2483 0.015
R14233 VDD.n2588 VDD.n2587 0.015
R14234 VDD.n2569 VDD.n2568 0.015
R14235 VDD.n149 VDD.n137 0.015
R14236 VDD.n151 VDD.n150 0.015
R14237 VDD.n5206 VDD.n5205 0.015
R14238 VDD.n5209 VDD.n5208 0.015
R14239 VDD.n5275 VDD.n5274 0.015
R14240 VDD.n5272 VDD.n5271 0.015
R14241 VDD.n5270 VDD.n5257 0.015
R14242 VDD.n2632 VDD.n2631 0.015
R14243 VDD.n2688 VDD.n2676 0.015
R14244 VDD.n2653 VDD.n2652 0.015
R14245 VDD.n2723 VDD.n2710 0.015
R14246 VDD.n2724 VDD.n2723 0.015
R14247 VDD.n2726 VDD.n2725 0.015
R14248 VDD.n5125 VDD.n5124 0.015
R14249 VDD.n5121 VDD.n5120 0.015
R14250 VDD.n2538 VDD.n2537 0.015
R14251 VDD.n2532 VDD.n2531 0.015
R14252 VDD.n163 VDD.n162 0.015
R14253 VDD.n96 VDD.n95 0.015
R14254 VDD.n99 VDD.n98 0.015
R14255 VDD.n5302 VDD.n5301 0.015
R14256 VDD.n2617 VDD.n2616 0.015
R14257 VDD.n2694 VDD.n2693 0.015
R14258 VDD.n5375 VDD.n5374 0.015
R14259 VDD.n5369 VDD.n5368 0.015
R14260 VDD.n5367 VDD.n5366 0.015
R14261 VDD.n5522 VDD.n5521 0.015
R14262 VDD.n5650 VDD.n5649 0.015
R14263 VDD.n5656 VDD.n5655 0.015
R14264 VDD.n5311 VDD.n5310 0.015
R14265 VDD.n5391 VDD.n5390 0.015
R14266 VDD.n5396 VDD.n5395 0.015
R14267 VDD.n5427 VDD.n5426 0.015
R14268 VDD.n5438 VDD.n5437 0.015
R14269 VDD.n5447 VDD.n5446 0.015
R14270 VDD.n5534 VDD.n5533 0.015
R14271 VDD.n5536 VDD.n5535 0.015
R14272 VDD.n5545 VDD.n5544 0.015
R14273 VDD.n5576 VDD.n5575 0.015
R14274 VDD.n5587 VDD.n5586 0.015
R14275 VDD.n5736 VDD.n5735 0.015
R14276 VDD.n5730 VDD.n5729 0.015
R14277 VDD.n5728 VDD.n5727 0.015
R14278 VDD.n5883 VDD.n5882 0.015
R14279 VDD.n6011 VDD.n6010 0.015
R14280 VDD.n6017 VDD.n6016 0.015
R14281 VDD.n5672 VDD.n5671 0.015
R14282 VDD.n5752 VDD.n5751 0.015
R14283 VDD.n5757 VDD.n5756 0.015
R14284 VDD.n5788 VDD.n5787 0.015
R14285 VDD.n5799 VDD.n5798 0.015
R14286 VDD.n5808 VDD.n5807 0.015
R14287 VDD.n5895 VDD.n5894 0.015
R14288 VDD.n5897 VDD.n5896 0.015
R14289 VDD.n5906 VDD.n5905 0.015
R14290 VDD.n5937 VDD.n5936 0.015
R14291 VDD.n5948 VDD.n5947 0.015
R14292 VDD.n6098 VDD.n6097 0.015
R14293 VDD.n6092 VDD.n6091 0.015
R14294 VDD.n6090 VDD.n6089 0.015
R14295 VDD.n6245 VDD.n6244 0.015
R14296 VDD.n6373 VDD.n6372 0.015
R14297 VDD.n6379 VDD.n6378 0.015
R14298 VDD.n6034 VDD.n6033 0.015
R14299 VDD.n6114 VDD.n6113 0.015
R14300 VDD.n6119 VDD.n6118 0.015
R14301 VDD.n6150 VDD.n6149 0.015
R14302 VDD.n6161 VDD.n6160 0.015
R14303 VDD.n6170 VDD.n6169 0.015
R14304 VDD.n6257 VDD.n6256 0.015
R14305 VDD.n6259 VDD.n6258 0.015
R14306 VDD.n6268 VDD.n6267 0.015
R14307 VDD.n6299 VDD.n6298 0.015
R14308 VDD.n6310 VDD.n6309 0.015
R14309 VDD.n6460 VDD.n6459 0.015
R14310 VDD.n6454 VDD.n6453 0.015
R14311 VDD.n6452 VDD.n6451 0.015
R14312 VDD.n6607 VDD.n6606 0.015
R14313 VDD.n6735 VDD.n6734 0.015
R14314 VDD.n6741 VDD.n6740 0.015
R14315 VDD.n6396 VDD.n6395 0.015
R14316 VDD.n6476 VDD.n6475 0.015
R14317 VDD.n6481 VDD.n6480 0.015
R14318 VDD.n6512 VDD.n6511 0.015
R14319 VDD.n6523 VDD.n6522 0.015
R14320 VDD.n6532 VDD.n6531 0.015
R14321 VDD.n6619 VDD.n6618 0.015
R14322 VDD.n6621 VDD.n6620 0.015
R14323 VDD.n6630 VDD.n6629 0.015
R14324 VDD.n6661 VDD.n6660 0.015
R14325 VDD.n6672 VDD.n6671 0.015
R14326 VDD.n6822 VDD.n6821 0.015
R14327 VDD.n6816 VDD.n6815 0.015
R14328 VDD.n6814 VDD.n6813 0.015
R14329 VDD.n6969 VDD.n6968 0.015
R14330 VDD.n7097 VDD.n7096 0.015
R14331 VDD.n7103 VDD.n7102 0.015
R14332 VDD.n6758 VDD.n6757 0.015
R14333 VDD.n6838 VDD.n6837 0.015
R14334 VDD.n6843 VDD.n6842 0.015
R14335 VDD.n6874 VDD.n6873 0.015
R14336 VDD.n6885 VDD.n6884 0.015
R14337 VDD.n6894 VDD.n6893 0.015
R14338 VDD.n6981 VDD.n6980 0.015
R14339 VDD.n6983 VDD.n6982 0.015
R14340 VDD.n6992 VDD.n6991 0.015
R14341 VDD.n7023 VDD.n7022 0.015
R14342 VDD.n7034 VDD.n7033 0.015
R14343 VDD.n7184 VDD.n7183 0.015
R14344 VDD.n7178 VDD.n7177 0.015
R14345 VDD.n7176 VDD.n7175 0.015
R14346 VDD.n7331 VDD.n7330 0.015
R14347 VDD.n7459 VDD.n7458 0.015
R14348 VDD.n7465 VDD.n7464 0.015
R14349 VDD.n7120 VDD.n7119 0.015
R14350 VDD.n7200 VDD.n7199 0.015
R14351 VDD.n7205 VDD.n7204 0.015
R14352 VDD.n7236 VDD.n7235 0.015
R14353 VDD.n7247 VDD.n7246 0.015
R14354 VDD.n7256 VDD.n7255 0.015
R14355 VDD.n7343 VDD.n7342 0.015
R14356 VDD.n7345 VDD.n7344 0.015
R14357 VDD.n7354 VDD.n7353 0.015
R14358 VDD.n7385 VDD.n7384 0.015
R14359 VDD.n7396 VDD.n7395 0.015
R14360 VDD.n7546 VDD.n7545 0.015
R14361 VDD.n7540 VDD.n7539 0.015
R14362 VDD.n7538 VDD.n7537 0.015
R14363 VDD.n7693 VDD.n7692 0.015
R14364 VDD.n7821 VDD.n7820 0.015
R14365 VDD.n7827 VDD.n7826 0.015
R14366 VDD.n7482 VDD.n7481 0.015
R14367 VDD.n7562 VDD.n7561 0.015
R14368 VDD.n7567 VDD.n7566 0.015
R14369 VDD.n7598 VDD.n7597 0.015
R14370 VDD.n7609 VDD.n7608 0.015
R14371 VDD.n7618 VDD.n7617 0.015
R14372 VDD.n7705 VDD.n7704 0.015
R14373 VDD.n7707 VDD.n7706 0.015
R14374 VDD.n7716 VDD.n7715 0.015
R14375 VDD.n7747 VDD.n7746 0.015
R14376 VDD.n7758 VDD.n7757 0.015
R14377 VDD.n7908 VDD.n7907 0.015
R14378 VDD.n7902 VDD.n7901 0.015
R14379 VDD.n7900 VDD.n7899 0.015
R14380 VDD.n8055 VDD.n8054 0.015
R14381 VDD.n8183 VDD.n8182 0.015
R14382 VDD.n8189 VDD.n8188 0.015
R14383 VDD.n7844 VDD.n7843 0.015
R14384 VDD.n7924 VDD.n7923 0.015
R14385 VDD.n7929 VDD.n7928 0.015
R14386 VDD.n7960 VDD.n7959 0.015
R14387 VDD.n7971 VDD.n7970 0.015
R14388 VDD.n7980 VDD.n7979 0.015
R14389 VDD.n8067 VDD.n8066 0.015
R14390 VDD.n8069 VDD.n8068 0.015
R14391 VDD.n8078 VDD.n8077 0.015
R14392 VDD.n8109 VDD.n8108 0.015
R14393 VDD.n8120 VDD.n8119 0.015
R14394 VDD.n8270 VDD.n8269 0.015
R14395 VDD.n8264 VDD.n8263 0.015
R14396 VDD.n8262 VDD.n8261 0.015
R14397 VDD.n8417 VDD.n8416 0.015
R14398 VDD.n8545 VDD.n8544 0.015
R14399 VDD.n8551 VDD.n8550 0.015
R14400 VDD.n8206 VDD.n8205 0.015
R14401 VDD.n8286 VDD.n8285 0.015
R14402 VDD.n8291 VDD.n8290 0.015
R14403 VDD.n8322 VDD.n8321 0.015
R14404 VDD.n8333 VDD.n8332 0.015
R14405 VDD.n8342 VDD.n8341 0.015
R14406 VDD.n8429 VDD.n8428 0.015
R14407 VDD.n8431 VDD.n8430 0.015
R14408 VDD.n8440 VDD.n8439 0.015
R14409 VDD.n8471 VDD.n8470 0.015
R14410 VDD.n8482 VDD.n8481 0.015
R14411 VDD.n8632 VDD.n8631 0.015
R14412 VDD.n8626 VDD.n8625 0.015
R14413 VDD.n8624 VDD.n8623 0.015
R14414 VDD.n8779 VDD.n8778 0.015
R14415 VDD.n8907 VDD.n8906 0.015
R14416 VDD.n8913 VDD.n8912 0.015
R14417 VDD.n8568 VDD.n8567 0.015
R14418 VDD.n8648 VDD.n8647 0.015
R14419 VDD.n8653 VDD.n8652 0.015
R14420 VDD.n8684 VDD.n8683 0.015
R14421 VDD.n8695 VDD.n8694 0.015
R14422 VDD.n8704 VDD.n8703 0.015
R14423 VDD.n8791 VDD.n8790 0.015
R14424 VDD.n8793 VDD.n8792 0.015
R14425 VDD.n8802 VDD.n8801 0.015
R14426 VDD.n8833 VDD.n8832 0.015
R14427 VDD.n8844 VDD.n8843 0.015
R14428 VDD.n8994 VDD.n8993 0.015
R14429 VDD.n8988 VDD.n8987 0.015
R14430 VDD.n8986 VDD.n8985 0.015
R14431 VDD.n9141 VDD.n9140 0.015
R14432 VDD.n9269 VDD.n9268 0.015
R14433 VDD.n9275 VDD.n9274 0.015
R14434 VDD.n8930 VDD.n8929 0.015
R14435 VDD.n9010 VDD.n9009 0.015
R14436 VDD.n9015 VDD.n9014 0.015
R14437 VDD.n9046 VDD.n9045 0.015
R14438 VDD.n9057 VDD.n9056 0.015
R14439 VDD.n9066 VDD.n9065 0.015
R14440 VDD.n9153 VDD.n9152 0.015
R14441 VDD.n9155 VDD.n9154 0.015
R14442 VDD.n9164 VDD.n9163 0.015
R14443 VDD.n9195 VDD.n9194 0.015
R14444 VDD.n9206 VDD.n9205 0.015
R14445 VDD.n9356 VDD.n9355 0.015
R14446 VDD.n9350 VDD.n9349 0.015
R14447 VDD.n9348 VDD.n9347 0.015
R14448 VDD.n9503 VDD.n9502 0.015
R14449 VDD.n9631 VDD.n9630 0.015
R14450 VDD.n9637 VDD.n9636 0.015
R14451 VDD.n9292 VDD.n9291 0.015
R14452 VDD.n9372 VDD.n9371 0.015
R14453 VDD.n9377 VDD.n9376 0.015
R14454 VDD.n9408 VDD.n9407 0.015
R14455 VDD.n9419 VDD.n9418 0.015
R14456 VDD.n9428 VDD.n9427 0.015
R14457 VDD.n9515 VDD.n9514 0.015
R14458 VDD.n9517 VDD.n9516 0.015
R14459 VDD.n9526 VDD.n9525 0.015
R14460 VDD.n9557 VDD.n9556 0.015
R14461 VDD.n9568 VDD.n9567 0.015
R14462 VDD.n9718 VDD.n9717 0.015
R14463 VDD.n9712 VDD.n9711 0.015
R14464 VDD.n9710 VDD.n9709 0.015
R14465 VDD.n9865 VDD.n9864 0.015
R14466 VDD.n9993 VDD.n9992 0.015
R14467 VDD.n9999 VDD.n9998 0.015
R14468 VDD.n9654 VDD.n9653 0.015
R14469 VDD.n9734 VDD.n9733 0.015
R14470 VDD.n9739 VDD.n9738 0.015
R14471 VDD.n9770 VDD.n9769 0.015
R14472 VDD.n9781 VDD.n9780 0.015
R14473 VDD.n9790 VDD.n9789 0.015
R14474 VDD.n9877 VDD.n9876 0.015
R14475 VDD.n9879 VDD.n9878 0.015
R14476 VDD.n9888 VDD.n9887 0.015
R14477 VDD.n9919 VDD.n9918 0.015
R14478 VDD.n9930 VDD.n9929 0.015
R14479 VDD.n10410 VDD.n10409 0.015
R14480 VDD.n10383 VDD.n10382 0.015
R14481 VDD.n11577 VDD.n11576 0.015
R14482 VDD.n11729 VDD.n11728 0.015
R14483 VDD.n10807 VDD.n10806 0.015
R14484 VDD.n10960 VDD.n10959 0.015
R14485 VDD.n10951 VDD.n10950 0.015
R14486 VDD.n11041 VDD.n11040 0.015
R14487 VDD.n10855 VDD.n10854 0.015
R14488 VDD.n10829 VDD.n10828 0.015
R14489 VDD.n11717 VDD.n11716 0.015
R14490 VDD.n11808 VDD.n11807 0.015
R14491 VDD.n11636 VDD.n11635 0.015
R14492 VDD.n11609 VDD.n11608 0.015
R14493 VDD.n12100 VDD.n12092 0.015
R14494 VDD.n12082 VDD.n12080 0.015
R14495 VDD.n11333 VDD.n11323 0.015
R14496 VDD.n11313 VDD.n11311 0.015
R14497 VDD.n2593 VDD.n2592 0.014
R14498 VDD.n5083 VDD.n5073 0.014
R14499 VDD.n4924 VDD.n4922 0.014
R14500 VDD.n4852 VDD.n4842 0.014
R14501 VDD.n4693 VDD.n4691 0.014
R14502 VDD.n2868 VDD.n2867 0.014
R14503 VDD.n3086 VDD.n3085 0.014
R14504 VDD.n3160 VDD.n3159 0.014
R14505 VDD.n3324 VDD.n3323 0.014
R14506 VDD.n3397 VDD.n3396 0.014
R14507 VDD.n3561 VDD.n3560 0.014
R14508 VDD.n3635 VDD.n3634 0.014
R14509 VDD.n3799 VDD.n3798 0.014
R14510 VDD.n3872 VDD.n3871 0.014
R14511 VDD.n4036 VDD.n4035 0.014
R14512 VDD.n4110 VDD.n4109 0.014
R14513 VDD.n4274 VDD.n4273 0.014
R14514 VDD.n4347 VDD.n4346 0.014
R14515 VDD.n4534 VDD.n4533 0.014
R14516 VDD.n281 VDD.n280 0.014
R14517 VDD.n506 VDD.n505 0.014
R14518 VDD.n573 VDD.n572 0.014
R14519 VDD.n740 VDD.n739 0.014
R14520 VDD.n806 VDD.n805 0.014
R14521 VDD.n973 VDD.n972 0.014
R14522 VDD.n1040 VDD.n1039 0.014
R14523 VDD.n1207 VDD.n1206 0.014
R14524 VDD.n1273 VDD.n1272 0.014
R14525 VDD.n1440 VDD.n1439 0.014
R14526 VDD.n1507 VDD.n1506 0.014
R14527 VDD.n1674 VDD.n1673 0.014
R14528 VDD.n1740 VDD.n1739 0.014
R14529 VDD.n1925 VDD.n1924 0.014
R14530 VDD.n2089 VDD.n2087 0.014
R14531 VDD.n2248 VDD.n2238 0.014
R14532 VDD.n2320 VDD.n2318 0.014
R14533 VDD.n2479 VDD.n2469 0.014
R14534 VDD.n12213 VDD.n12211 0.014
R14535 VDD.n12167 VDD.n12165 0.014
R14536 VDD.n12009 VDD.n12007 0.014
R14537 VDD.n11963 VDD.n11961 0.014
R14538 VDD.n11441 VDD.n11439 0.014
R14539 VDD.n11397 VDD.n11395 0.014
R14540 VDD.n11243 VDD.n11241 0.014
R14541 VDD.n11198 VDD.n11196 0.014
R14542 VDD.n2608 VDD.n2607 0.014
R14543 VDD.n102 VDD.n99 0.014
R14544 VDD.n5129 VDD.n2757 0.014
R14545 VDD.n164 VDD.n163 0.013
R14546 VDD.n10443 VDD.n10439 0.013
R14547 VDD.n10417 VDD.n10413 0.013
R14548 VDD.n10413 VDD.n10412 0.013
R14549 VDD.n10390 VDD.n10386 0.013
R14550 VDD.n10386 VDD.n10385 0.013
R14551 VDD.n10363 VDD.n10359 0.013
R14552 VDD.n4580 VDD.n4579 0.013
R14553 VDD.n4615 VDD.n4598 0.013
R14554 VDD.n2847 VDD.n2846 0.013
R14555 VDD.n2950 VDD.n2937 0.013
R14556 VDD.n263 VDD.n262 0.013
R14557 VDD.n367 VDD.n355 0.013
R14558 VDD.n1974 VDD.n1973 0.013
R14559 VDD.n2009 VDD.n1992 0.013
R14560 VDD.n2517 VDD.n2516 0.013
R14561 VDD.n2527 VDD.n2520 0.013
R14562 VDD.n2566 VDD.n2565 0.013
R14563 VDD.n2563 VDD.n2550 0.013
R14564 VDD.n2550 VDD.n2549 0.013
R14565 VDD.n137 VDD.n136 0.013
R14566 VDD.n5166 VDD.n5165 0.013
R14567 VDD.n5210 VDD.n5209 0.013
R14568 VDD.n5224 VDD.n5212 0.013
R14569 VDD.n5274 VDD.n5273 0.013
R14570 VDD.n5250 VDD.n5249 0.013
R14571 VDD.n2645 VDD.n2633 0.013
R14572 VDD.n2676 VDD.n2675 0.013
R14573 VDD.n2710 VDD.n2709 0.013
R14574 VDD.n2729 VDD.n2728 0.013
R14575 VDD.n2748 VDD.n2747 0.013
R14576 VDD.n5100 VDD.n5087 0.013
R14577 VDD.n97 VDD.n96 0.013
R14578 VDD.n5304 VDD.n5303 0.013
R14579 VDD.n5301 VDD.n5300 0.013
R14580 VDD.n2702 VDD.n2701 0.013
R14581 VDD.n2708 VDD.n2707 0.013
R14582 VDD.n5376 VDD.n5375 0.013
R14583 VDD.n5479 VDD.n5478 0.013
R14584 VDD.n5659 VDD.n5656 0.013
R14585 VDD.n5313 VDD.n5312 0.013
R14586 VDD.n5433 VDD.n5432 0.013
R14587 VDD.n5590 VDD.n5589 0.013
R14588 VDD.n5737 VDD.n5736 0.013
R14589 VDD.n5840 VDD.n5839 0.013
R14590 VDD.n6020 VDD.n6017 0.013
R14591 VDD.n5674 VDD.n5673 0.013
R14592 VDD.n5794 VDD.n5793 0.013
R14593 VDD.n5951 VDD.n5950 0.013
R14594 VDD.n6099 VDD.n6098 0.013
R14595 VDD.n6202 VDD.n6201 0.013
R14596 VDD.n6382 VDD.n6379 0.013
R14597 VDD.n6036 VDD.n6035 0.013
R14598 VDD.n6156 VDD.n6155 0.013
R14599 VDD.n6313 VDD.n6312 0.013
R14600 VDD.n6461 VDD.n6460 0.013
R14601 VDD.n6564 VDD.n6563 0.013
R14602 VDD.n6744 VDD.n6741 0.013
R14603 VDD.n6398 VDD.n6397 0.013
R14604 VDD.n6518 VDD.n6517 0.013
R14605 VDD.n6675 VDD.n6674 0.013
R14606 VDD.n6823 VDD.n6822 0.013
R14607 VDD.n6926 VDD.n6925 0.013
R14608 VDD.n7106 VDD.n7103 0.013
R14609 VDD.n6760 VDD.n6759 0.013
R14610 VDD.n6880 VDD.n6879 0.013
R14611 VDD.n7037 VDD.n7036 0.013
R14612 VDD.n7185 VDD.n7184 0.013
R14613 VDD.n7288 VDD.n7287 0.013
R14614 VDD.n7468 VDD.n7465 0.013
R14615 VDD.n7122 VDD.n7121 0.013
R14616 VDD.n7242 VDD.n7241 0.013
R14617 VDD.n7399 VDD.n7398 0.013
R14618 VDD.n7547 VDD.n7546 0.013
R14619 VDD.n7650 VDD.n7649 0.013
R14620 VDD.n7830 VDD.n7827 0.013
R14621 VDD.n7484 VDD.n7483 0.013
R14622 VDD.n7604 VDD.n7603 0.013
R14623 VDD.n7761 VDD.n7760 0.013
R14624 VDD.n7909 VDD.n7908 0.013
R14625 VDD.n8012 VDD.n8011 0.013
R14626 VDD.n8192 VDD.n8189 0.013
R14627 VDD.n7846 VDD.n7845 0.013
R14628 VDD.n7966 VDD.n7965 0.013
R14629 VDD.n8123 VDD.n8122 0.013
R14630 VDD.n8271 VDD.n8270 0.013
R14631 VDD.n8374 VDD.n8373 0.013
R14632 VDD.n8554 VDD.n8551 0.013
R14633 VDD.n8208 VDD.n8207 0.013
R14634 VDD.n8328 VDD.n8327 0.013
R14635 VDD.n8485 VDD.n8484 0.013
R14636 VDD.n8633 VDD.n8632 0.013
R14637 VDD.n8736 VDD.n8735 0.013
R14638 VDD.n8916 VDD.n8913 0.013
R14639 VDD.n8570 VDD.n8569 0.013
R14640 VDD.n8690 VDD.n8689 0.013
R14641 VDD.n8847 VDD.n8846 0.013
R14642 VDD.n8995 VDD.n8994 0.013
R14643 VDD.n9098 VDD.n9097 0.013
R14644 VDD.n9278 VDD.n9275 0.013
R14645 VDD.n8932 VDD.n8931 0.013
R14646 VDD.n9052 VDD.n9051 0.013
R14647 VDD.n9209 VDD.n9208 0.013
R14648 VDD.n9357 VDD.n9356 0.013
R14649 VDD.n9460 VDD.n9459 0.013
R14650 VDD.n9640 VDD.n9637 0.013
R14651 VDD.n9294 VDD.n9293 0.013
R14652 VDD.n9414 VDD.n9413 0.013
R14653 VDD.n9571 VDD.n9570 0.013
R14654 VDD.n9719 VDD.n9718 0.013
R14655 VDD.n9822 VDD.n9821 0.013
R14656 VDD.n10002 VDD.n9999 0.013
R14657 VDD.n9656 VDD.n9655 0.013
R14658 VDD.n9776 VDD.n9775 0.013
R14659 VDD.n9933 VDD.n9932 0.013
R14660 VDD.n10324 VDD.n10322 0.013
R14661 VDD.n10260 VDD.n10251 0.013
R14662 VDD.n10205 VDD.n10203 0.013
R14663 VDD.n10143 VDD.n10135 0.013
R14664 VDD.n10671 VDD.n10669 0.013
R14665 VDD.n10607 VDD.n10598 0.013
R14666 VDD.n10551 VDD.n10549 0.013
R14667 VDD.n10489 VDD.n10481 0.013
R14668 VDD.n11555 VDD.n11554 0.013
R14669 VDD.n10785 VDD.n10784 0.013
R14670 VDD.n10892 VDD.n10890 0.013
R14671 VDD.n10955 VDD.n10954 0.013
R14672 VDD.n10764 VDD.n10763 0.013
R14673 VDD.n10771 VDD.n10770 0.013
R14674 VDD.n10718 VDD.n10716 0.013
R14675 VDD.n11661 VDD.n11659 0.013
R14676 VDD.n11724 VDD.n11723 0.013
R14677 VDD.n11534 VDD.n11533 0.013
R14678 VDD.n11541 VDD.n11540 0.013
R14679 VDD.n11488 VDD.n11486 0.013
R14680 VDD.n12113 VDD.n12104 0.013
R14681 VDD.n12070 VDD.n12068 0.013
R14682 VDD.n11345 VDD.n11337 0.013
R14683 VDD.n11301 VDD.n11299 0.013
R14684 VDD.n5031 VDD.n5029 0.012
R14685 VDD.n4968 VDD.n4966 0.012
R14686 VDD.n4800 VDD.n4798 0.012
R14687 VDD.n4737 VDD.n4735 0.012
R14688 VDD.n2976 VDD.n2964 0.012
R14689 VDD.n3043 VDD.n3042 0.012
R14690 VDD.n3214 VDD.n3202 0.012
R14691 VDD.n3280 VDD.n3279 0.012
R14692 VDD.n3451 VDD.n3439 0.012
R14693 VDD.n3518 VDD.n3517 0.012
R14694 VDD.n3689 VDD.n3677 0.012
R14695 VDD.n3755 VDD.n3754 0.012
R14696 VDD.n3926 VDD.n3914 0.012
R14697 VDD.n3993 VDD.n3992 0.012
R14698 VDD.n4164 VDD.n4152 0.012
R14699 VDD.n4230 VDD.n4229 0.012
R14700 VDD.n4401 VDD.n4389 0.012
R14701 VDD.n4473 VDD.n4472 0.012
R14702 VDD.n393 VDD.n381 0.012
R14703 VDD.n463 VDD.n462 0.012
R14704 VDD.n627 VDD.n615 0.012
R14705 VDD.n696 VDD.n695 0.012
R14706 VDD.n860 VDD.n848 0.012
R14707 VDD.n930 VDD.n929 0.012
R14708 VDD.n1094 VDD.n1082 0.012
R14709 VDD.n1163 VDD.n1162 0.012
R14710 VDD.n1327 VDD.n1315 0.012
R14711 VDD.n1397 VDD.n1396 0.012
R14712 VDD.n1561 VDD.n1549 0.012
R14713 VDD.n1630 VDD.n1629 0.012
R14714 VDD.n1794 VDD.n1782 0.012
R14715 VDD.n1868 VDD.n1867 0.012
R14716 VDD.n2133 VDD.n2131 0.012
R14717 VDD.n2196 VDD.n2194 0.012
R14718 VDD.n2364 VDD.n2362 0.012
R14719 VDD.n2427 VDD.n2425 0.012
R14720 VDD.n12225 VDD.n12223 0.012
R14721 VDD.n12154 VDD.n12152 0.012
R14722 VDD.n12022 VDD.n12020 0.012
R14723 VDD.n11453 VDD.n11451 0.012
R14724 VDD.n11385 VDD.n11383 0.012
R14725 VDD.n11255 VDD.n11253 0.012
R14726 VDD.n4572 VDD.n4571 0.011
R14727 VDD.n4594 VDD.n4593 0.011
R14728 VDD.n2819 VDD.n2818 0.011
R14729 VDD.n2933 VDD.n2932 0.011
R14730 VDD.n243 VDD.n242 0.011
R14731 VDD.n1966 VDD.n1965 0.011
R14732 VDD.n1988 VDD.n1987 0.011
R14733 VDD.n2503 VDD.n2502 0.011
R14734 VDD.n5153 VDD.n5152 0.011
R14735 VDD.n5185 VDD.n5184 0.011
R14736 VDD.n5186 VDD.n5185 0.011
R14737 VDD.n5289 VDD.n5277 0.011
R14738 VDD.n5251 VDD.n5250 0.011
R14739 VDD.n2647 VDD.n2646 0.011
R14740 VDD.n2741 VDD.n2731 0.011
R14741 VDD.n5107 VDD.n5106 0.011
R14742 VDD.n5101 VDD.n5100 0.011
R14743 VDD.n5366 VDD.n5365 0.011
R14744 VDD.n5342 VDD.n5341 0.011
R14745 VDD.n5610 VDD.n5609 0.011
R14746 VDD.n5644 VDD.n5643 0.011
R14747 VDD.n5727 VDD.n5726 0.011
R14748 VDD.n5703 VDD.n5702 0.011
R14749 VDD.n5971 VDD.n5970 0.011
R14750 VDD.n6005 VDD.n6004 0.011
R14751 VDD.n6089 VDD.n6088 0.011
R14752 VDD.n6065 VDD.n6064 0.011
R14753 VDD.n6333 VDD.n6332 0.011
R14754 VDD.n6367 VDD.n6366 0.011
R14755 VDD.n6451 VDD.n6450 0.011
R14756 VDD.n6427 VDD.n6426 0.011
R14757 VDD.n6695 VDD.n6694 0.011
R14758 VDD.n6729 VDD.n6728 0.011
R14759 VDD.n6813 VDD.n6812 0.011
R14760 VDD.n6789 VDD.n6788 0.011
R14761 VDD.n7057 VDD.n7056 0.011
R14762 VDD.n7091 VDD.n7090 0.011
R14763 VDD.n7175 VDD.n7174 0.011
R14764 VDD.n7151 VDD.n7150 0.011
R14765 VDD.n7419 VDD.n7418 0.011
R14766 VDD.n7453 VDD.n7452 0.011
R14767 VDD.n7537 VDD.n7536 0.011
R14768 VDD.n7513 VDD.n7512 0.011
R14769 VDD.n7781 VDD.n7780 0.011
R14770 VDD.n7815 VDD.n7814 0.011
R14771 VDD.n7899 VDD.n7898 0.011
R14772 VDD.n7875 VDD.n7874 0.011
R14773 VDD.n8143 VDD.n8142 0.011
R14774 VDD.n8177 VDD.n8176 0.011
R14775 VDD.n8261 VDD.n8260 0.011
R14776 VDD.n8237 VDD.n8236 0.011
R14777 VDD.n8505 VDD.n8504 0.011
R14778 VDD.n8539 VDD.n8538 0.011
R14779 VDD.n8623 VDD.n8622 0.011
R14780 VDD.n8599 VDD.n8598 0.011
R14781 VDD.n8867 VDD.n8866 0.011
R14782 VDD.n8901 VDD.n8900 0.011
R14783 VDD.n8985 VDD.n8984 0.011
R14784 VDD.n8961 VDD.n8960 0.011
R14785 VDD.n9229 VDD.n9228 0.011
R14786 VDD.n9263 VDD.n9262 0.011
R14787 VDD.n9347 VDD.n9346 0.011
R14788 VDD.n9323 VDD.n9322 0.011
R14789 VDD.n9591 VDD.n9590 0.011
R14790 VDD.n9625 VDD.n9624 0.011
R14791 VDD.n9709 VDD.n9708 0.011
R14792 VDD.n9685 VDD.n9684 0.011
R14793 VDD.n9953 VDD.n9952 0.011
R14794 VDD.n9987 VDD.n9986 0.011
R14795 VDD.n10896 VDD.n10895 0.011
R14796 VDD.n10909 VDD.n10897 0.011
R14797 VDD.n11013 VDD.n11012 0.011
R14798 VDD.n11103 VDD.n11102 0.011
R14799 VDD.n11665 VDD.n11664 0.011
R14800 VDD.n11677 VDD.n11666 0.011
R14801 VDD.n11781 VDD.n11780 0.011
R14802 VDD.n11877 VDD.n11876 0.011
R14803 VDD.n12125 VDD.n12117 0.011
R14804 VDD.n12057 VDD.n12055 0.011
R14805 VDD.n11357 VDD.n11349 0.011
R14806 VDD.n11289 VDD.n11287 0.011
R14807 VDD.n12142 VDD.n12140 0.01
R14808 VDD.n12034 VDD.n12032 0.01
R14809 VDD.n11373 VDD.n11371 0.01
R14810 VDD.n11267 VDD.n11265 0.01
R14811 VDD.n11462 VDD.n10689 0.01
R14812 VDD.n180 VDD.n179 0.01
R14813 VDD.n1965 VDD.n1964 0.009
R14814 VDD.n4571 VDD.n4570 0.009
R14815 VDD.n2818 VDD.n2817 0.009
R14816 VDD.n242 VDD.n241 0.009
R14817 VDD.n4910 VDD.n4908 0.009
R14818 VDD.n4866 VDD.n4856 0.009
R14819 VDD.n4679 VDD.n4677 0.009
R14820 VDD.n4577 VDD.n4576 0.009
R14821 VDD.n2824 VDD.n2823 0.009
R14822 VDD.n2842 VDD.n2841 0.009
R14823 VDD.n3100 VDD.n3099 0.009
R14824 VDD.n3145 VDD.n3144 0.009
R14825 VDD.n3338 VDD.n3337 0.009
R14826 VDD.n3383 VDD.n3382 0.009
R14827 VDD.n3575 VDD.n3574 0.009
R14828 VDD.n3620 VDD.n3619 0.009
R14829 VDD.n3813 VDD.n3812 0.009
R14830 VDD.n3858 VDD.n3857 0.009
R14831 VDD.n4050 VDD.n4049 0.009
R14832 VDD.n4095 VDD.n4094 0.009
R14833 VDD.n4288 VDD.n4287 0.009
R14834 VDD.n4333 VDD.n4332 0.009
R14835 VDD.n4562 VDD.n4561 0.009
R14836 VDD.n248 VDD.n247 0.009
R14837 VDD.n1971 VDD.n1970 0.009
R14838 VDD.n258 VDD.n257 0.009
R14839 VDD.n520 VDD.n519 0.009
R14840 VDD.n558 VDD.n557 0.009
R14841 VDD.n754 VDD.n753 0.009
R14842 VDD.n792 VDD.n791 0.009
R14843 VDD.n987 VDD.n986 0.009
R14844 VDD.n1025 VDD.n1024 0.009
R14845 VDD.n1221 VDD.n1220 0.009
R14846 VDD.n1259 VDD.n1258 0.009
R14847 VDD.n1454 VDD.n1453 0.009
R14848 VDD.n1492 VDD.n1491 0.009
R14849 VDD.n1688 VDD.n1687 0.009
R14850 VDD.n1726 VDD.n1725 0.009
R14851 VDD.n1947 VDD.n1946 0.009
R14852 VDD.n2075 VDD.n2073 0.009
R14853 VDD.n2262 VDD.n2252 0.009
R14854 VDD.n2306 VDD.n2304 0.009
R14855 VDD.n2497 VDD.n2496 0.009
R14856 VDD.n2502 VDD.n2501 0.009
R14857 VDD.n2574 VDD.n2571 0.009
R14858 VDD.n134 VDD.n133 0.009
R14859 VDD.n155 VDD.n154 0.009
R14860 VDD.n5187 VDD.n5186 0.009
R14861 VDD.n2648 VDD.n2647 0.009
R14862 VDD.n2689 VDD.n2651 0.009
R14863 VDD.n2675 VDD.n2674 0.009
R14864 VDD.n5106 VDD.n5105 0.009
R14865 VDD.n166 VDD.n165 0.009
R14866 VDD.n169 VDD.n168 0.009
R14867 VDD.n2629 VDD.n2628 0.009
R14868 VDD.n5374 VDD.n5372 0.009
R14869 VDD.n5349 VDD.n5348 0.009
R14870 VDD.n5623 VDD.n5622 0.009
R14871 VDD.n5631 VDD.n5630 0.009
R14872 VDD.n5662 VDD.n5661 0.009
R14873 VDD.n5414 VDD.n5413 0.009
R14874 VDD.n5429 VDD.n5428 0.009
R14875 VDD.n5557 VDD.n5555 0.009
R14876 VDD.n5561 VDD.n5560 0.009
R14877 VDD.n5563 VDD.n5562 0.009
R14878 VDD.n5595 VDD.n5594 0.009
R14879 VDD.n5667 VDD.n5598 0.009
R14880 VDD.n5386 VDD.n5385 0.009
R14881 VDD.n5388 VDD.n5387 0.009
R14882 VDD.n5393 VDD.n5392 0.009
R14883 VDD.n5398 VDD.n5394 0.009
R14884 VDD.n5424 VDD.n5423 0.009
R14885 VDD.n5430 VDD.n5425 0.009
R14886 VDD.n5435 VDD.n5434 0.009
R14887 VDD.n5441 VDD.n5436 0.009
R14888 VDD.n5531 VDD.n5530 0.009
R14889 VDD.n5537 VDD.n5532 0.009
R14890 VDD.n5542 VDD.n5541 0.009
R14891 VDD.n5548 VDD.n5543 0.009
R14892 VDD.n5573 VDD.n5572 0.009
R14893 VDD.n5579 VDD.n5574 0.009
R14894 VDD.n5584 VDD.n5583 0.009
R14895 VDD.n5591 VDD.n5585 0.009
R14896 VDD.n5735 VDD.n5733 0.009
R14897 VDD.n5710 VDD.n5709 0.009
R14898 VDD.n5984 VDD.n5983 0.009
R14899 VDD.n5992 VDD.n5991 0.009
R14900 VDD.n6023 VDD.n6022 0.009
R14901 VDD.n5775 VDD.n5774 0.009
R14902 VDD.n5790 VDD.n5789 0.009
R14903 VDD.n5918 VDD.n5916 0.009
R14904 VDD.n5922 VDD.n5921 0.009
R14905 VDD.n5924 VDD.n5923 0.009
R14906 VDD.n5956 VDD.n5955 0.009
R14907 VDD.n6028 VDD.n5959 0.009
R14908 VDD.n5747 VDD.n5746 0.009
R14909 VDD.n5749 VDD.n5748 0.009
R14910 VDD.n5754 VDD.n5753 0.009
R14911 VDD.n5759 VDD.n5755 0.009
R14912 VDD.n5785 VDD.n5784 0.009
R14913 VDD.n5791 VDD.n5786 0.009
R14914 VDD.n5796 VDD.n5795 0.009
R14915 VDD.n5802 VDD.n5797 0.009
R14916 VDD.n5892 VDD.n5891 0.009
R14917 VDD.n5898 VDD.n5893 0.009
R14918 VDD.n5903 VDD.n5902 0.009
R14919 VDD.n5909 VDD.n5904 0.009
R14920 VDD.n5934 VDD.n5933 0.009
R14921 VDD.n5940 VDD.n5935 0.009
R14922 VDD.n5945 VDD.n5944 0.009
R14923 VDD.n5952 VDD.n5946 0.009
R14924 VDD.n6097 VDD.n6095 0.009
R14925 VDD.n6072 VDD.n6071 0.009
R14926 VDD.n6346 VDD.n6345 0.009
R14927 VDD.n6354 VDD.n6353 0.009
R14928 VDD.n6385 VDD.n6384 0.009
R14929 VDD.n6137 VDD.n6136 0.009
R14930 VDD.n6152 VDD.n6151 0.009
R14931 VDD.n6280 VDD.n6278 0.009
R14932 VDD.n6284 VDD.n6283 0.009
R14933 VDD.n6286 VDD.n6285 0.009
R14934 VDD.n6318 VDD.n6317 0.009
R14935 VDD.n6390 VDD.n6321 0.009
R14936 VDD.n6109 VDD.n6108 0.009
R14937 VDD.n6111 VDD.n6110 0.009
R14938 VDD.n6116 VDD.n6115 0.009
R14939 VDD.n6121 VDD.n6117 0.009
R14940 VDD.n6147 VDD.n6146 0.009
R14941 VDD.n6153 VDD.n6148 0.009
R14942 VDD.n6158 VDD.n6157 0.009
R14943 VDD.n6164 VDD.n6159 0.009
R14944 VDD.n6254 VDD.n6253 0.009
R14945 VDD.n6260 VDD.n6255 0.009
R14946 VDD.n6265 VDD.n6264 0.009
R14947 VDD.n6271 VDD.n6266 0.009
R14948 VDD.n6296 VDD.n6295 0.009
R14949 VDD.n6302 VDD.n6297 0.009
R14950 VDD.n6307 VDD.n6306 0.009
R14951 VDD.n6314 VDD.n6308 0.009
R14952 VDD.n6459 VDD.n6457 0.009
R14953 VDD.n6434 VDD.n6433 0.009
R14954 VDD.n6708 VDD.n6707 0.009
R14955 VDD.n6716 VDD.n6715 0.009
R14956 VDD.n6747 VDD.n6746 0.009
R14957 VDD.n6499 VDD.n6498 0.009
R14958 VDD.n6514 VDD.n6513 0.009
R14959 VDD.n6642 VDD.n6640 0.009
R14960 VDD.n6646 VDD.n6645 0.009
R14961 VDD.n6648 VDD.n6647 0.009
R14962 VDD.n6680 VDD.n6679 0.009
R14963 VDD.n6752 VDD.n6683 0.009
R14964 VDD.n6471 VDD.n6470 0.009
R14965 VDD.n6473 VDD.n6472 0.009
R14966 VDD.n6478 VDD.n6477 0.009
R14967 VDD.n6483 VDD.n6479 0.009
R14968 VDD.n6509 VDD.n6508 0.009
R14969 VDD.n6515 VDD.n6510 0.009
R14970 VDD.n6520 VDD.n6519 0.009
R14971 VDD.n6526 VDD.n6521 0.009
R14972 VDD.n6616 VDD.n6615 0.009
R14973 VDD.n6622 VDD.n6617 0.009
R14974 VDD.n6627 VDD.n6626 0.009
R14975 VDD.n6633 VDD.n6628 0.009
R14976 VDD.n6658 VDD.n6657 0.009
R14977 VDD.n6664 VDD.n6659 0.009
R14978 VDD.n6669 VDD.n6668 0.009
R14979 VDD.n6676 VDD.n6670 0.009
R14980 VDD.n6821 VDD.n6819 0.009
R14981 VDD.n6796 VDD.n6795 0.009
R14982 VDD.n7070 VDD.n7069 0.009
R14983 VDD.n7078 VDD.n7077 0.009
R14984 VDD.n7109 VDD.n7108 0.009
R14985 VDD.n6861 VDD.n6860 0.009
R14986 VDD.n6876 VDD.n6875 0.009
R14987 VDD.n7004 VDD.n7002 0.009
R14988 VDD.n7008 VDD.n7007 0.009
R14989 VDD.n7010 VDD.n7009 0.009
R14990 VDD.n7042 VDD.n7041 0.009
R14991 VDD.n7114 VDD.n7045 0.009
R14992 VDD.n6833 VDD.n6832 0.009
R14993 VDD.n6835 VDD.n6834 0.009
R14994 VDD.n6840 VDD.n6839 0.009
R14995 VDD.n6845 VDD.n6841 0.009
R14996 VDD.n6871 VDD.n6870 0.009
R14997 VDD.n6877 VDD.n6872 0.009
R14998 VDD.n6882 VDD.n6881 0.009
R14999 VDD.n6888 VDD.n6883 0.009
R15000 VDD.n6978 VDD.n6977 0.009
R15001 VDD.n6984 VDD.n6979 0.009
R15002 VDD.n6989 VDD.n6988 0.009
R15003 VDD.n6995 VDD.n6990 0.009
R15004 VDD.n7020 VDD.n7019 0.009
R15005 VDD.n7026 VDD.n7021 0.009
R15006 VDD.n7031 VDD.n7030 0.009
R15007 VDD.n7038 VDD.n7032 0.009
R15008 VDD.n7183 VDD.n7181 0.009
R15009 VDD.n7158 VDD.n7157 0.009
R15010 VDD.n7432 VDD.n7431 0.009
R15011 VDD.n7440 VDD.n7439 0.009
R15012 VDD.n7471 VDD.n7470 0.009
R15013 VDD.n7223 VDD.n7222 0.009
R15014 VDD.n7238 VDD.n7237 0.009
R15015 VDD.n7366 VDD.n7364 0.009
R15016 VDD.n7370 VDD.n7369 0.009
R15017 VDD.n7372 VDD.n7371 0.009
R15018 VDD.n7404 VDD.n7403 0.009
R15019 VDD.n7476 VDD.n7407 0.009
R15020 VDD.n7195 VDD.n7194 0.009
R15021 VDD.n7197 VDD.n7196 0.009
R15022 VDD.n7202 VDD.n7201 0.009
R15023 VDD.n7207 VDD.n7203 0.009
R15024 VDD.n7233 VDD.n7232 0.009
R15025 VDD.n7239 VDD.n7234 0.009
R15026 VDD.n7244 VDD.n7243 0.009
R15027 VDD.n7250 VDD.n7245 0.009
R15028 VDD.n7340 VDD.n7339 0.009
R15029 VDD.n7346 VDD.n7341 0.009
R15030 VDD.n7351 VDD.n7350 0.009
R15031 VDD.n7357 VDD.n7352 0.009
R15032 VDD.n7382 VDD.n7381 0.009
R15033 VDD.n7388 VDD.n7383 0.009
R15034 VDD.n7393 VDD.n7392 0.009
R15035 VDD.n7400 VDD.n7394 0.009
R15036 VDD.n7545 VDD.n7543 0.009
R15037 VDD.n7520 VDD.n7519 0.009
R15038 VDD.n7794 VDD.n7793 0.009
R15039 VDD.n7802 VDD.n7801 0.009
R15040 VDD.n7833 VDD.n7832 0.009
R15041 VDD.n7585 VDD.n7584 0.009
R15042 VDD.n7600 VDD.n7599 0.009
R15043 VDD.n7728 VDD.n7726 0.009
R15044 VDD.n7732 VDD.n7731 0.009
R15045 VDD.n7734 VDD.n7733 0.009
R15046 VDD.n7766 VDD.n7765 0.009
R15047 VDD.n7838 VDD.n7769 0.009
R15048 VDD.n7557 VDD.n7556 0.009
R15049 VDD.n7559 VDD.n7558 0.009
R15050 VDD.n7564 VDD.n7563 0.009
R15051 VDD.n7569 VDD.n7565 0.009
R15052 VDD.n7595 VDD.n7594 0.009
R15053 VDD.n7601 VDD.n7596 0.009
R15054 VDD.n7606 VDD.n7605 0.009
R15055 VDD.n7612 VDD.n7607 0.009
R15056 VDD.n7702 VDD.n7701 0.009
R15057 VDD.n7708 VDD.n7703 0.009
R15058 VDD.n7713 VDD.n7712 0.009
R15059 VDD.n7719 VDD.n7714 0.009
R15060 VDD.n7744 VDD.n7743 0.009
R15061 VDD.n7750 VDD.n7745 0.009
R15062 VDD.n7755 VDD.n7754 0.009
R15063 VDD.n7762 VDD.n7756 0.009
R15064 VDD.n7907 VDD.n7905 0.009
R15065 VDD.n7882 VDD.n7881 0.009
R15066 VDD.n8156 VDD.n8155 0.009
R15067 VDD.n8164 VDD.n8163 0.009
R15068 VDD.n8195 VDD.n8194 0.009
R15069 VDD.n7947 VDD.n7946 0.009
R15070 VDD.n7962 VDD.n7961 0.009
R15071 VDD.n8090 VDD.n8088 0.009
R15072 VDD.n8094 VDD.n8093 0.009
R15073 VDD.n8096 VDD.n8095 0.009
R15074 VDD.n8128 VDD.n8127 0.009
R15075 VDD.n8200 VDD.n8131 0.009
R15076 VDD.n7919 VDD.n7918 0.009
R15077 VDD.n7921 VDD.n7920 0.009
R15078 VDD.n7926 VDD.n7925 0.009
R15079 VDD.n7931 VDD.n7927 0.009
R15080 VDD.n7957 VDD.n7956 0.009
R15081 VDD.n7963 VDD.n7958 0.009
R15082 VDD.n7968 VDD.n7967 0.009
R15083 VDD.n7974 VDD.n7969 0.009
R15084 VDD.n8064 VDD.n8063 0.009
R15085 VDD.n8070 VDD.n8065 0.009
R15086 VDD.n8075 VDD.n8074 0.009
R15087 VDD.n8081 VDD.n8076 0.009
R15088 VDD.n8106 VDD.n8105 0.009
R15089 VDD.n8112 VDD.n8107 0.009
R15090 VDD.n8117 VDD.n8116 0.009
R15091 VDD.n8124 VDD.n8118 0.009
R15092 VDD.n8269 VDD.n8267 0.009
R15093 VDD.n8244 VDD.n8243 0.009
R15094 VDD.n8518 VDD.n8517 0.009
R15095 VDD.n8526 VDD.n8525 0.009
R15096 VDD.n8557 VDD.n8556 0.009
R15097 VDD.n8309 VDD.n8308 0.009
R15098 VDD.n8324 VDD.n8323 0.009
R15099 VDD.n8452 VDD.n8450 0.009
R15100 VDD.n8456 VDD.n8455 0.009
R15101 VDD.n8458 VDD.n8457 0.009
R15102 VDD.n8490 VDD.n8489 0.009
R15103 VDD.n8562 VDD.n8493 0.009
R15104 VDD.n8281 VDD.n8280 0.009
R15105 VDD.n8283 VDD.n8282 0.009
R15106 VDD.n8288 VDD.n8287 0.009
R15107 VDD.n8293 VDD.n8289 0.009
R15108 VDD.n8319 VDD.n8318 0.009
R15109 VDD.n8325 VDD.n8320 0.009
R15110 VDD.n8330 VDD.n8329 0.009
R15111 VDD.n8336 VDD.n8331 0.009
R15112 VDD.n8426 VDD.n8425 0.009
R15113 VDD.n8432 VDD.n8427 0.009
R15114 VDD.n8437 VDD.n8436 0.009
R15115 VDD.n8443 VDD.n8438 0.009
R15116 VDD.n8468 VDD.n8467 0.009
R15117 VDD.n8474 VDD.n8469 0.009
R15118 VDD.n8479 VDD.n8478 0.009
R15119 VDD.n8486 VDD.n8480 0.009
R15120 VDD.n8631 VDD.n8629 0.009
R15121 VDD.n8606 VDD.n8605 0.009
R15122 VDD.n8880 VDD.n8879 0.009
R15123 VDD.n8888 VDD.n8887 0.009
R15124 VDD.n8919 VDD.n8918 0.009
R15125 VDD.n8671 VDD.n8670 0.009
R15126 VDD.n8686 VDD.n8685 0.009
R15127 VDD.n8814 VDD.n8812 0.009
R15128 VDD.n8818 VDD.n8817 0.009
R15129 VDD.n8820 VDD.n8819 0.009
R15130 VDD.n8852 VDD.n8851 0.009
R15131 VDD.n8924 VDD.n8855 0.009
R15132 VDD.n8643 VDD.n8642 0.009
R15133 VDD.n8645 VDD.n8644 0.009
R15134 VDD.n8650 VDD.n8649 0.009
R15135 VDD.n8655 VDD.n8651 0.009
R15136 VDD.n8681 VDD.n8680 0.009
R15137 VDD.n8687 VDD.n8682 0.009
R15138 VDD.n8692 VDD.n8691 0.009
R15139 VDD.n8698 VDD.n8693 0.009
R15140 VDD.n8788 VDD.n8787 0.009
R15141 VDD.n8794 VDD.n8789 0.009
R15142 VDD.n8799 VDD.n8798 0.009
R15143 VDD.n8805 VDD.n8800 0.009
R15144 VDD.n8830 VDD.n8829 0.009
R15145 VDD.n8836 VDD.n8831 0.009
R15146 VDD.n8841 VDD.n8840 0.009
R15147 VDD.n8848 VDD.n8842 0.009
R15148 VDD.n8993 VDD.n8991 0.009
R15149 VDD.n8968 VDD.n8967 0.009
R15150 VDD.n9242 VDD.n9241 0.009
R15151 VDD.n9250 VDD.n9249 0.009
R15152 VDD.n9281 VDD.n9280 0.009
R15153 VDD.n9033 VDD.n9032 0.009
R15154 VDD.n9048 VDD.n9047 0.009
R15155 VDD.n9176 VDD.n9174 0.009
R15156 VDD.n9180 VDD.n9179 0.009
R15157 VDD.n9182 VDD.n9181 0.009
R15158 VDD.n9214 VDD.n9213 0.009
R15159 VDD.n9286 VDD.n9217 0.009
R15160 VDD.n9005 VDD.n9004 0.009
R15161 VDD.n9007 VDD.n9006 0.009
R15162 VDD.n9012 VDD.n9011 0.009
R15163 VDD.n9017 VDD.n9013 0.009
R15164 VDD.n9043 VDD.n9042 0.009
R15165 VDD.n9049 VDD.n9044 0.009
R15166 VDD.n9054 VDD.n9053 0.009
R15167 VDD.n9060 VDD.n9055 0.009
R15168 VDD.n9150 VDD.n9149 0.009
R15169 VDD.n9156 VDD.n9151 0.009
R15170 VDD.n9161 VDD.n9160 0.009
R15171 VDD.n9167 VDD.n9162 0.009
R15172 VDD.n9192 VDD.n9191 0.009
R15173 VDD.n9198 VDD.n9193 0.009
R15174 VDD.n9203 VDD.n9202 0.009
R15175 VDD.n9210 VDD.n9204 0.009
R15176 VDD.n9355 VDD.n9353 0.009
R15177 VDD.n9330 VDD.n9329 0.009
R15178 VDD.n9604 VDD.n9603 0.009
R15179 VDD.n9612 VDD.n9611 0.009
R15180 VDD.n9643 VDD.n9642 0.009
R15181 VDD.n9395 VDD.n9394 0.009
R15182 VDD.n9410 VDD.n9409 0.009
R15183 VDD.n9538 VDD.n9536 0.009
R15184 VDD.n9542 VDD.n9541 0.009
R15185 VDD.n9544 VDD.n9543 0.009
R15186 VDD.n9576 VDD.n9575 0.009
R15187 VDD.n9648 VDD.n9579 0.009
R15188 VDD.n9367 VDD.n9366 0.009
R15189 VDD.n9369 VDD.n9368 0.009
R15190 VDD.n9374 VDD.n9373 0.009
R15191 VDD.n9379 VDD.n9375 0.009
R15192 VDD.n9405 VDD.n9404 0.009
R15193 VDD.n9411 VDD.n9406 0.009
R15194 VDD.n9416 VDD.n9415 0.009
R15195 VDD.n9422 VDD.n9417 0.009
R15196 VDD.n9512 VDD.n9511 0.009
R15197 VDD.n9518 VDD.n9513 0.009
R15198 VDD.n9523 VDD.n9522 0.009
R15199 VDD.n9529 VDD.n9524 0.009
R15200 VDD.n9554 VDD.n9553 0.009
R15201 VDD.n9560 VDD.n9555 0.009
R15202 VDD.n9565 VDD.n9564 0.009
R15203 VDD.n9572 VDD.n9566 0.009
R15204 VDD.n9717 VDD.n9715 0.009
R15205 VDD.n9692 VDD.n9691 0.009
R15206 VDD.n9966 VDD.n9965 0.009
R15207 VDD.n9974 VDD.n9973 0.009
R15208 VDD.n10005 VDD.n10004 0.009
R15209 VDD.n9757 VDD.n9756 0.009
R15210 VDD.n9772 VDD.n9771 0.009
R15211 VDD.n9900 VDD.n9898 0.009
R15212 VDD.n9904 VDD.n9903 0.009
R15213 VDD.n9906 VDD.n9905 0.009
R15214 VDD.n9938 VDD.n9937 0.009
R15215 VDD.n10010 VDD.n9941 0.009
R15216 VDD.n9729 VDD.n9728 0.009
R15217 VDD.n9731 VDD.n9730 0.009
R15218 VDD.n9736 VDD.n9735 0.009
R15219 VDD.n9741 VDD.n9737 0.009
R15220 VDD.n9767 VDD.n9766 0.009
R15221 VDD.n9773 VDD.n9768 0.009
R15222 VDD.n9778 VDD.n9777 0.009
R15223 VDD.n9784 VDD.n9779 0.009
R15224 VDD.n9874 VDD.n9873 0.009
R15225 VDD.n9880 VDD.n9875 0.009
R15226 VDD.n9885 VDD.n9884 0.009
R15227 VDD.n9891 VDD.n9886 0.009
R15228 VDD.n9916 VDD.n9915 0.009
R15229 VDD.n9922 VDD.n9917 0.009
R15230 VDD.n9927 VDD.n9926 0.009
R15231 VDD.n9934 VDD.n9928 0.009
R15232 VDD.n10445 VDD.n10438 0.009
R15233 VDD.n10444 VDD.n10443 0.009
R15234 VDD.n10426 VDD.n10425 0.009
R15235 VDD.n10419 VDD.n10402 0.009
R15236 VDD.n10418 VDD.n10417 0.009
R15237 VDD.n10412 VDD.n10408 0.009
R15238 VDD.n10392 VDD.n10375 0.009
R15239 VDD.n10391 VDD.n10390 0.009
R15240 VDD.n10385 VDD.n10381 0.009
R15241 VDD.n10365 VDD.n10358 0.009
R15242 VDD.n10364 VDD.n10363 0.009
R15243 VDD.n10345 VDD.n10344 0.009
R15244 VDD.n10351 VDD.n10350 0.009
R15245 VDD.n10312 VDD.n10310 0.009
R15246 VDD.n10272 VDD.n10264 0.009
R15247 VDD.n10193 VDD.n10191 0.009
R15248 VDD.n10155 VDD.n10147 0.009
R15249 VDD.n10659 VDD.n10657 0.009
R15250 VDD.n10619 VDD.n10611 0.009
R15251 VDD.n10539 VDD.n10537 0.009
R15252 VDD.n10501 VDD.n10493 0.009
R15253 VDD.n11038 VDD.n11037 0.009
R15254 VDD.n11076 VDD.n11075 0.009
R15255 VDD.n11087 VDD.n11076 0.009
R15256 VDD.n10861 VDD.n10860 0.009
R15257 VDD.n10724 VDD.n10723 0.009
R15258 VDD.n10722 VDD.n10721 0.009
R15259 VDD.n11805 VDD.n11804 0.009
R15260 VDD.n11844 VDD.n11843 0.009
R15261 VDD.n11854 VDD.n11844 0.009
R15262 VDD.n11642 VDD.n11641 0.009
R15263 VDD.n11494 VDD.n11493 0.009
R15264 VDD.n11492 VDD.n11491 0.009
R15265 VDD.n12138 VDD.n12129 0.009
R15266 VDD.n12045 VDD.n12043 0.009
R15267 VDD.n11369 VDD.n11361 0.009
R15268 VDD.n11277 VDD.n11275 0.009
R15269 VDD.n2009 VDD.n2008 0.009
R15270 VDD.n367 VDD.n366 0.009
R15271 VDD.n21 VDD.n16 0.008
R15272 VDD.n12129 VDD.n12127 0.008
R15273 VDD.n12047 VDD.n12045 0.008
R15274 VDD.n11361 VDD.n11359 0.008
R15275 VDD.n11279 VDD.n11277 0.008
R15276 VDD.n15 VDD.n14 0.008
R15277 VDD.n12246 VDD.n12245 0.008
R15278 VDD.n2699 VDD.n2698 0.008
R15279 VDD.n2534 VDD.n2533 0.008
R15280 VDD.n180 VDD.n177 0.008
R15281 VDD.n117 VDD.n113 0.008
R15282 VDD.n109 VDD.n106 0.008
R15283 VDD.n2608 VDD.n2605 0.008
R15284 VDD.n2613 VDD.n2612 0.008
R15285 VDD.n2699 VDD.n2696 0.008
R15286 VDD.n2704 VDD.n2703 0.008
R15287 VDD.n5135 VDD.n5134 0.008
R15288 VDD.n4615 VDD.n4614 0.008
R15289 VDD.n2950 VDD.n2949 0.008
R15290 VDD.n184 VDD.n183 0.008
R15291 VDD.n183 VDD.n182 0.007
R15292 VDD.n5017 VDD.n5015 0.007
R15293 VDD.n4982 VDD.n4980 0.007
R15294 VDD.n4786 VDD.n4784 0.007
R15295 VDD.n4751 VDD.n4749 0.007
R15296 VDD.n4583 VDD.n4582 0.007
R15297 VDD.n4588 VDD.n4587 0.007
R15298 VDD.n2879 VDD.n2878 0.007
R15299 VDD.n2990 VDD.n2978 0.007
R15300 VDD.n3029 VDD.n3028 0.007
R15301 VDD.n3228 VDD.n3216 0.007
R15302 VDD.n3266 VDD.n3265 0.007
R15303 VDD.n3465 VDD.n3453 0.007
R15304 VDD.n3504 VDD.n3503 0.007
R15305 VDD.n3703 VDD.n3691 0.007
R15306 VDD.n3741 VDD.n3740 0.007
R15307 VDD.n3940 VDD.n3928 0.007
R15308 VDD.n3979 VDD.n3978 0.007
R15309 VDD.n4178 VDD.n4166 0.007
R15310 VDD.n4216 VDD.n4215 0.007
R15311 VDD.n4415 VDD.n4403 0.007
R15312 VDD.n4454 VDD.n4453 0.007
R15313 VDD.n285 VDD.n284 0.007
R15314 VDD.n294 VDD.n293 0.007
R15315 VDD.n1977 VDD.n1976 0.007
R15316 VDD.n1982 VDD.n1981 0.007
R15317 VDD.n407 VDD.n395 0.007
R15318 VDD.n449 VDD.n448 0.007
R15319 VDD.n641 VDD.n629 0.007
R15320 VDD.n682 VDD.n681 0.007
R15321 VDD.n874 VDD.n862 0.007
R15322 VDD.n916 VDD.n915 0.007
R15323 VDD.n1108 VDD.n1096 0.007
R15324 VDD.n1149 VDD.n1148 0.007
R15325 VDD.n1341 VDD.n1329 0.007
R15326 VDD.n1383 VDD.n1382 0.007
R15327 VDD.n1575 VDD.n1563 0.007
R15328 VDD.n1616 VDD.n1615 0.007
R15329 VDD.n1808 VDD.n1796 0.007
R15330 VDD.n1850 VDD.n1849 0.007
R15331 VDD.n2147 VDD.n2145 0.007
R15332 VDD.n2182 VDD.n2180 0.007
R15333 VDD.n2378 VDD.n2376 0.007
R15334 VDD.n2413 VDD.n2411 0.007
R15335 VDD.n2500 VDD.n2499 0.007
R15336 VDD.n2516 VDD.n2503 0.007
R15337 VDD.n136 VDD.n135 0.007
R15338 VDD.n155 VDD.n149 0.007
R15339 VDD.n5165 VDD.n5153 0.007
R15340 VDD.n5167 VDD.n5166 0.007
R15341 VDD.n5295 VDD.n5294 0.007
R15342 VDD.n5252 VDD.n5251 0.007
R15343 VDD.n2633 VDD.n2632 0.007
R15344 VDD.n2646 VDD.n2645 0.007
R15345 VDD.n2689 VDD.n2688 0.007
R15346 VDD.n2673 VDD.n2672 0.007
R15347 VDD.n2669 VDD.n2656 0.007
R15348 VDD.n187 VDD.n186 0.007
R15349 VDD.n190 VDD.n189 0.007
R15350 VDD.n172 VDD.n171 0.007
R15351 VDD.n161 VDD.n160 0.007
R15352 VDD.n5299 VDD.n5298 0.007
R15353 VDD.n2619 VDD.n2618 0.007
R15354 VDD.n2690 VDD.n2630 0.007
R15355 VDD.n2626 VDD.n2625 0.007
R15356 VDD.n2623 VDD.n2622 0.007
R15357 VDD.n5379 VDD.n5378 0.007
R15358 VDD.n5371 VDD.n5370 0.007
R15359 VDD.n5354 VDD.n5353 0.007
R15360 VDD.n5348 VDD.n5347 0.007
R15361 VDD.n5473 VDD.n5472 0.007
R15362 VDD.n5503 VDD.n5502 0.007
R15363 VDD.n5512 VDD.n5511 0.007
R15364 VDD.n5519 VDD.n5518 0.007
R15365 VDD.n5603 VDD.n5602 0.007
R15366 VDD.n5607 VDD.n5604 0.007
R15367 VDD.n5615 VDD.n5610 0.007
R15368 VDD.n5622 VDD.n5621 0.007
R15369 VDD.n5655 VDD.n5653 0.007
R15370 VDD.n5315 VDD.n5314 0.007
R15371 VDD.n5309 VDD.n5308 0.007
R15372 VDD.n5405 VDD.n5404 0.007
R15373 VDD.n5408 VDD.n5407 0.007
R15374 VDD.n5449 VDD.n5448 0.007
R15375 VDD.n5455 VDD.n5454 0.007
R15376 VDD.n5458 VDD.n5457 0.007
R15377 VDD.n5540 VDD.n5539 0.007
R15378 VDD.n5547 VDD.n5546 0.007
R15379 VDD.n5552 VDD.n5551 0.007
R15380 VDD.n5740 VDD.n5739 0.007
R15381 VDD.n5732 VDD.n5731 0.007
R15382 VDD.n5715 VDD.n5714 0.007
R15383 VDD.n5709 VDD.n5708 0.007
R15384 VDD.n5834 VDD.n5833 0.007
R15385 VDD.n5864 VDD.n5863 0.007
R15386 VDD.n5873 VDD.n5872 0.007
R15387 VDD.n5880 VDD.n5879 0.007
R15388 VDD.n5964 VDD.n5963 0.007
R15389 VDD.n5968 VDD.n5965 0.007
R15390 VDD.n5976 VDD.n5971 0.007
R15391 VDD.n5983 VDD.n5982 0.007
R15392 VDD.n6016 VDD.n6014 0.007
R15393 VDD.n5676 VDD.n5675 0.007
R15394 VDD.n5670 VDD.n5669 0.007
R15395 VDD.n5766 VDD.n5765 0.007
R15396 VDD.n5769 VDD.n5768 0.007
R15397 VDD.n5810 VDD.n5809 0.007
R15398 VDD.n5816 VDD.n5815 0.007
R15399 VDD.n5819 VDD.n5818 0.007
R15400 VDD.n5901 VDD.n5900 0.007
R15401 VDD.n5908 VDD.n5907 0.007
R15402 VDD.n5913 VDD.n5912 0.007
R15403 VDD.n6102 VDD.n6101 0.007
R15404 VDD.n6094 VDD.n6093 0.007
R15405 VDD.n6077 VDD.n6076 0.007
R15406 VDD.n6071 VDD.n6070 0.007
R15407 VDD.n6196 VDD.n6195 0.007
R15408 VDD.n6226 VDD.n6225 0.007
R15409 VDD.n6235 VDD.n6234 0.007
R15410 VDD.n6242 VDD.n6241 0.007
R15411 VDD.n6326 VDD.n6325 0.007
R15412 VDD.n6330 VDD.n6327 0.007
R15413 VDD.n6338 VDD.n6333 0.007
R15414 VDD.n6345 VDD.n6344 0.007
R15415 VDD.n6378 VDD.n6376 0.007
R15416 VDD.n6038 VDD.n6037 0.007
R15417 VDD.n6032 VDD.n6031 0.007
R15418 VDD.n6128 VDD.n6127 0.007
R15419 VDD.n6131 VDD.n6130 0.007
R15420 VDD.n6172 VDD.n6171 0.007
R15421 VDD.n6178 VDD.n6177 0.007
R15422 VDD.n6181 VDD.n6180 0.007
R15423 VDD.n6263 VDD.n6262 0.007
R15424 VDD.n6270 VDD.n6269 0.007
R15425 VDD.n6275 VDD.n6274 0.007
R15426 VDD.n6464 VDD.n6463 0.007
R15427 VDD.n6456 VDD.n6455 0.007
R15428 VDD.n6439 VDD.n6438 0.007
R15429 VDD.n6433 VDD.n6432 0.007
R15430 VDD.n6558 VDD.n6557 0.007
R15431 VDD.n6588 VDD.n6587 0.007
R15432 VDD.n6597 VDD.n6596 0.007
R15433 VDD.n6604 VDD.n6603 0.007
R15434 VDD.n6688 VDD.n6687 0.007
R15435 VDD.n6692 VDD.n6689 0.007
R15436 VDD.n6700 VDD.n6695 0.007
R15437 VDD.n6707 VDD.n6706 0.007
R15438 VDD.n6740 VDD.n6738 0.007
R15439 VDD.n6400 VDD.n6399 0.007
R15440 VDD.n6394 VDD.n6393 0.007
R15441 VDD.n6490 VDD.n6489 0.007
R15442 VDD.n6493 VDD.n6492 0.007
R15443 VDD.n6534 VDD.n6533 0.007
R15444 VDD.n6540 VDD.n6539 0.007
R15445 VDD.n6543 VDD.n6542 0.007
R15446 VDD.n6625 VDD.n6624 0.007
R15447 VDD.n6632 VDD.n6631 0.007
R15448 VDD.n6637 VDD.n6636 0.007
R15449 VDD.n6826 VDD.n6825 0.007
R15450 VDD.n6818 VDD.n6817 0.007
R15451 VDD.n6801 VDD.n6800 0.007
R15452 VDD.n6795 VDD.n6794 0.007
R15453 VDD.n6920 VDD.n6919 0.007
R15454 VDD.n6950 VDD.n6949 0.007
R15455 VDD.n6959 VDD.n6958 0.007
R15456 VDD.n6966 VDD.n6965 0.007
R15457 VDD.n7050 VDD.n7049 0.007
R15458 VDD.n7054 VDD.n7051 0.007
R15459 VDD.n7062 VDD.n7057 0.007
R15460 VDD.n7069 VDD.n7068 0.007
R15461 VDD.n7102 VDD.n7100 0.007
R15462 VDD.n6762 VDD.n6761 0.007
R15463 VDD.n6756 VDD.n6755 0.007
R15464 VDD.n6852 VDD.n6851 0.007
R15465 VDD.n6855 VDD.n6854 0.007
R15466 VDD.n6896 VDD.n6895 0.007
R15467 VDD.n6902 VDD.n6901 0.007
R15468 VDD.n6905 VDD.n6904 0.007
R15469 VDD.n6987 VDD.n6986 0.007
R15470 VDD.n6994 VDD.n6993 0.007
R15471 VDD.n6999 VDD.n6998 0.007
R15472 VDD.n7188 VDD.n7187 0.007
R15473 VDD.n7180 VDD.n7179 0.007
R15474 VDD.n7163 VDD.n7162 0.007
R15475 VDD.n7157 VDD.n7156 0.007
R15476 VDD.n7282 VDD.n7281 0.007
R15477 VDD.n7312 VDD.n7311 0.007
R15478 VDD.n7321 VDD.n7320 0.007
R15479 VDD.n7328 VDD.n7327 0.007
R15480 VDD.n7412 VDD.n7411 0.007
R15481 VDD.n7416 VDD.n7413 0.007
R15482 VDD.n7424 VDD.n7419 0.007
R15483 VDD.n7431 VDD.n7430 0.007
R15484 VDD.n7464 VDD.n7462 0.007
R15485 VDD.n7124 VDD.n7123 0.007
R15486 VDD.n7118 VDD.n7117 0.007
R15487 VDD.n7214 VDD.n7213 0.007
R15488 VDD.n7217 VDD.n7216 0.007
R15489 VDD.n7258 VDD.n7257 0.007
R15490 VDD.n7264 VDD.n7263 0.007
R15491 VDD.n7267 VDD.n7266 0.007
R15492 VDD.n7349 VDD.n7348 0.007
R15493 VDD.n7356 VDD.n7355 0.007
R15494 VDD.n7361 VDD.n7360 0.007
R15495 VDD.n7550 VDD.n7549 0.007
R15496 VDD.n7542 VDD.n7541 0.007
R15497 VDD.n7525 VDD.n7524 0.007
R15498 VDD.n7519 VDD.n7518 0.007
R15499 VDD.n7644 VDD.n7643 0.007
R15500 VDD.n7674 VDD.n7673 0.007
R15501 VDD.n7683 VDD.n7682 0.007
R15502 VDD.n7690 VDD.n7689 0.007
R15503 VDD.n7774 VDD.n7773 0.007
R15504 VDD.n7778 VDD.n7775 0.007
R15505 VDD.n7786 VDD.n7781 0.007
R15506 VDD.n7793 VDD.n7792 0.007
R15507 VDD.n7826 VDD.n7824 0.007
R15508 VDD.n7486 VDD.n7485 0.007
R15509 VDD.n7480 VDD.n7479 0.007
R15510 VDD.n7576 VDD.n7575 0.007
R15511 VDD.n7579 VDD.n7578 0.007
R15512 VDD.n7620 VDD.n7619 0.007
R15513 VDD.n7626 VDD.n7625 0.007
R15514 VDD.n7629 VDD.n7628 0.007
R15515 VDD.n7711 VDD.n7710 0.007
R15516 VDD.n7718 VDD.n7717 0.007
R15517 VDD.n7723 VDD.n7722 0.007
R15518 VDD.n7912 VDD.n7911 0.007
R15519 VDD.n7904 VDD.n7903 0.007
R15520 VDD.n7887 VDD.n7886 0.007
R15521 VDD.n7881 VDD.n7880 0.007
R15522 VDD.n8006 VDD.n8005 0.007
R15523 VDD.n8036 VDD.n8035 0.007
R15524 VDD.n8045 VDD.n8044 0.007
R15525 VDD.n8052 VDD.n8051 0.007
R15526 VDD.n8136 VDD.n8135 0.007
R15527 VDD.n8140 VDD.n8137 0.007
R15528 VDD.n8148 VDD.n8143 0.007
R15529 VDD.n8155 VDD.n8154 0.007
R15530 VDD.n8188 VDD.n8186 0.007
R15531 VDD.n7848 VDD.n7847 0.007
R15532 VDD.n7842 VDD.n7841 0.007
R15533 VDD.n7938 VDD.n7937 0.007
R15534 VDD.n7941 VDD.n7940 0.007
R15535 VDD.n7982 VDD.n7981 0.007
R15536 VDD.n7988 VDD.n7987 0.007
R15537 VDD.n7991 VDD.n7990 0.007
R15538 VDD.n8073 VDD.n8072 0.007
R15539 VDD.n8080 VDD.n8079 0.007
R15540 VDD.n8085 VDD.n8084 0.007
R15541 VDD.n8274 VDD.n8273 0.007
R15542 VDD.n8266 VDD.n8265 0.007
R15543 VDD.n8249 VDD.n8248 0.007
R15544 VDD.n8243 VDD.n8242 0.007
R15545 VDD.n8368 VDD.n8367 0.007
R15546 VDD.n8398 VDD.n8397 0.007
R15547 VDD.n8407 VDD.n8406 0.007
R15548 VDD.n8414 VDD.n8413 0.007
R15549 VDD.n8498 VDD.n8497 0.007
R15550 VDD.n8502 VDD.n8499 0.007
R15551 VDD.n8510 VDD.n8505 0.007
R15552 VDD.n8517 VDD.n8516 0.007
R15553 VDD.n8550 VDD.n8548 0.007
R15554 VDD.n8210 VDD.n8209 0.007
R15555 VDD.n8204 VDD.n8203 0.007
R15556 VDD.n8300 VDD.n8299 0.007
R15557 VDD.n8303 VDD.n8302 0.007
R15558 VDD.n8344 VDD.n8343 0.007
R15559 VDD.n8350 VDD.n8349 0.007
R15560 VDD.n8353 VDD.n8352 0.007
R15561 VDD.n8435 VDD.n8434 0.007
R15562 VDD.n8442 VDD.n8441 0.007
R15563 VDD.n8447 VDD.n8446 0.007
R15564 VDD.n8636 VDD.n8635 0.007
R15565 VDD.n8628 VDD.n8627 0.007
R15566 VDD.n8611 VDD.n8610 0.007
R15567 VDD.n8605 VDD.n8604 0.007
R15568 VDD.n8730 VDD.n8729 0.007
R15569 VDD.n8760 VDD.n8759 0.007
R15570 VDD.n8769 VDD.n8768 0.007
R15571 VDD.n8776 VDD.n8775 0.007
R15572 VDD.n8860 VDD.n8859 0.007
R15573 VDD.n8864 VDD.n8861 0.007
R15574 VDD.n8872 VDD.n8867 0.007
R15575 VDD.n8879 VDD.n8878 0.007
R15576 VDD.n8912 VDD.n8910 0.007
R15577 VDD.n8572 VDD.n8571 0.007
R15578 VDD.n8566 VDD.n8565 0.007
R15579 VDD.n8662 VDD.n8661 0.007
R15580 VDD.n8665 VDD.n8664 0.007
R15581 VDD.n8706 VDD.n8705 0.007
R15582 VDD.n8712 VDD.n8711 0.007
R15583 VDD.n8715 VDD.n8714 0.007
R15584 VDD.n8797 VDD.n8796 0.007
R15585 VDD.n8804 VDD.n8803 0.007
R15586 VDD.n8809 VDD.n8808 0.007
R15587 VDD.n8998 VDD.n8997 0.007
R15588 VDD.n8990 VDD.n8989 0.007
R15589 VDD.n8973 VDD.n8972 0.007
R15590 VDD.n8967 VDD.n8966 0.007
R15591 VDD.n9092 VDD.n9091 0.007
R15592 VDD.n9122 VDD.n9121 0.007
R15593 VDD.n9131 VDD.n9130 0.007
R15594 VDD.n9138 VDD.n9137 0.007
R15595 VDD.n9222 VDD.n9221 0.007
R15596 VDD.n9226 VDD.n9223 0.007
R15597 VDD.n9234 VDD.n9229 0.007
R15598 VDD.n9241 VDD.n9240 0.007
R15599 VDD.n9274 VDD.n9272 0.007
R15600 VDD.n8934 VDD.n8933 0.007
R15601 VDD.n8928 VDD.n8927 0.007
R15602 VDD.n9024 VDD.n9023 0.007
R15603 VDD.n9027 VDD.n9026 0.007
R15604 VDD.n9068 VDD.n9067 0.007
R15605 VDD.n9074 VDD.n9073 0.007
R15606 VDD.n9077 VDD.n9076 0.007
R15607 VDD.n9159 VDD.n9158 0.007
R15608 VDD.n9166 VDD.n9165 0.007
R15609 VDD.n9171 VDD.n9170 0.007
R15610 VDD.n9360 VDD.n9359 0.007
R15611 VDD.n9352 VDD.n9351 0.007
R15612 VDD.n9335 VDD.n9334 0.007
R15613 VDD.n9329 VDD.n9328 0.007
R15614 VDD.n9454 VDD.n9453 0.007
R15615 VDD.n9484 VDD.n9483 0.007
R15616 VDD.n9493 VDD.n9492 0.007
R15617 VDD.n9500 VDD.n9499 0.007
R15618 VDD.n9584 VDD.n9583 0.007
R15619 VDD.n9588 VDD.n9585 0.007
R15620 VDD.n9596 VDD.n9591 0.007
R15621 VDD.n9603 VDD.n9602 0.007
R15622 VDD.n9636 VDD.n9634 0.007
R15623 VDD.n9296 VDD.n9295 0.007
R15624 VDD.n9290 VDD.n9289 0.007
R15625 VDD.n9386 VDD.n9385 0.007
R15626 VDD.n9389 VDD.n9388 0.007
R15627 VDD.n9430 VDD.n9429 0.007
R15628 VDD.n9436 VDD.n9435 0.007
R15629 VDD.n9439 VDD.n9438 0.007
R15630 VDD.n9521 VDD.n9520 0.007
R15631 VDD.n9528 VDD.n9527 0.007
R15632 VDD.n9533 VDD.n9532 0.007
R15633 VDD.n9722 VDD.n9721 0.007
R15634 VDD.n9714 VDD.n9713 0.007
R15635 VDD.n9697 VDD.n9696 0.007
R15636 VDD.n9691 VDD.n9690 0.007
R15637 VDD.n9816 VDD.n9815 0.007
R15638 VDD.n9846 VDD.n9845 0.007
R15639 VDD.n9855 VDD.n9854 0.007
R15640 VDD.n9862 VDD.n9861 0.007
R15641 VDD.n9946 VDD.n9945 0.007
R15642 VDD.n9950 VDD.n9947 0.007
R15643 VDD.n9958 VDD.n9953 0.007
R15644 VDD.n9965 VDD.n9964 0.007
R15645 VDD.n9998 VDD.n9996 0.007
R15646 VDD.n9658 VDD.n9657 0.007
R15647 VDD.n9652 VDD.n9651 0.007
R15648 VDD.n9748 VDD.n9747 0.007
R15649 VDD.n9751 VDD.n9750 0.007
R15650 VDD.n9792 VDD.n9791 0.007
R15651 VDD.n9798 VDD.n9797 0.007
R15652 VDD.n9801 VDD.n9800 0.007
R15653 VDD.n9883 VDD.n9882 0.007
R15654 VDD.n9890 VDD.n9889 0.007
R15655 VDD.n9895 VDD.n9894 0.007
R15656 VDD.n10433 VDD.n10422 0.007
R15657 VDD.n11568 VDD.n11567 0.007
R15658 VDD.n11564 VDD.n11563 0.007
R15659 VDD.n11738 VDD.n11737 0.007
R15660 VDD.n11742 VDD.n11741 0.007
R15661 VDD.n10798 VDD.n10797 0.007
R15662 VDD.n10794 VDD.n10793 0.007
R15663 VDD.n10969 VDD.n10968 0.007
R15664 VDD.n10973 VDD.n10972 0.007
R15665 VDD.n10953 VDD.n10952 0.007
R15666 VDD.n11022 VDD.n11021 0.007
R15667 VDD.n11102 VDD.n11101 0.007
R15668 VDD.n10872 VDD.n10861 0.007
R15669 VDD.n10826 VDD.n10825 0.007
R15670 VDD.n10729 VDD.n10725 0.007
R15671 VDD.n11722 VDD.n11721 0.007
R15672 VDD.n11789 VDD.n11788 0.007
R15673 VDD.n11876 VDD.n11875 0.007
R15674 VDD.n11643 VDD.n11642 0.007
R15675 VDD.n11606 VDD.n11605 0.007
R15676 VDD.n11500 VDD.n11495 0.007
R15677 VDD.n12150 VDD.n12142 0.007
R15678 VDD.n12032 VDD.n12030 0.007
R15679 VDD.n11381 VDD.n11373 0.007
R15680 VDD.n11265 VDD.n11263 0.007
R15681 VDD.n92 VDD.n91 0.007
R15682 VDD.n12250 VDD.n12249 0.007
R15683 VDD.n12117 VDD.n12115 0.006
R15684 VDD.n12059 VDD.n12057 0.006
R15685 VDD.n11349 VDD.n11347 0.006
R15686 VDD.n11291 VDD.n11289 0.006
R15687 VDD.n5136 VDD.n5135 0.006
R15688 VDD.n94 VDD.n93 0.006
R15689 VDD.n10367 VDD.n10366 0.005
R15690 VDD.n10394 VDD.n10393 0.005
R15691 VDD.n10421 VDD.n10420 0.005
R15692 VDD.n10447 VDD.n10446 0.005
R15693 VDD.n7 VDD.n5 0.005
R15694 VDD.n2483 VDD.n2482 0.005
R15695 VDD.n2570 VDD.n2569 0.005
R15696 VDD.n2549 VDD.n2548 0.005
R15697 VDD.n2545 VDD.n2544 0.005
R15698 VDD.n5171 VDD.n5170 0.005
R15699 VDD.n5191 VDD.n5190 0.005
R15700 VDD.n5192 VDD.n5191 0.005
R15701 VDD.n5226 VDD.n5225 0.005
R15702 VDD.n5233 VDD.n5232 0.005
R15703 VDD.n5291 VDD.n5290 0.005
R15704 VDD.n5257 VDD.n5256 0.005
R15705 VDD.n5256 VDD.n5255 0.005
R15706 VDD.n5236 VDD.n5235 0.005
R15707 VDD.n2656 VDD.n2655 0.005
R15708 VDD.n2730 VDD.n2729 0.005
R15709 VDD.n5120 VDD.n5107 0.005
R15710 VDD.n5104 VDD.n5103 0.005
R15711 VDD.n5087 VDD.n5086 0.005
R15712 VDD.n182 VDD.n181 0.005
R15713 VDD.n2533 VDD.n2532 0.005
R15714 VDD.n177 VDD.n176 0.005
R15715 VDD.n113 VDD.n112 0.005
R15716 VDD.n106 VDD.n105 0.005
R15717 VDD.n101 VDD.n100 0.005
R15718 VDD.n2605 VDD.n2604 0.005
R15719 VDD.n2612 VDD.n2611 0.005
R15720 VDD.n2696 VDD.n2695 0.005
R15721 VDD.n2703 VDD.n2702 0.005
R15722 VDD.n5142 VDD.n5141 0.005
R15723 VDD.n5139 VDD.n5138 0.005
R15724 VDD.n5134 VDD.n5133 0.005
R15725 VDD.n5368 VDD.n5367 0.005
R15726 VDD.n5365 VDD.n5363 0.005
R15727 VDD.n5351 VDD.n5350 0.005
R15728 VDD.n5345 VDD.n5344 0.005
R15729 VDD.n5343 VDD.n5342 0.005
R15730 VDD.n5340 VDD.n5339 0.005
R15731 VDD.n5339 VDD.n5336 0.005
R15732 VDD.n5466 VDD.n5465 0.005
R15733 VDD.n5495 VDD.n5492 0.005
R15734 VDD.n5501 VDD.n5500 0.005
R15735 VDD.n5617 VDD.n5616 0.005
R15736 VDD.n5625 VDD.n5624 0.005
R15737 VDD.n5652 VDD.n5651 0.005
R15738 VDD.n5414 VDD.n5411 0.005
R15739 VDD.n5420 VDD.n5419 0.005
R15740 VDD.n5422 VDD.n5421 0.005
R15741 VDD.n5453 VDD.n5452 0.005
R15742 VDD.n5557 VDD.n5556 0.005
R15743 VDD.n5582 VDD.n5581 0.005
R15744 VDD.n5387 VDD.n5386 0.005
R15745 VDD.n5394 VDD.n5393 0.005
R15746 VDD.n5425 VDD.n5424 0.005
R15747 VDD.n5436 VDD.n5435 0.005
R15748 VDD.n5532 VDD.n5531 0.005
R15749 VDD.n5543 VDD.n5542 0.005
R15750 VDD.n5574 VDD.n5573 0.005
R15751 VDD.n5585 VDD.n5584 0.005
R15752 VDD.n5729 VDD.n5728 0.005
R15753 VDD.n5726 VDD.n5724 0.005
R15754 VDD.n5712 VDD.n5711 0.005
R15755 VDD.n5706 VDD.n5705 0.005
R15756 VDD.n5704 VDD.n5703 0.005
R15757 VDD.n5701 VDD.n5700 0.005
R15758 VDD.n5700 VDD.n5697 0.005
R15759 VDD.n5827 VDD.n5826 0.005
R15760 VDD.n5856 VDD.n5853 0.005
R15761 VDD.n5862 VDD.n5861 0.005
R15762 VDD.n5978 VDD.n5977 0.005
R15763 VDD.n5986 VDD.n5985 0.005
R15764 VDD.n6013 VDD.n6012 0.005
R15765 VDD.n5775 VDD.n5772 0.005
R15766 VDD.n5781 VDD.n5780 0.005
R15767 VDD.n5783 VDD.n5782 0.005
R15768 VDD.n5814 VDD.n5813 0.005
R15769 VDD.n5918 VDD.n5917 0.005
R15770 VDD.n5943 VDD.n5942 0.005
R15771 VDD.n5748 VDD.n5747 0.005
R15772 VDD.n5755 VDD.n5754 0.005
R15773 VDD.n5786 VDD.n5785 0.005
R15774 VDD.n5797 VDD.n5796 0.005
R15775 VDD.n5893 VDD.n5892 0.005
R15776 VDD.n5904 VDD.n5903 0.005
R15777 VDD.n5935 VDD.n5934 0.005
R15778 VDD.n5946 VDD.n5945 0.005
R15779 VDD.n6091 VDD.n6090 0.005
R15780 VDD.n6088 VDD.n6086 0.005
R15781 VDD.n6074 VDD.n6073 0.005
R15782 VDD.n6068 VDD.n6067 0.005
R15783 VDD.n6066 VDD.n6065 0.005
R15784 VDD.n6063 VDD.n6062 0.005
R15785 VDD.n6062 VDD.n6059 0.005
R15786 VDD.n6189 VDD.n6188 0.005
R15787 VDD.n6218 VDD.n6215 0.005
R15788 VDD.n6224 VDD.n6223 0.005
R15789 VDD.n6340 VDD.n6339 0.005
R15790 VDD.n6348 VDD.n6347 0.005
R15791 VDD.n6375 VDD.n6374 0.005
R15792 VDD.n6137 VDD.n6134 0.005
R15793 VDD.n6143 VDD.n6142 0.005
R15794 VDD.n6145 VDD.n6144 0.005
R15795 VDD.n6176 VDD.n6175 0.005
R15796 VDD.n6280 VDD.n6279 0.005
R15797 VDD.n6305 VDD.n6304 0.005
R15798 VDD.n6110 VDD.n6109 0.005
R15799 VDD.n6117 VDD.n6116 0.005
R15800 VDD.n6148 VDD.n6147 0.005
R15801 VDD.n6159 VDD.n6158 0.005
R15802 VDD.n6255 VDD.n6254 0.005
R15803 VDD.n6266 VDD.n6265 0.005
R15804 VDD.n6297 VDD.n6296 0.005
R15805 VDD.n6308 VDD.n6307 0.005
R15806 VDD.n6453 VDD.n6452 0.005
R15807 VDD.n6450 VDD.n6448 0.005
R15808 VDD.n6436 VDD.n6435 0.005
R15809 VDD.n6430 VDD.n6429 0.005
R15810 VDD.n6428 VDD.n6427 0.005
R15811 VDD.n6425 VDD.n6424 0.005
R15812 VDD.n6424 VDD.n6421 0.005
R15813 VDD.n6551 VDD.n6550 0.005
R15814 VDD.n6580 VDD.n6577 0.005
R15815 VDD.n6586 VDD.n6585 0.005
R15816 VDD.n6702 VDD.n6701 0.005
R15817 VDD.n6710 VDD.n6709 0.005
R15818 VDD.n6737 VDD.n6736 0.005
R15819 VDD.n6499 VDD.n6496 0.005
R15820 VDD.n6505 VDD.n6504 0.005
R15821 VDD.n6507 VDD.n6506 0.005
R15822 VDD.n6538 VDD.n6537 0.005
R15823 VDD.n6642 VDD.n6641 0.005
R15824 VDD.n6667 VDD.n6666 0.005
R15825 VDD.n6472 VDD.n6471 0.005
R15826 VDD.n6479 VDD.n6478 0.005
R15827 VDD.n6510 VDD.n6509 0.005
R15828 VDD.n6521 VDD.n6520 0.005
R15829 VDD.n6617 VDD.n6616 0.005
R15830 VDD.n6628 VDD.n6627 0.005
R15831 VDD.n6659 VDD.n6658 0.005
R15832 VDD.n6670 VDD.n6669 0.005
R15833 VDD.n6815 VDD.n6814 0.005
R15834 VDD.n6812 VDD.n6810 0.005
R15835 VDD.n6798 VDD.n6797 0.005
R15836 VDD.n6792 VDD.n6791 0.005
R15837 VDD.n6790 VDD.n6789 0.005
R15838 VDD.n6787 VDD.n6786 0.005
R15839 VDD.n6786 VDD.n6783 0.005
R15840 VDD.n6913 VDD.n6912 0.005
R15841 VDD.n6942 VDD.n6939 0.005
R15842 VDD.n6948 VDD.n6947 0.005
R15843 VDD.n7064 VDD.n7063 0.005
R15844 VDD.n7072 VDD.n7071 0.005
R15845 VDD.n7099 VDD.n7098 0.005
R15846 VDD.n6861 VDD.n6858 0.005
R15847 VDD.n6867 VDD.n6866 0.005
R15848 VDD.n6869 VDD.n6868 0.005
R15849 VDD.n6900 VDD.n6899 0.005
R15850 VDD.n7004 VDD.n7003 0.005
R15851 VDD.n7029 VDD.n7028 0.005
R15852 VDD.n6834 VDD.n6833 0.005
R15853 VDD.n6841 VDD.n6840 0.005
R15854 VDD.n6872 VDD.n6871 0.005
R15855 VDD.n6883 VDD.n6882 0.005
R15856 VDD.n6979 VDD.n6978 0.005
R15857 VDD.n6990 VDD.n6989 0.005
R15858 VDD.n7021 VDD.n7020 0.005
R15859 VDD.n7032 VDD.n7031 0.005
R15860 VDD.n7177 VDD.n7176 0.005
R15861 VDD.n7174 VDD.n7172 0.005
R15862 VDD.n7160 VDD.n7159 0.005
R15863 VDD.n7154 VDD.n7153 0.005
R15864 VDD.n7152 VDD.n7151 0.005
R15865 VDD.n7149 VDD.n7148 0.005
R15866 VDD.n7148 VDD.n7145 0.005
R15867 VDD.n7275 VDD.n7274 0.005
R15868 VDD.n7304 VDD.n7301 0.005
R15869 VDD.n7310 VDD.n7309 0.005
R15870 VDD.n7426 VDD.n7425 0.005
R15871 VDD.n7434 VDD.n7433 0.005
R15872 VDD.n7461 VDD.n7460 0.005
R15873 VDD.n7223 VDD.n7220 0.005
R15874 VDD.n7229 VDD.n7228 0.005
R15875 VDD.n7231 VDD.n7230 0.005
R15876 VDD.n7262 VDD.n7261 0.005
R15877 VDD.n7366 VDD.n7365 0.005
R15878 VDD.n7391 VDD.n7390 0.005
R15879 VDD.n7196 VDD.n7195 0.005
R15880 VDD.n7203 VDD.n7202 0.005
R15881 VDD.n7234 VDD.n7233 0.005
R15882 VDD.n7245 VDD.n7244 0.005
R15883 VDD.n7341 VDD.n7340 0.005
R15884 VDD.n7352 VDD.n7351 0.005
R15885 VDD.n7383 VDD.n7382 0.005
R15886 VDD.n7394 VDD.n7393 0.005
R15887 VDD.n7539 VDD.n7538 0.005
R15888 VDD.n7536 VDD.n7534 0.005
R15889 VDD.n7522 VDD.n7521 0.005
R15890 VDD.n7516 VDD.n7515 0.005
R15891 VDD.n7514 VDD.n7513 0.005
R15892 VDD.n7511 VDD.n7510 0.005
R15893 VDD.n7510 VDD.n7507 0.005
R15894 VDD.n7637 VDD.n7636 0.005
R15895 VDD.n7666 VDD.n7663 0.005
R15896 VDD.n7672 VDD.n7671 0.005
R15897 VDD.n7788 VDD.n7787 0.005
R15898 VDD.n7796 VDD.n7795 0.005
R15899 VDD.n7823 VDD.n7822 0.005
R15900 VDD.n7585 VDD.n7582 0.005
R15901 VDD.n7591 VDD.n7590 0.005
R15902 VDD.n7593 VDD.n7592 0.005
R15903 VDD.n7624 VDD.n7623 0.005
R15904 VDD.n7728 VDD.n7727 0.005
R15905 VDD.n7753 VDD.n7752 0.005
R15906 VDD.n7558 VDD.n7557 0.005
R15907 VDD.n7565 VDD.n7564 0.005
R15908 VDD.n7596 VDD.n7595 0.005
R15909 VDD.n7607 VDD.n7606 0.005
R15910 VDD.n7703 VDD.n7702 0.005
R15911 VDD.n7714 VDD.n7713 0.005
R15912 VDD.n7745 VDD.n7744 0.005
R15913 VDD.n7756 VDD.n7755 0.005
R15914 VDD.n7901 VDD.n7900 0.005
R15915 VDD.n7898 VDD.n7896 0.005
R15916 VDD.n7884 VDD.n7883 0.005
R15917 VDD.n7878 VDD.n7877 0.005
R15918 VDD.n7876 VDD.n7875 0.005
R15919 VDD.n7873 VDD.n7872 0.005
R15920 VDD.n7872 VDD.n7869 0.005
R15921 VDD.n7999 VDD.n7998 0.005
R15922 VDD.n8028 VDD.n8025 0.005
R15923 VDD.n8034 VDD.n8033 0.005
R15924 VDD.n8150 VDD.n8149 0.005
R15925 VDD.n8158 VDD.n8157 0.005
R15926 VDD.n8185 VDD.n8184 0.005
R15927 VDD.n7947 VDD.n7944 0.005
R15928 VDD.n7953 VDD.n7952 0.005
R15929 VDD.n7955 VDD.n7954 0.005
R15930 VDD.n7986 VDD.n7985 0.005
R15931 VDD.n8090 VDD.n8089 0.005
R15932 VDD.n8115 VDD.n8114 0.005
R15933 VDD.n7920 VDD.n7919 0.005
R15934 VDD.n7927 VDD.n7926 0.005
R15935 VDD.n7958 VDD.n7957 0.005
R15936 VDD.n7969 VDD.n7968 0.005
R15937 VDD.n8065 VDD.n8064 0.005
R15938 VDD.n8076 VDD.n8075 0.005
R15939 VDD.n8107 VDD.n8106 0.005
R15940 VDD.n8118 VDD.n8117 0.005
R15941 VDD.n8263 VDD.n8262 0.005
R15942 VDD.n8260 VDD.n8258 0.005
R15943 VDD.n8246 VDD.n8245 0.005
R15944 VDD.n8240 VDD.n8239 0.005
R15945 VDD.n8238 VDD.n8237 0.005
R15946 VDD.n8235 VDD.n8234 0.005
R15947 VDD.n8234 VDD.n8231 0.005
R15948 VDD.n8361 VDD.n8360 0.005
R15949 VDD.n8390 VDD.n8387 0.005
R15950 VDD.n8396 VDD.n8395 0.005
R15951 VDD.n8512 VDD.n8511 0.005
R15952 VDD.n8520 VDD.n8519 0.005
R15953 VDD.n8547 VDD.n8546 0.005
R15954 VDD.n8309 VDD.n8306 0.005
R15955 VDD.n8315 VDD.n8314 0.005
R15956 VDD.n8317 VDD.n8316 0.005
R15957 VDD.n8348 VDD.n8347 0.005
R15958 VDD.n8452 VDD.n8451 0.005
R15959 VDD.n8477 VDD.n8476 0.005
R15960 VDD.n8282 VDD.n8281 0.005
R15961 VDD.n8289 VDD.n8288 0.005
R15962 VDD.n8320 VDD.n8319 0.005
R15963 VDD.n8331 VDD.n8330 0.005
R15964 VDD.n8427 VDD.n8426 0.005
R15965 VDD.n8438 VDD.n8437 0.005
R15966 VDD.n8469 VDD.n8468 0.005
R15967 VDD.n8480 VDD.n8479 0.005
R15968 VDD.n8625 VDD.n8624 0.005
R15969 VDD.n8622 VDD.n8620 0.005
R15970 VDD.n8608 VDD.n8607 0.005
R15971 VDD.n8602 VDD.n8601 0.005
R15972 VDD.n8600 VDD.n8599 0.005
R15973 VDD.n8597 VDD.n8596 0.005
R15974 VDD.n8596 VDD.n8593 0.005
R15975 VDD.n8723 VDD.n8722 0.005
R15976 VDD.n8752 VDD.n8749 0.005
R15977 VDD.n8758 VDD.n8757 0.005
R15978 VDD.n8874 VDD.n8873 0.005
R15979 VDD.n8882 VDD.n8881 0.005
R15980 VDD.n8909 VDD.n8908 0.005
R15981 VDD.n8671 VDD.n8668 0.005
R15982 VDD.n8677 VDD.n8676 0.005
R15983 VDD.n8679 VDD.n8678 0.005
R15984 VDD.n8710 VDD.n8709 0.005
R15985 VDD.n8814 VDD.n8813 0.005
R15986 VDD.n8839 VDD.n8838 0.005
R15987 VDD.n8644 VDD.n8643 0.005
R15988 VDD.n8651 VDD.n8650 0.005
R15989 VDD.n8682 VDD.n8681 0.005
R15990 VDD.n8693 VDD.n8692 0.005
R15991 VDD.n8789 VDD.n8788 0.005
R15992 VDD.n8800 VDD.n8799 0.005
R15993 VDD.n8831 VDD.n8830 0.005
R15994 VDD.n8842 VDD.n8841 0.005
R15995 VDD.n8987 VDD.n8986 0.005
R15996 VDD.n8984 VDD.n8982 0.005
R15997 VDD.n8970 VDD.n8969 0.005
R15998 VDD.n8964 VDD.n8963 0.005
R15999 VDD.n8962 VDD.n8961 0.005
R16000 VDD.n8959 VDD.n8958 0.005
R16001 VDD.n8958 VDD.n8955 0.005
R16002 VDD.n9085 VDD.n9084 0.005
R16003 VDD.n9114 VDD.n9111 0.005
R16004 VDD.n9120 VDD.n9119 0.005
R16005 VDD.n9236 VDD.n9235 0.005
R16006 VDD.n9244 VDD.n9243 0.005
R16007 VDD.n9271 VDD.n9270 0.005
R16008 VDD.n9033 VDD.n9030 0.005
R16009 VDD.n9039 VDD.n9038 0.005
R16010 VDD.n9041 VDD.n9040 0.005
R16011 VDD.n9072 VDD.n9071 0.005
R16012 VDD.n9176 VDD.n9175 0.005
R16013 VDD.n9201 VDD.n9200 0.005
R16014 VDD.n9006 VDD.n9005 0.005
R16015 VDD.n9013 VDD.n9012 0.005
R16016 VDD.n9044 VDD.n9043 0.005
R16017 VDD.n9055 VDD.n9054 0.005
R16018 VDD.n9151 VDD.n9150 0.005
R16019 VDD.n9162 VDD.n9161 0.005
R16020 VDD.n9193 VDD.n9192 0.005
R16021 VDD.n9204 VDD.n9203 0.005
R16022 VDD.n9349 VDD.n9348 0.005
R16023 VDD.n9346 VDD.n9344 0.005
R16024 VDD.n9332 VDD.n9331 0.005
R16025 VDD.n9326 VDD.n9325 0.005
R16026 VDD.n9324 VDD.n9323 0.005
R16027 VDD.n9321 VDD.n9320 0.005
R16028 VDD.n9320 VDD.n9317 0.005
R16029 VDD.n9447 VDD.n9446 0.005
R16030 VDD.n9476 VDD.n9473 0.005
R16031 VDD.n9482 VDD.n9481 0.005
R16032 VDD.n9598 VDD.n9597 0.005
R16033 VDD.n9606 VDD.n9605 0.005
R16034 VDD.n9633 VDD.n9632 0.005
R16035 VDD.n9395 VDD.n9392 0.005
R16036 VDD.n9401 VDD.n9400 0.005
R16037 VDD.n9403 VDD.n9402 0.005
R16038 VDD.n9434 VDD.n9433 0.005
R16039 VDD.n9538 VDD.n9537 0.005
R16040 VDD.n9563 VDD.n9562 0.005
R16041 VDD.n9368 VDD.n9367 0.005
R16042 VDD.n9375 VDD.n9374 0.005
R16043 VDD.n9406 VDD.n9405 0.005
R16044 VDD.n9417 VDD.n9416 0.005
R16045 VDD.n9513 VDD.n9512 0.005
R16046 VDD.n9524 VDD.n9523 0.005
R16047 VDD.n9555 VDD.n9554 0.005
R16048 VDD.n9566 VDD.n9565 0.005
R16049 VDD.n9711 VDD.n9710 0.005
R16050 VDD.n9708 VDD.n9706 0.005
R16051 VDD.n9694 VDD.n9693 0.005
R16052 VDD.n9688 VDD.n9687 0.005
R16053 VDD.n9686 VDD.n9685 0.005
R16054 VDD.n9683 VDD.n9682 0.005
R16055 VDD.n9682 VDD.n9679 0.005
R16056 VDD.n9809 VDD.n9808 0.005
R16057 VDD.n9838 VDD.n9835 0.005
R16058 VDD.n9844 VDD.n9843 0.005
R16059 VDD.n9960 VDD.n9959 0.005
R16060 VDD.n9968 VDD.n9967 0.005
R16061 VDD.n9995 VDD.n9994 0.005
R16062 VDD.n9757 VDD.n9754 0.005
R16063 VDD.n9763 VDD.n9762 0.005
R16064 VDD.n9765 VDD.n9764 0.005
R16065 VDD.n9796 VDD.n9795 0.005
R16066 VDD.n9900 VDD.n9899 0.005
R16067 VDD.n9925 VDD.n9924 0.005
R16068 VDD.n9730 VDD.n9729 0.005
R16069 VDD.n9737 VDD.n9736 0.005
R16070 VDD.n9768 VDD.n9767 0.005
R16071 VDD.n9779 VDD.n9778 0.005
R16072 VDD.n9875 VDD.n9874 0.005
R16073 VDD.n9886 VDD.n9885 0.005
R16074 VDD.n9917 VDD.n9916 0.005
R16075 VDD.n9928 VDD.n9927 0.005
R16076 VDD.n10445 VDD.n10444 0.005
R16077 VDD.n10427 VDD.n10426 0.005
R16078 VDD.n10419 VDD.n10418 0.005
R16079 VDD.n10408 VDD.n10407 0.005
R16080 VDD.n10392 VDD.n10391 0.005
R16081 VDD.n10381 VDD.n10380 0.005
R16082 VDD.n10365 VDD.n10364 0.005
R16083 VDD.n10351 VDD.n10345 0.005
R16084 VDD.n11053 VDD.n11041 0.005
R16085 VDD.n11055 VDD.n11054 0.005
R16086 VDD.n11014 VDD.n11013 0.005
R16087 VDD.n11011 VDD.n11010 0.005
R16088 VDD.n10769 VDD.n10768 0.005
R16089 VDD.n10781 VDD.n10771 0.005
R16090 VDD.n11819 VDD.n11808 0.005
R16091 VDD.n11821 VDD.n11820 0.005
R16092 VDD.n11782 VDD.n11781 0.005
R16093 VDD.n11779 VDD.n11778 0.005
R16094 VDD.n11539 VDD.n11538 0.005
R16095 VDD.n11551 VDD.n11541 0.005
R16096 VDD.n12223 VDD.n12221 0.005
R16097 VDD.n12163 VDD.n12154 0.005
R16098 VDD.n12020 VDD.n12018 0.005
R16099 VDD.n11451 VDD.n11449 0.005
R16100 VDD.n11393 VDD.n11385 0.005
R16101 VDD.n11253 VDD.n11251 0.005
R16102 VDD.n12238 VDD.n12236 0.005
R16103 VDD.n10380 VDD.n10379 0.005
R16104 VDD.n10407 VDD.n10406 0.005
R16105 VDD.n12248 VDD.n12247 0.004
R16106 VDD.n12326 VDD.n12325 0.004
R16107 VDD.n12324 VDD.n12248 0.004
R16108 VDD.n12325 VDD.n12324 0.004
R16109 VDD.n84 VDD.n82 0.004
R16110 VDD.n48 VDD.n39 0.004
R16111 VDD.n4896 VDD.n4894 0.004
R16112 VDD.n4880 VDD.n4870 0.004
R16113 VDD.n4665 VDD.n4663 0.004
R16114 VDD.n4649 VDD.n4639 0.004
R16115 VDD.n2789 VDD.n2788 0.004
R16116 VDD.n2810 VDD.n2809 0.004
R16117 VDD.n3114 VDD.n3113 0.004
R16118 VDD.n3131 VDD.n3130 0.004
R16119 VDD.n3352 VDD.n3351 0.004
R16120 VDD.n3369 VDD.n3368 0.004
R16121 VDD.n3589 VDD.n3588 0.004
R16122 VDD.n3606 VDD.n3605 0.004
R16123 VDD.n3827 VDD.n3826 0.004
R16124 VDD.n3844 VDD.n3843 0.004
R16125 VDD.n4064 VDD.n4063 0.004
R16126 VDD.n4081 VDD.n4080 0.004
R16127 VDD.n4302 VDD.n4301 0.004
R16128 VDD.n4319 VDD.n4318 0.004
R16129 VDD.n4625 VDD.n4624 0.004
R16130 VDD.n2926 VDD.n2925 0.004
R16131 VDD.n2925 VDD.n2924 0.004
R16132 VDD.n2921 VDD.n2920 0.004
R16133 VDD.n2924 VDD.n2921 0.004
R16134 VDD.n2923 VDD.n2922 0.004
R16135 VDD.n2924 VDD.n2923 0.004
R16136 VDD.n2919 VDD.n2918 0.004
R16137 VDD.n2924 VDD.n2919 0.004
R16138 VDD.n4549 VDD.n4548 0.004
R16139 VDD.n4548 VDD.n4547 0.004
R16140 VDD.n4544 VDD.n4543 0.004
R16141 VDD.n4547 VDD.n4544 0.004
R16142 VDD.n4546 VDD.n4545 0.004
R16143 VDD.n4547 VDD.n4546 0.004
R16144 VDD.n4542 VDD.n4541 0.004
R16145 VDD.n4547 VDD.n4542 0.004
R16146 VDD.n217 VDD.n216 0.004
R16147 VDD.n227 VDD.n226 0.004
R16148 VDD.n534 VDD.n533 0.004
R16149 VDD.n544 VDD.n543 0.004
R16150 VDD.n768 VDD.n767 0.004
R16151 VDD.n778 VDD.n777 0.004
R16152 VDD.n1001 VDD.n1000 0.004
R16153 VDD.n1011 VDD.n1010 0.004
R16154 VDD.n1235 VDD.n1234 0.004
R16155 VDD.n1245 VDD.n1244 0.004
R16156 VDD.n1468 VDD.n1467 0.004
R16157 VDD.n1478 VDD.n1477 0.004
R16158 VDD.n1702 VDD.n1701 0.004
R16159 VDD.n1712 VDD.n1711 0.004
R16160 VDD.n2020 VDD.n2019 0.004
R16161 VDD.n1949 VDD.n1948 0.004
R16162 VDD.n1956 VDD.n1949 0.004
R16163 VDD.n1954 VDD.n1953 0.004
R16164 VDD.n1951 VDD.n1950 0.004
R16165 VDD.n1958 VDD.n1957 0.004
R16166 VDD.n1957 VDD.n1956 0.004
R16167 VDD.n336 VDD.n335 0.004
R16168 VDD.n343 VDD.n336 0.004
R16169 VDD.n341 VDD.n340 0.004
R16170 VDD.n338 VDD.n337 0.004
R16171 VDD.n345 VDD.n344 0.004
R16172 VDD.n344 VDD.n343 0.004
R16173 VDD.n2045 VDD.n2035 0.004
R16174 VDD.n2061 VDD.n2059 0.004
R16175 VDD.n2276 VDD.n2266 0.004
R16176 VDD.n2292 VDD.n2290 0.004
R16177 VDD.n10299 VDD.n10297 0.004
R16178 VDD.n10285 VDD.n10276 0.004
R16179 VDD.n10181 VDD.n10179 0.004
R16180 VDD.n10167 VDD.n10159 0.004
R16181 VDD.n10099 VDD.n10097 0.004
R16182 VDD.n10084 VDD.n10076 0.004
R16183 VDD.n10054 VDD.n10052 0.004
R16184 VDD.n10040 VDD.n10031 0.004
R16185 VDD.n10646 VDD.n10644 0.004
R16186 VDD.n10632 VDD.n10623 0.004
R16187 VDD.n10527 VDD.n10525 0.004
R16188 VDD.n10513 VDD.n10505 0.004
R16189 VDD.n12104 VDD.n12102 0.004
R16190 VDD.n12072 VDD.n12070 0.004
R16191 VDD.n11337 VDD.n11335 0.004
R16192 VDD.n11303 VDD.n11301 0.004
R16193 VDD.n12315 VDD.n12313 0.004
R16194 VDD.n12279 VDD.n12270 0.004
R16195 VDD.n10370 VDD.n10369 0.004
R16196 VDD.n10397 VDD.n10396 0.004
R16197 VDD.n10369 VDD.n10368 0.004
R16198 VDD.n10396 VDD.n10395 0.004
R16199 VDD.n10432 VDD.n10427 0.004
R16200 VDD.n13 VDD.n1 0.004
R16201 VDD.n12244 VDD.n12232 0.004
R16202 VDD.n10353 VDD.n10352 0.003
R16203 VDD.n93 VDD.n21 0.003
R16204 VDD.n20 VDD.n19 0.003
R16205 VDD.n12323 VDD.n12322 0.003
R16206 VDD.n2576 VDD.n2575 0.003
R16207 VDD.n2743 VDD.n2742 0.003
R16208 VDD.n5377 VDD.n5376 0.003
R16209 VDD.n5528 VDD.n5514 0.003
R16210 VDD.n5527 VDD.n5525 0.003
R16211 VDD.n5608 VDD.n5607 0.003
R16212 VDD.n5629 VDD.n5625 0.003
R16213 VDD.n5643 VDD.n5641 0.003
R16214 VDD.n5649 VDD.n5648 0.003
R16215 VDD.n5660 VDD.n5659 0.003
R16216 VDD.n5406 VDD.n5400 0.003
R16217 VDD.n5416 VDD.n5415 0.003
R16218 VDD.n5451 VDD.n5443 0.003
R16219 VDD.n5461 VDD.n5460 0.003
R16220 VDD.n5558 VDD.n5550 0.003
R16221 VDD.n5565 VDD.n5564 0.003
R16222 VDD.n5668 VDD.n5593 0.003
R16223 VDD.n5738 VDD.n5737 0.003
R16224 VDD.n5889 VDD.n5875 0.003
R16225 VDD.n5888 VDD.n5886 0.003
R16226 VDD.n5969 VDD.n5968 0.003
R16227 VDD.n5990 VDD.n5986 0.003
R16228 VDD.n6004 VDD.n6002 0.003
R16229 VDD.n6010 VDD.n6009 0.003
R16230 VDD.n6021 VDD.n6020 0.003
R16231 VDD.n5767 VDD.n5761 0.003
R16232 VDD.n5777 VDD.n5776 0.003
R16233 VDD.n5812 VDD.n5804 0.003
R16234 VDD.n5822 VDD.n5821 0.003
R16235 VDD.n5919 VDD.n5911 0.003
R16236 VDD.n5926 VDD.n5925 0.003
R16237 VDD.n6029 VDD.n5954 0.003
R16238 VDD.n6100 VDD.n6099 0.003
R16239 VDD.n6251 VDD.n6237 0.003
R16240 VDD.n6250 VDD.n6248 0.003
R16241 VDD.n6331 VDD.n6330 0.003
R16242 VDD.n6352 VDD.n6348 0.003
R16243 VDD.n6366 VDD.n6364 0.003
R16244 VDD.n6372 VDD.n6371 0.003
R16245 VDD.n6383 VDD.n6382 0.003
R16246 VDD.n6129 VDD.n6123 0.003
R16247 VDD.n6139 VDD.n6138 0.003
R16248 VDD.n6174 VDD.n6166 0.003
R16249 VDD.n6184 VDD.n6183 0.003
R16250 VDD.n6281 VDD.n6273 0.003
R16251 VDD.n6288 VDD.n6287 0.003
R16252 VDD.n6391 VDD.n6316 0.003
R16253 VDD.n6462 VDD.n6461 0.003
R16254 VDD.n6613 VDD.n6599 0.003
R16255 VDD.n6612 VDD.n6610 0.003
R16256 VDD.n6693 VDD.n6692 0.003
R16257 VDD.n6714 VDD.n6710 0.003
R16258 VDD.n6728 VDD.n6726 0.003
R16259 VDD.n6734 VDD.n6733 0.003
R16260 VDD.n6745 VDD.n6744 0.003
R16261 VDD.n6491 VDD.n6485 0.003
R16262 VDD.n6501 VDD.n6500 0.003
R16263 VDD.n6536 VDD.n6528 0.003
R16264 VDD.n6546 VDD.n6545 0.003
R16265 VDD.n6643 VDD.n6635 0.003
R16266 VDD.n6650 VDD.n6649 0.003
R16267 VDD.n6753 VDD.n6678 0.003
R16268 VDD.n6824 VDD.n6823 0.003
R16269 VDD.n6975 VDD.n6961 0.003
R16270 VDD.n6974 VDD.n6972 0.003
R16271 VDD.n7055 VDD.n7054 0.003
R16272 VDD.n7076 VDD.n7072 0.003
R16273 VDD.n7090 VDD.n7088 0.003
R16274 VDD.n7096 VDD.n7095 0.003
R16275 VDD.n7107 VDD.n7106 0.003
R16276 VDD.n6853 VDD.n6847 0.003
R16277 VDD.n6863 VDD.n6862 0.003
R16278 VDD.n6898 VDD.n6890 0.003
R16279 VDD.n6908 VDD.n6907 0.003
R16280 VDD.n7005 VDD.n6997 0.003
R16281 VDD.n7012 VDD.n7011 0.003
R16282 VDD.n7115 VDD.n7040 0.003
R16283 VDD.n7186 VDD.n7185 0.003
R16284 VDD.n7337 VDD.n7323 0.003
R16285 VDD.n7336 VDD.n7334 0.003
R16286 VDD.n7417 VDD.n7416 0.003
R16287 VDD.n7438 VDD.n7434 0.003
R16288 VDD.n7452 VDD.n7450 0.003
R16289 VDD.n7458 VDD.n7457 0.003
R16290 VDD.n7469 VDD.n7468 0.003
R16291 VDD.n7215 VDD.n7209 0.003
R16292 VDD.n7225 VDD.n7224 0.003
R16293 VDD.n7260 VDD.n7252 0.003
R16294 VDD.n7270 VDD.n7269 0.003
R16295 VDD.n7367 VDD.n7359 0.003
R16296 VDD.n7374 VDD.n7373 0.003
R16297 VDD.n7477 VDD.n7402 0.003
R16298 VDD.n7548 VDD.n7547 0.003
R16299 VDD.n7699 VDD.n7685 0.003
R16300 VDD.n7698 VDD.n7696 0.003
R16301 VDD.n7779 VDD.n7778 0.003
R16302 VDD.n7800 VDD.n7796 0.003
R16303 VDD.n7814 VDD.n7812 0.003
R16304 VDD.n7820 VDD.n7819 0.003
R16305 VDD.n7831 VDD.n7830 0.003
R16306 VDD.n7577 VDD.n7571 0.003
R16307 VDD.n7587 VDD.n7586 0.003
R16308 VDD.n7622 VDD.n7614 0.003
R16309 VDD.n7632 VDD.n7631 0.003
R16310 VDD.n7729 VDD.n7721 0.003
R16311 VDD.n7736 VDD.n7735 0.003
R16312 VDD.n7839 VDD.n7764 0.003
R16313 VDD.n7910 VDD.n7909 0.003
R16314 VDD.n8061 VDD.n8047 0.003
R16315 VDD.n8060 VDD.n8058 0.003
R16316 VDD.n8141 VDD.n8140 0.003
R16317 VDD.n8162 VDD.n8158 0.003
R16318 VDD.n8176 VDD.n8174 0.003
R16319 VDD.n8182 VDD.n8181 0.003
R16320 VDD.n8193 VDD.n8192 0.003
R16321 VDD.n7939 VDD.n7933 0.003
R16322 VDD.n7949 VDD.n7948 0.003
R16323 VDD.n7984 VDD.n7976 0.003
R16324 VDD.n7994 VDD.n7993 0.003
R16325 VDD.n8091 VDD.n8083 0.003
R16326 VDD.n8098 VDD.n8097 0.003
R16327 VDD.n8201 VDD.n8126 0.003
R16328 VDD.n8272 VDD.n8271 0.003
R16329 VDD.n8423 VDD.n8409 0.003
R16330 VDD.n8422 VDD.n8420 0.003
R16331 VDD.n8503 VDD.n8502 0.003
R16332 VDD.n8524 VDD.n8520 0.003
R16333 VDD.n8538 VDD.n8536 0.003
R16334 VDD.n8544 VDD.n8543 0.003
R16335 VDD.n8555 VDD.n8554 0.003
R16336 VDD.n8301 VDD.n8295 0.003
R16337 VDD.n8311 VDD.n8310 0.003
R16338 VDD.n8346 VDD.n8338 0.003
R16339 VDD.n8356 VDD.n8355 0.003
R16340 VDD.n8453 VDD.n8445 0.003
R16341 VDD.n8460 VDD.n8459 0.003
R16342 VDD.n8563 VDD.n8488 0.003
R16343 VDD.n8634 VDD.n8633 0.003
R16344 VDD.n8785 VDD.n8771 0.003
R16345 VDD.n8784 VDD.n8782 0.003
R16346 VDD.n8865 VDD.n8864 0.003
R16347 VDD.n8886 VDD.n8882 0.003
R16348 VDD.n8900 VDD.n8898 0.003
R16349 VDD.n8906 VDD.n8905 0.003
R16350 VDD.n8917 VDD.n8916 0.003
R16351 VDD.n8663 VDD.n8657 0.003
R16352 VDD.n8673 VDD.n8672 0.003
R16353 VDD.n8708 VDD.n8700 0.003
R16354 VDD.n8718 VDD.n8717 0.003
R16355 VDD.n8815 VDD.n8807 0.003
R16356 VDD.n8822 VDD.n8821 0.003
R16357 VDD.n8925 VDD.n8850 0.003
R16358 VDD.n8996 VDD.n8995 0.003
R16359 VDD.n9147 VDD.n9133 0.003
R16360 VDD.n9146 VDD.n9144 0.003
R16361 VDD.n9227 VDD.n9226 0.003
R16362 VDD.n9248 VDD.n9244 0.003
R16363 VDD.n9262 VDD.n9260 0.003
R16364 VDD.n9268 VDD.n9267 0.003
R16365 VDD.n9279 VDD.n9278 0.003
R16366 VDD.n9025 VDD.n9019 0.003
R16367 VDD.n9035 VDD.n9034 0.003
R16368 VDD.n9070 VDD.n9062 0.003
R16369 VDD.n9080 VDD.n9079 0.003
R16370 VDD.n9177 VDD.n9169 0.003
R16371 VDD.n9184 VDD.n9183 0.003
R16372 VDD.n9287 VDD.n9212 0.003
R16373 VDD.n9358 VDD.n9357 0.003
R16374 VDD.n9509 VDD.n9495 0.003
R16375 VDD.n9508 VDD.n9506 0.003
R16376 VDD.n9589 VDD.n9588 0.003
R16377 VDD.n9610 VDD.n9606 0.003
R16378 VDD.n9624 VDD.n9622 0.003
R16379 VDD.n9630 VDD.n9629 0.003
R16380 VDD.n9641 VDD.n9640 0.003
R16381 VDD.n9387 VDD.n9381 0.003
R16382 VDD.n9397 VDD.n9396 0.003
R16383 VDD.n9432 VDD.n9424 0.003
R16384 VDD.n9442 VDD.n9441 0.003
R16385 VDD.n9539 VDD.n9531 0.003
R16386 VDD.n9546 VDD.n9545 0.003
R16387 VDD.n9649 VDD.n9574 0.003
R16388 VDD.n9720 VDD.n9719 0.003
R16389 VDD.n9871 VDD.n9857 0.003
R16390 VDD.n9870 VDD.n9868 0.003
R16391 VDD.n9951 VDD.n9950 0.003
R16392 VDD.n9972 VDD.n9968 0.003
R16393 VDD.n9986 VDD.n9984 0.003
R16394 VDD.n9992 VDD.n9991 0.003
R16395 VDD.n10003 VDD.n10002 0.003
R16396 VDD.n9749 VDD.n9743 0.003
R16397 VDD.n9759 VDD.n9758 0.003
R16398 VDD.n9794 VDD.n9786 0.003
R16399 VDD.n9804 VDD.n9803 0.003
R16400 VDD.n9901 VDD.n9893 0.003
R16401 VDD.n9908 VDD.n9907 0.003
R16402 VDD.n10011 VDD.n9936 0.003
R16403 VDD.n11940 VDD.n11748 0.003
R16404 VDD.n11183 VDD.n10979 0.003
R16405 VDD.n10956 VDD.n10955 0.003
R16406 VDD.n10949 VDD.n10948 0.003
R16407 VDD.n10947 VDD.n10946 0.003
R16408 VDD.n11026 VDD.n11025 0.003
R16409 VDD.n11036 VDD.n11026 0.003
R16410 VDD.n11139 VDD.n11138 0.003
R16411 VDD.n11137 VDD.n11136 0.003
R16412 VDD.n11105 VDD.n11104 0.003
R16413 VDD.n10859 VDD.n10858 0.003
R16414 VDD.n10842 VDD.n10841 0.003
R16415 VDD.n10840 VDD.n10829 0.003
R16416 VDD.n10824 VDD.n10823 0.003
R16417 VDD.n10823 VDD.n10822 0.003
R16418 VDD.n11725 VDD.n11724 0.003
R16419 VDD.n11715 VDD.n11714 0.003
R16420 VDD.n11713 VDD.n11712 0.003
R16421 VDD.n11793 VDD.n11792 0.003
R16422 VDD.n11803 VDD.n11793 0.003
R16423 VDD.n11898 VDD.n11897 0.003
R16424 VDD.n11886 VDD.n11885 0.003
R16425 VDD.n11879 VDD.n11878 0.003
R16426 VDD.n11640 VDD.n11639 0.003
R16427 VDD.n11621 VDD.n11620 0.003
R16428 VDD.n11619 VDD.n11609 0.003
R16429 VDD.n11604 VDD.n11592 0.003
R16430 VDD.n11592 VDD.n11591 0.003
R16431 VDD.n12211 VDD.n12209 0.003
R16432 VDD.n12175 VDD.n12167 0.003
R16433 VDD.n12007 VDD.n12005 0.003
R16434 VDD.n11971 VDD.n11963 0.003
R16435 VDD.n11439 VDD.n11437 0.003
R16436 VDD.n11405 VDD.n11397 0.003
R16437 VDD.n11241 VDD.n11239 0.003
R16438 VDD.n11207 VDD.n11198 0.003
R16439 VDD.n10366 VDD.n10353 0.003
R16440 VDD.n10393 VDD.n10370 0.003
R16441 VDD.n10420 VDD.n10397 0.003
R16442 VDD.n10446 VDD.n10433 0.003
R16443 VDD.n342 VDD.n341 0.002
R16444 VDD.n339 VDD.n338 0.002
R16445 VDD.n1955 VDD.n1954 0.002
R16446 VDD.n1952 VDD.n1951 0.002
R16447 VDD.n1956 VDD.n1955 0.002
R16448 VDD.n1956 VDD.n1952 0.002
R16449 VDD.n343 VDD.n342 0.002
R16450 VDD.n343 VDD.n339 0.002
R16451 VDD.n10981 VDD.n10980 0.002
R16452 VDD.n11183 VDD.n10981 0.002
R16453 VDD.n11941 VDD.n11940 0.002
R16454 VDD.n11942 VDD.n11941 0.002
R16455 VDD.n19 VDD.n18 0.002
R16456 VDD.n92 VDD.n90 0.002
R16457 VDD.n5002 VDD.n5000 0.002
R16458 VDD.n4996 VDD.n4994 0.002
R16459 VDD.n4771 VDD.n4769 0.002
R16460 VDD.n4765 VDD.n4763 0.002
R16461 VDD.n3002 VDD.n2992 0.002
R16462 VDD.n3015 VDD.n3014 0.002
R16463 VDD.n3239 VDD.n3230 0.002
R16464 VDD.n3252 VDD.n3251 0.002
R16465 VDD.n3477 VDD.n3467 0.002
R16466 VDD.n3490 VDD.n3489 0.002
R16467 VDD.n3714 VDD.n3705 0.002
R16468 VDD.n3727 VDD.n3726 0.002
R16469 VDD.n3952 VDD.n3942 0.002
R16470 VDD.n3965 VDD.n3964 0.002
R16471 VDD.n4189 VDD.n4180 0.002
R16472 VDD.n4202 VDD.n4201 0.002
R16473 VDD.n4427 VDD.n4417 0.002
R16474 VDD.n4440 VDD.n4439 0.002
R16475 VDD.n422 VDD.n409 0.002
R16476 VDD.n435 VDD.n434 0.002
R16477 VDD.n655 VDD.n643 0.002
R16478 VDD.n668 VDD.n667 0.002
R16479 VDD.n889 VDD.n876 0.002
R16480 VDD.n902 VDD.n901 0.002
R16481 VDD.n1122 VDD.n1110 0.002
R16482 VDD.n1135 VDD.n1134 0.002
R16483 VDD.n1356 VDD.n1343 0.002
R16484 VDD.n1369 VDD.n1368 0.002
R16485 VDD.n1589 VDD.n1577 0.002
R16486 VDD.n1602 VDD.n1601 0.002
R16487 VDD.n1823 VDD.n1810 0.002
R16488 VDD.n1836 VDD.n1835 0.002
R16489 VDD.n2161 VDD.n2159 0.002
R16490 VDD.n2167 VDD.n2165 0.002
R16491 VDD.n2392 VDD.n2390 0.002
R16492 VDD.n2398 VDD.n2396 0.002
R16493 VDD.n2596 VDD.n2595 0.002
R16494 VDD.n2600 VDD.n2599 0.002
R16495 VDD.n5151 VDD.n5150 0.002
R16496 VDD.n5147 VDD.n5146 0.002
R16497 VDD.n12092 VDD.n12090 0.002
R16498 VDD.n12084 VDD.n12082 0.002
R16499 VDD.n11323 VDD.n11321 0.002
R16500 VDD.n11315 VDD.n11313 0.002
R16501 VDD.n12322 VDD.n12321 0.002
R16502 VDD.n12252 VDD.n12250 0.002
R16503 VDD.n11184 VDD.n11183 0.002
R16504 VDD.n11185 VDD.n11184 0.002
R16505 VDD.n11940 VDD.n11750 0.002
R16506 VDD.n11750 VDD.n11749 0.002
R16507 VDD.n71 VDD.n69 0.001
R16508 VDD.n60 VDD.n52 0.001
R16509 VDD.n2482 VDD.n2481 0.001
R16510 VDD.n2565 VDD.n2564 0.001
R16511 VDD.n132 VDD.n131 0.001
R16512 VDD.n153 VDD.n152 0.001
R16513 VDD.n5212 VDD.n5211 0.001
R16514 VDD.n5277 VDD.n5276 0.001
R16515 VDD.n2671 VDD.n2670 0.001
R16516 VDD.n2725 VDD.n2724 0.001
R16517 VDD.n2764 VDD.n2759 0.001
R16518 VDD.n5086 VDD.n5085 0.001
R16519 VDD.n158 VDD.n157 0.001
R16520 VDD.n5128 VDD.n5127 0.001
R16521 VDD.n195 VDD.n194 0.001
R16522 VDD.n2594 VDD.n195 0.001
R16523 VDD.n2595 VDD.n2594 0.001
R16524 VDD.n2597 VDD.n2596 0.001
R16525 VDD.n2598 VDD.n2597 0.001
R16526 VDD.n2599 VDD.n2598 0.001
R16527 VDD.n2601 VDD.n2600 0.001
R16528 VDD.n5306 VDD.n2601 0.001
R16529 VDD.n5306 VDD.n5151 0.001
R16530 VDD.n5150 VDD.n5149 0.001
R16531 VDD.n5149 VDD.n5148 0.001
R16532 VDD.n5148 VDD.n5147 0.001
R16533 VDD.n5146 VDD.n5145 0.001
R16534 VDD.n5145 VDD.n5144 0.001
R16535 VDD.n5144 VDD.n5130 0.001
R16536 VDD.n5360 VDD.n5359 0.001
R16537 VDD.n5358 VDD.n5356 0.001
R16538 VDD.n5352 VDD.n5351 0.001
R16539 VDD.n5347 VDD.n5346 0.001
R16540 VDD.n5471 VDD.n5469 0.001
R16541 VDD.n5476 VDD.n5473 0.001
R16542 VDD.n5484 VDD.n5482 0.001
R16543 VDD.n5488 VDD.n5485 0.001
R16544 VDD.n5489 VDD.n5488 0.001
R16545 VDD.n5491 VDD.n5490 0.001
R16546 VDD.n5499 VDD.n5498 0.001
R16547 VDD.n5508 VDD.n5504 0.001
R16548 VDD.n5637 VDD.n5634 0.001
R16549 VDD.n5639 VDD.n5638 0.001
R16550 VDD.n5404 VDD.n5403 0.001
R16551 VDD.n5410 VDD.n5409 0.001
R16552 VDD.n5440 VDD.n5439 0.001
R16553 VDD.n5445 VDD.n5444 0.001
R16554 VDD.n5450 VDD.n5449 0.001
R16555 VDD.n5459 VDD.n5458 0.001
R16556 VDD.n5569 VDD.n5568 0.001
R16557 VDD.n5571 VDD.n5570 0.001
R16558 VDD.n5588 VDD.n5587 0.001
R16559 VDD.n5721 VDD.n5720 0.001
R16560 VDD.n5719 VDD.n5717 0.001
R16561 VDD.n5713 VDD.n5712 0.001
R16562 VDD.n5708 VDD.n5707 0.001
R16563 VDD.n5832 VDD.n5830 0.001
R16564 VDD.n5837 VDD.n5834 0.001
R16565 VDD.n5845 VDD.n5843 0.001
R16566 VDD.n5849 VDD.n5846 0.001
R16567 VDD.n5850 VDD.n5849 0.001
R16568 VDD.n5852 VDD.n5851 0.001
R16569 VDD.n5860 VDD.n5859 0.001
R16570 VDD.n5869 VDD.n5865 0.001
R16571 VDD.n5998 VDD.n5995 0.001
R16572 VDD.n6000 VDD.n5999 0.001
R16573 VDD.n5765 VDD.n5764 0.001
R16574 VDD.n5771 VDD.n5770 0.001
R16575 VDD.n5801 VDD.n5800 0.001
R16576 VDD.n5806 VDD.n5805 0.001
R16577 VDD.n5811 VDD.n5810 0.001
R16578 VDD.n5820 VDD.n5819 0.001
R16579 VDD.n5930 VDD.n5929 0.001
R16580 VDD.n5932 VDD.n5931 0.001
R16581 VDD.n5949 VDD.n5948 0.001
R16582 VDD.n6083 VDD.n6082 0.001
R16583 VDD.n6081 VDD.n6079 0.001
R16584 VDD.n6075 VDD.n6074 0.001
R16585 VDD.n6070 VDD.n6069 0.001
R16586 VDD.n6194 VDD.n6192 0.001
R16587 VDD.n6199 VDD.n6196 0.001
R16588 VDD.n6207 VDD.n6205 0.001
R16589 VDD.n6211 VDD.n6208 0.001
R16590 VDD.n6212 VDD.n6211 0.001
R16591 VDD.n6214 VDD.n6213 0.001
R16592 VDD.n6222 VDD.n6221 0.001
R16593 VDD.n6231 VDD.n6227 0.001
R16594 VDD.n6360 VDD.n6357 0.001
R16595 VDD.n6362 VDD.n6361 0.001
R16596 VDD.n6127 VDD.n6126 0.001
R16597 VDD.n6133 VDD.n6132 0.001
R16598 VDD.n6163 VDD.n6162 0.001
R16599 VDD.n6168 VDD.n6167 0.001
R16600 VDD.n6173 VDD.n6172 0.001
R16601 VDD.n6182 VDD.n6181 0.001
R16602 VDD.n6292 VDD.n6291 0.001
R16603 VDD.n6294 VDD.n6293 0.001
R16604 VDD.n6311 VDD.n6310 0.001
R16605 VDD.n6445 VDD.n6444 0.001
R16606 VDD.n6443 VDD.n6441 0.001
R16607 VDD.n6437 VDD.n6436 0.001
R16608 VDD.n6432 VDD.n6431 0.001
R16609 VDD.n6556 VDD.n6554 0.001
R16610 VDD.n6561 VDD.n6558 0.001
R16611 VDD.n6569 VDD.n6567 0.001
R16612 VDD.n6573 VDD.n6570 0.001
R16613 VDD.n6574 VDD.n6573 0.001
R16614 VDD.n6576 VDD.n6575 0.001
R16615 VDD.n6584 VDD.n6583 0.001
R16616 VDD.n6593 VDD.n6589 0.001
R16617 VDD.n6722 VDD.n6719 0.001
R16618 VDD.n6724 VDD.n6723 0.001
R16619 VDD.n6489 VDD.n6488 0.001
R16620 VDD.n6495 VDD.n6494 0.001
R16621 VDD.n6525 VDD.n6524 0.001
R16622 VDD.n6530 VDD.n6529 0.001
R16623 VDD.n6535 VDD.n6534 0.001
R16624 VDD.n6544 VDD.n6543 0.001
R16625 VDD.n6654 VDD.n6653 0.001
R16626 VDD.n6656 VDD.n6655 0.001
R16627 VDD.n6673 VDD.n6672 0.001
R16628 VDD.n6807 VDD.n6806 0.001
R16629 VDD.n6805 VDD.n6803 0.001
R16630 VDD.n6799 VDD.n6798 0.001
R16631 VDD.n6794 VDD.n6793 0.001
R16632 VDD.n6918 VDD.n6916 0.001
R16633 VDD.n6923 VDD.n6920 0.001
R16634 VDD.n6931 VDD.n6929 0.001
R16635 VDD.n6935 VDD.n6932 0.001
R16636 VDD.n6936 VDD.n6935 0.001
R16637 VDD.n6938 VDD.n6937 0.001
R16638 VDD.n6946 VDD.n6945 0.001
R16639 VDD.n6955 VDD.n6951 0.001
R16640 VDD.n7084 VDD.n7081 0.001
R16641 VDD.n7086 VDD.n7085 0.001
R16642 VDD.n6851 VDD.n6850 0.001
R16643 VDD.n6857 VDD.n6856 0.001
R16644 VDD.n6887 VDD.n6886 0.001
R16645 VDD.n6892 VDD.n6891 0.001
R16646 VDD.n6897 VDD.n6896 0.001
R16647 VDD.n6906 VDD.n6905 0.001
R16648 VDD.n7016 VDD.n7015 0.001
R16649 VDD.n7018 VDD.n7017 0.001
R16650 VDD.n7035 VDD.n7034 0.001
R16651 VDD.n7169 VDD.n7168 0.001
R16652 VDD.n7167 VDD.n7165 0.001
R16653 VDD.n7161 VDD.n7160 0.001
R16654 VDD.n7156 VDD.n7155 0.001
R16655 VDD.n7280 VDD.n7278 0.001
R16656 VDD.n7285 VDD.n7282 0.001
R16657 VDD.n7293 VDD.n7291 0.001
R16658 VDD.n7297 VDD.n7294 0.001
R16659 VDD.n7298 VDD.n7297 0.001
R16660 VDD.n7300 VDD.n7299 0.001
R16661 VDD.n7308 VDD.n7307 0.001
R16662 VDD.n7317 VDD.n7313 0.001
R16663 VDD.n7446 VDD.n7443 0.001
R16664 VDD.n7448 VDD.n7447 0.001
R16665 VDD.n7213 VDD.n7212 0.001
R16666 VDD.n7219 VDD.n7218 0.001
R16667 VDD.n7249 VDD.n7248 0.001
R16668 VDD.n7254 VDD.n7253 0.001
R16669 VDD.n7259 VDD.n7258 0.001
R16670 VDD.n7268 VDD.n7267 0.001
R16671 VDD.n7378 VDD.n7377 0.001
R16672 VDD.n7380 VDD.n7379 0.001
R16673 VDD.n7397 VDD.n7396 0.001
R16674 VDD.n7531 VDD.n7530 0.001
R16675 VDD.n7529 VDD.n7527 0.001
R16676 VDD.n7523 VDD.n7522 0.001
R16677 VDD.n7518 VDD.n7517 0.001
R16678 VDD.n7642 VDD.n7640 0.001
R16679 VDD.n7647 VDD.n7644 0.001
R16680 VDD.n7655 VDD.n7653 0.001
R16681 VDD.n7659 VDD.n7656 0.001
R16682 VDD.n7660 VDD.n7659 0.001
R16683 VDD.n7662 VDD.n7661 0.001
R16684 VDD.n7670 VDD.n7669 0.001
R16685 VDD.n7679 VDD.n7675 0.001
R16686 VDD.n7808 VDD.n7805 0.001
R16687 VDD.n7810 VDD.n7809 0.001
R16688 VDD.n7575 VDD.n7574 0.001
R16689 VDD.n7581 VDD.n7580 0.001
R16690 VDD.n7611 VDD.n7610 0.001
R16691 VDD.n7616 VDD.n7615 0.001
R16692 VDD.n7621 VDD.n7620 0.001
R16693 VDD.n7630 VDD.n7629 0.001
R16694 VDD.n7740 VDD.n7739 0.001
R16695 VDD.n7742 VDD.n7741 0.001
R16696 VDD.n7759 VDD.n7758 0.001
R16697 VDD.n7893 VDD.n7892 0.001
R16698 VDD.n7891 VDD.n7889 0.001
R16699 VDD.n7885 VDD.n7884 0.001
R16700 VDD.n7880 VDD.n7879 0.001
R16701 VDD.n8004 VDD.n8002 0.001
R16702 VDD.n8009 VDD.n8006 0.001
R16703 VDD.n8017 VDD.n8015 0.001
R16704 VDD.n8021 VDD.n8018 0.001
R16705 VDD.n8022 VDD.n8021 0.001
R16706 VDD.n8024 VDD.n8023 0.001
R16707 VDD.n8032 VDD.n8031 0.001
R16708 VDD.n8041 VDD.n8037 0.001
R16709 VDD.n8170 VDD.n8167 0.001
R16710 VDD.n8172 VDD.n8171 0.001
R16711 VDD.n7937 VDD.n7936 0.001
R16712 VDD.n7943 VDD.n7942 0.001
R16713 VDD.n7973 VDD.n7972 0.001
R16714 VDD.n7978 VDD.n7977 0.001
R16715 VDD.n7983 VDD.n7982 0.001
R16716 VDD.n7992 VDD.n7991 0.001
R16717 VDD.n8102 VDD.n8101 0.001
R16718 VDD.n8104 VDD.n8103 0.001
R16719 VDD.n8121 VDD.n8120 0.001
R16720 VDD.n8255 VDD.n8254 0.001
R16721 VDD.n8253 VDD.n8251 0.001
R16722 VDD.n8247 VDD.n8246 0.001
R16723 VDD.n8242 VDD.n8241 0.001
R16724 VDD.n8366 VDD.n8364 0.001
R16725 VDD.n8371 VDD.n8368 0.001
R16726 VDD.n8379 VDD.n8377 0.001
R16727 VDD.n8383 VDD.n8380 0.001
R16728 VDD.n8384 VDD.n8383 0.001
R16729 VDD.n8386 VDD.n8385 0.001
R16730 VDD.n8394 VDD.n8393 0.001
R16731 VDD.n8403 VDD.n8399 0.001
R16732 VDD.n8532 VDD.n8529 0.001
R16733 VDD.n8534 VDD.n8533 0.001
R16734 VDD.n8299 VDD.n8298 0.001
R16735 VDD.n8305 VDD.n8304 0.001
R16736 VDD.n8335 VDD.n8334 0.001
R16737 VDD.n8340 VDD.n8339 0.001
R16738 VDD.n8345 VDD.n8344 0.001
R16739 VDD.n8354 VDD.n8353 0.001
R16740 VDD.n8464 VDD.n8463 0.001
R16741 VDD.n8466 VDD.n8465 0.001
R16742 VDD.n8483 VDD.n8482 0.001
R16743 VDD.n8617 VDD.n8616 0.001
R16744 VDD.n8615 VDD.n8613 0.001
R16745 VDD.n8609 VDD.n8608 0.001
R16746 VDD.n8604 VDD.n8603 0.001
R16747 VDD.n8728 VDD.n8726 0.001
R16748 VDD.n8733 VDD.n8730 0.001
R16749 VDD.n8741 VDD.n8739 0.001
R16750 VDD.n8745 VDD.n8742 0.001
R16751 VDD.n8746 VDD.n8745 0.001
R16752 VDD.n8748 VDD.n8747 0.001
R16753 VDD.n8756 VDD.n8755 0.001
R16754 VDD.n8765 VDD.n8761 0.001
R16755 VDD.n8894 VDD.n8891 0.001
R16756 VDD.n8896 VDD.n8895 0.001
R16757 VDD.n8661 VDD.n8660 0.001
R16758 VDD.n8667 VDD.n8666 0.001
R16759 VDD.n8697 VDD.n8696 0.001
R16760 VDD.n8702 VDD.n8701 0.001
R16761 VDD.n8707 VDD.n8706 0.001
R16762 VDD.n8716 VDD.n8715 0.001
R16763 VDD.n8826 VDD.n8825 0.001
R16764 VDD.n8828 VDD.n8827 0.001
R16765 VDD.n8845 VDD.n8844 0.001
R16766 VDD.n8979 VDD.n8978 0.001
R16767 VDD.n8977 VDD.n8975 0.001
R16768 VDD.n8971 VDD.n8970 0.001
R16769 VDD.n8966 VDD.n8965 0.001
R16770 VDD.n9090 VDD.n9088 0.001
R16771 VDD.n9095 VDD.n9092 0.001
R16772 VDD.n9103 VDD.n9101 0.001
R16773 VDD.n9107 VDD.n9104 0.001
R16774 VDD.n9108 VDD.n9107 0.001
R16775 VDD.n9110 VDD.n9109 0.001
R16776 VDD.n9118 VDD.n9117 0.001
R16777 VDD.n9127 VDD.n9123 0.001
R16778 VDD.n9256 VDD.n9253 0.001
R16779 VDD.n9258 VDD.n9257 0.001
R16780 VDD.n9023 VDD.n9022 0.001
R16781 VDD.n9029 VDD.n9028 0.001
R16782 VDD.n9059 VDD.n9058 0.001
R16783 VDD.n9064 VDD.n9063 0.001
R16784 VDD.n9069 VDD.n9068 0.001
R16785 VDD.n9078 VDD.n9077 0.001
R16786 VDD.n9188 VDD.n9187 0.001
R16787 VDD.n9190 VDD.n9189 0.001
R16788 VDD.n9207 VDD.n9206 0.001
R16789 VDD.n9341 VDD.n9340 0.001
R16790 VDD.n9339 VDD.n9337 0.001
R16791 VDD.n9333 VDD.n9332 0.001
R16792 VDD.n9328 VDD.n9327 0.001
R16793 VDD.n9452 VDD.n9450 0.001
R16794 VDD.n9457 VDD.n9454 0.001
R16795 VDD.n9465 VDD.n9463 0.001
R16796 VDD.n9469 VDD.n9466 0.001
R16797 VDD.n9470 VDD.n9469 0.001
R16798 VDD.n9472 VDD.n9471 0.001
R16799 VDD.n9480 VDD.n9479 0.001
R16800 VDD.n9489 VDD.n9485 0.001
R16801 VDD.n9618 VDD.n9615 0.001
R16802 VDD.n9620 VDD.n9619 0.001
R16803 VDD.n9385 VDD.n9384 0.001
R16804 VDD.n9391 VDD.n9390 0.001
R16805 VDD.n9421 VDD.n9420 0.001
R16806 VDD.n9426 VDD.n9425 0.001
R16807 VDD.n9431 VDD.n9430 0.001
R16808 VDD.n9440 VDD.n9439 0.001
R16809 VDD.n9550 VDD.n9549 0.001
R16810 VDD.n9552 VDD.n9551 0.001
R16811 VDD.n9569 VDD.n9568 0.001
R16812 VDD.n9703 VDD.n9702 0.001
R16813 VDD.n9701 VDD.n9699 0.001
R16814 VDD.n9695 VDD.n9694 0.001
R16815 VDD.n9690 VDD.n9689 0.001
R16816 VDD.n9814 VDD.n9812 0.001
R16817 VDD.n9819 VDD.n9816 0.001
R16818 VDD.n9827 VDD.n9825 0.001
R16819 VDD.n9831 VDD.n9828 0.001
R16820 VDD.n9832 VDD.n9831 0.001
R16821 VDD.n9834 VDD.n9833 0.001
R16822 VDD.n9842 VDD.n9841 0.001
R16823 VDD.n9851 VDD.n9847 0.001
R16824 VDD.n9980 VDD.n9977 0.001
R16825 VDD.n9982 VDD.n9981 0.001
R16826 VDD.n9747 VDD.n9746 0.001
R16827 VDD.n9753 VDD.n9752 0.001
R16828 VDD.n9783 VDD.n9782 0.001
R16829 VDD.n9788 VDD.n9787 0.001
R16830 VDD.n9793 VDD.n9792 0.001
R16831 VDD.n9802 VDD.n9801 0.001
R16832 VDD.n9912 VDD.n9911 0.001
R16833 VDD.n9914 VDD.n9913 0.001
R16834 VDD.n9931 VDD.n9930 0.001
R16835 VDD.n11069 VDD.n11058 0.001
R16836 VDD.n11071 VDD.n11070 0.001
R16837 VDD.n11074 VDD.n11073 0.001
R16838 VDD.n11000 VDD.n10999 0.001
R16839 VDD.n10998 VDD.n10997 0.001
R16840 VDD.n11155 VDD.n11154 0.001
R16841 VDD.n11167 VDD.n11166 0.001
R16842 VDD.n11181 VDD.n11180 0.001
R16843 VDD.n11153 VDD.n11152 0.001
R16844 VDD.n10744 VDD.n10733 0.001
R16845 VDD.n10746 VDD.n10745 0.001
R16846 VDD.n10760 VDD.n10759 0.001
R16847 VDD.n10762 VDD.n10761 0.001
R16848 VDD.n11835 VDD.n11824 0.001
R16849 VDD.n11837 VDD.n11836 0.001
R16850 VDD.n11842 VDD.n11841 0.001
R16851 VDD.n11768 VDD.n11767 0.001
R16852 VDD.n11766 VDD.n11765 0.001
R16853 VDD.n11913 VDD.n11912 0.001
R16854 VDD.n11925 VDD.n11924 0.001
R16855 VDD.n11938 VDD.n11937 0.001
R16856 VDD.n11911 VDD.n11910 0.001
R16857 VDD.n11515 VDD.n11504 0.001
R16858 VDD.n11517 VDD.n11516 0.001
R16859 VDD.n11530 VDD.n11529 0.001
R16860 VDD.n11532 VDD.n11531 0.001
R16861 VDD.n12199 VDD.n12197 0.001
R16862 VDD.n12188 VDD.n12179 0.001
R16863 VDD.n11995 VDD.n11993 0.001
R16864 VDD.n11984 VDD.n11975 0.001
R16865 VDD.n11427 VDD.n11425 0.001
R16866 VDD.n11417 VDD.n11409 0.001
R16867 VDD.n11229 VDD.n11227 0.001
R16868 VDD.n11219 VDD.n11211 0.001
R16869 VDD.n12302 VDD.n12300 0.001
R16870 VDD.n12291 VDD.n12283 0.001
R16871 VBN.n12 VBN.t12 234.071
R16872 VBN.n12 VBN.t17 233.984
R16873 VBN.n250 VBN.n249 175.251
R16874 VBN.n173 VBN.n172 175.251
R16875 VBN.n80 VBN.n79 175.251
R16876 VBN.n249 VBN.t0 122.709
R16877 VBN.n172 VBN.t1 122.709
R16878 VBN.n79 VBN.t2 122.709
R16879 VBN.n0 VBN.t16 117.49
R16880 VBN.n10 VBN.t3 117.249
R16881 VBN.n8 VBN.t4 117.249
R16882 VBN.n6 VBN.t7 117.249
R16883 VBN.n4 VBN.t9 117.249
R16884 VBN.n2 VBN.t10 117.249
R16885 VBN.n0 VBN.t13 117.249
R16886 VBN.n1 VBN.t15 117.247
R16887 VBN.n3 VBN.t14 117.247
R16888 VBN.n5 VBN.t11 117.247
R16889 VBN.n7 VBN.t8 117.247
R16890 VBN.n9 VBN.t6 117.247
R16891 VBN.n11 VBN.t5 117.247
R16892 VBN.n57 VBN.n56 9.3
R16893 VBN.n233 VBN.n232 9.013
R16894 VBN.n193 VBN.n192 9.013
R16895 VBN.n107 VBN.n106 9.013
R16896 VBN.n223 VBN.n222 9.013
R16897 VBN.n92 VBN.n91 9.013
R16898 VBN.n28 VBN.n27 9.013
R16899 VBN.n13 VBN.n12 8.779
R16900 VBN.n251 VBN.n250 6.413
R16901 VBN.n174 VBN.n173 6.413
R16902 VBN.n81 VBN.n80 6.413
R16903 VBN.n177 VBN.n176 4.5
R16904 VBN.n159 VBN.n149 4.5
R16905 VBN.n164 VBN.n145 4.5
R16906 VBN.n161 VBN.n147 4.5
R16907 VBN.n156 VBN.n153 4.5
R16908 VBN.n214 VBN.n212 4.5
R16909 VBN.n86 VBN.n83 4.5
R16910 VBN.n43 VBN.n42 4.5
R16911 VBN.n34 VBN.n33 4.5
R16912 VBN.n39 VBN.n38 4.5
R16913 VBN.n49 VBN.n48 4.5
R16914 VBN.n60 VBN.n59 4.5
R16915 VBN.n254 VBN.n253 4.5
R16916 VBN.n139 VBN.n136 4.5
R16917 VBN.n264 VBN.n263 4.5
R16918 VBN.n281 VBN.n279 4.5
R16919 VBN.n133 VBN.n130 4.5
R16920 VBN.n122 VBN.n119 4.5
R16921 VBN.n108 VBN.n107 3.992
R16922 VBN.n224 VBN.n223 3.992
R16923 VBN.n234 VBN.n233 3.882
R16924 VBN.n93 VBN.n92 3.882
R16925 VBN.n64 VBN.n28 2.792
R16926 VBN.n250 VBN.n248 2.787
R16927 VBN.n173 VBN.n171 2.787
R16928 VBN.n194 VBN.n193 2.738
R16929 VBN.n251 VBN.n247 2.695
R16930 VBN.n174 VBN.n170 2.695
R16931 VBN.n57 VBN.n55 2.695
R16932 VBN.n279 VBN.n278 2.656
R16933 VBN.n26 VBN.n25 2.535
R16934 VBN.n191 VBN.n190 2.415
R16935 VBN.n262 VBN.n261 2.082
R16936 VBN.n129 VBN.n128 2.082
R16937 VBN.n252 VBN.n251 2.082
R16938 VBN.n118 VBN.n117 2.082
R16939 VBN.n144 VBN.n143 2.082
R16940 VBN.n152 VBN.n151 2.082
R16941 VBN.n175 VBN.n174 2.082
R16942 VBN.n211 VBN.n210 2.082
R16943 VBN.n82 VBN.n81 2.082
R16944 VBN.n32 VBN.n31 2.082
R16945 VBN.n47 VBN.n46 2.082
R16946 VBN.n58 VBN.n57 2.082
R16947 VBN.n288 VBN.n287 1.957
R16948 VBN.n282 VBN.n281 1.501
R16949 VBN.n140 VBN.n139 1.501
R16950 VBN.n215 VBN.n214 1.5
R16951 VBN.n226 VBN.n225 1.5
R16952 VBN.n87 VBN.n86 1.5
R16953 VBN.n98 VBN.n97 1.5
R16954 VBN.n265 VBN.n264 1.5
R16955 VBN.n134 VBN.n133 1.5
R16956 VBN.n255 VBN.n254 1.5
R16957 VBN.n123 VBN.n122 1.5
R16958 VBN.n110 VBN.n109 1.5
R16959 VBN.n238 VBN.n237 1.5
R16960 VBN.n252 VBN.n246 1.449
R16961 VBN.n175 VBN.n169 1.449
R16962 VBN.n82 VBN.n78 1.449
R16963 VBN.n233 VBN.n231 1.328
R16964 VBN.n118 VBN.n116 1.328
R16965 VBN.n193 VBN.n191 1.328
R16966 VBN.n211 VBN.n209 1.328
R16967 VBN.n92 VBN.n90 1.328
R16968 VBN.n58 VBN.n54 1.328
R16969 VBN.n279 VBN.n268 1.207
R16970 VBN.n130 VBN.n129 1.207
R16971 VBN.n107 VBN.n105 1.207
R16972 VBN.n147 VBN.n146 1.207
R16973 VBN.n153 VBN.n152 1.207
R16974 VBN.n223 VBN.n221 1.207
R16975 VBN.n38 VBN.n37 1.207
R16976 VBN.n48 VBN.n47 1.207
R16977 VBN.n28 VBN.n26 1.207
R16978 VBN.n286 VBN.n285 1.137
R16979 VBN.n283 VBN.n14 1.137
R16980 VBN.n263 VBN.n262 1.086
R16981 VBN.n136 VBN.n135 1.086
R16982 VBN.n145 VBN.n144 1.086
R16983 VBN.n149 VBN.n148 1.086
R16984 VBN.n33 VBN.n32 1.086
R16985 VBN.n42 VBN.n41 1.086
R16986 VBN.n65 VBN.n64 0.935
R16987 VBN.n195 VBN.n194 0.935
R16988 VBN.n287 VBN.n13 0.884
R16989 VBN.n119 VBN.n118 0.724
R16990 VBN.n212 VBN.n211 0.724
R16991 VBN.n59 VBN.n58 0.724
R16992 VBN.n253 VBN.n252 0.603
R16993 VBN.n176 VBN.n175 0.603
R16994 VBN.n83 VBN.n82 0.603
R16995 VBN.n128 VBN.n127 0.557
R16996 VBN.n151 VBN.n150 0.557
R16997 VBN.n13 VBN.n11 0.51
R16998 VBN VBN.n288 0.333
R16999 VBN.n288 VBN 0.33
R17000 VBN.n100 VBN.n99 0.245
R17001 VBN.n228 VBN.n227 0.245
R17002 VBN.n11 VBN.n10 0.241
R17003 VBN.n10 VBN.n9 0.241
R17004 VBN.n9 VBN.n8 0.241
R17005 VBN.n8 VBN.n7 0.241
R17006 VBN.n7 VBN.n6 0.241
R17007 VBN.n6 VBN.n5 0.241
R17008 VBN.n5 VBN.n4 0.241
R17009 VBN.n4 VBN.n3 0.241
R17010 VBN.n3 VBN.n2 0.241
R17011 VBN.n2 VBN.n1 0.241
R17012 VBN.n1 VBN.n0 0.241
R17013 VBN.n287 VBN.n286 0.14
R17014 VBN.n180 VBN.n179 0.048
R17015 VBN.n167 VBN.n166 0.048
R17016 VBN.n219 VBN.n218 0.048
R17017 VBN.n95 VBN.n94 0.048
R17018 VBN.n52 VBN.n51 0.048
R17019 VBN.n63 VBN.n62 0.048
R17020 VBN.n160 VBN.n159 0.044
R17021 VBN.n43 VBN.n40 0.044
R17022 VBN.n281 VBN.n280 0.042
R17023 VBN.n161 VBN.n160 0.042
R17024 VBN.n40 VBN.n39 0.042
R17025 VBN.n264 VBN.n260 0.036
R17026 VBN.n165 VBN.n164 0.036
R17027 VBN.n34 VBN.n30 0.036
R17028 VBN.n133 VBN.n132 0.034
R17029 VBN.n156 VBN.n155 0.034
R17030 VBN.n50 VBN.n49 0.034
R17031 VBN.n194 VBN.n180 0.031
R17032 VBN.n64 VBN.n63 0.031
R17033 VBN.n254 VBN.n243 0.028
R17034 VBN.n178 VBN.n177 0.028
R17035 VBN.n86 VBN.n77 0.028
R17036 VBN.n122 VBN.n121 0.026
R17037 VBN.n214 VBN.n213 0.026
R17038 VBN.n198 VBN.n197 0.026
R17039 VBN.n215 VBN.n206 0.026
R17040 VBN.n226 VBN.n217 0.026
R17041 VBN.n61 VBN.n60 0.026
R17042 VBN.n98 VBN.n89 0.026
R17043 VBN.n87 VBN.n76 0.026
R17044 VBN.n68 VBN.n67 0.026
R17045 VBN.n245 VBN.n244 0.023
R17046 VBN.n121 VBN.n120 0.023
R17047 VBN.n168 VBN.n167 0.023
R17048 VBN.n85 VBN.n84 0.023
R17049 VBN.n62 VBN.n61 0.023
R17050 VBN.n236 VBN.n235 0.021
R17051 VBN.n243 VBN.n242 0.021
R17052 VBN.n115 VBN.n114 0.021
R17053 VBN.n179 VBN.n178 0.021
R17054 VBN.n208 VBN.n207 0.021
R17055 VBN.n96 VBN.n95 0.021
R17056 VBN.n53 VBN.n52 0.021
R17057 VBN.n281 VBN.n267 0.019
R17058 VBN.n104 VBN.n103 0.019
R17059 VBN.n162 VBN.n161 0.019
R17060 VBN.n157 VBN.n156 0.019
R17061 VBN.n220 VBN.n219 0.019
R17062 VBN.n39 VBN.n36 0.019
R17063 VBN.n49 VBN.n45 0.019
R17064 VBN.n139 VBN.n138 0.017
R17065 VBN.n164 VBN.n163 0.017
R17066 VBN.n159 VBN.n158 0.017
R17067 VBN.n35 VBN.n34 0.017
R17068 VBN.n44 VBN.n43 0.017
R17069 VBN.n132 VBN.n131 0.015
R17070 VBN.n155 VBN.n154 0.015
R17071 VBN.n51 VBN.n50 0.015
R17072 VBN.n257 VBN.n256 0.015
R17073 VBN.n101 VBN.n100 0.015
R17074 VBN.n229 VBN.n228 0.015
R17075 VBN.n201 VBN.n200 0.014
R17076 VBN.n202 VBN.n201 0.014
R17077 VBN.n203 VBN.n202 0.014
R17078 VBN.n204 VBN.n203 0.014
R17079 VBN.n74 VBN.n73 0.014
R17080 VBN.n73 VBN.n72 0.014
R17081 VBN.n72 VBN.n71 0.014
R17082 VBN.n71 VBN.n70 0.014
R17083 VBN.n125 VBN.n124 0.014
R17084 VBN.n140 VBN.n134 0.013
R17085 VBN.n282 VBN.n265 0.013
R17086 VBN.n283 VBN.n140 0.013
R17087 VBN.n283 VBN.n282 0.013
R17088 VBN.n260 VBN.n259 0.013
R17089 VBN.n109 VBN.n104 0.013
R17090 VBN.n166 VBN.n165 0.013
R17091 VBN.n225 VBN.n220 0.013
R17092 VBN.n30 VBN.n29 0.013
R17093 VBN.n111 VBN.n110 0.013
R17094 VBN.n200 VBN.n199 0.012
R17095 VBN.n75 VBN.n74 0.012
R17096 VBN.n239 VBN.n238 0.012
R17097 VBN.n240 VBN.n239 0.012
R17098 VBN.n112 VBN.n111 0.012
R17099 VBN.n99 VBN.n98 0.012
R17100 VBN.n227 VBN.n226 0.011
R17101 VBN.n237 VBN.n236 0.011
R17102 VBN.n122 VBN.n115 0.011
R17103 VBN.n214 VBN.n208 0.011
R17104 VBN.n205 VBN.n204 0.011
R17105 VBN.n97 VBN.n96 0.011
R17106 VBN.n60 VBN.n53 0.011
R17107 VBN.n70 VBN.n69 0.011
R17108 VBN.n265 VBN.n258 0.011
R17109 VBN.n256 VBN.n255 0.01
R17110 VBN.n134 VBN.n126 0.01
R17111 VBN.n124 VBN.n123 0.01
R17112 VBN.n254 VBN.n245 0.009
R17113 VBN.n177 VBN.n168 0.009
R17114 VBN.n197 VBN.n196 0.009
R17115 VBN.n86 VBN.n85 0.009
R17116 VBN.n88 VBN.n87 0.009
R17117 VBN.n255 VBN.n241 0.009
R17118 VBN.n216 VBN.n215 0.008
R17119 VBN.n67 VBN.n66 0.008
R17120 VBN.n123 VBN.n113 0.008
R17121 VBN.n267 VBN.n266 0.007
R17122 VBN.n138 VBN.n137 0.007
R17123 VBN.n163 VBN.n162 0.007
R17124 VBN.n158 VBN.n157 0.007
R17125 VBN.n196 VBN.n195 0.007
R17126 VBN.n217 VBN.n216 0.007
R17127 VBN.n36 VBN.n35 0.007
R17128 VBN.n45 VBN.n44 0.007
R17129 VBN.n89 VBN.n88 0.007
R17130 VBN.n66 VBN.n65 0.007
R17131 VBN.n113 VBN.n112 0.007
R17132 VBN.n97 VBN.n93 0.007
R17133 VBN.n237 VBN.n234 0.007
R17134 VBN.n109 VBN.n108 0.006
R17135 VBN.n225 VBN.n224 0.006
R17136 VBN.n238 VBN.n230 0.006
R17137 VBN.n241 VBN.n240 0.006
R17138 VBN.n110 VBN.n102 0.006
R17139 VBN.n206 VBN.n205 0.005
R17140 VBN.n69 VBN.n68 0.005
R17141 VBN.n230 VBN.n229 0.004
R17142 VBN.n102 VBN.n101 0.004
R17143 VBN.n270 VBN.n269 0.004
R17144 VBN.n278 VBN.n270 0.004
R17145 VBN.n274 VBN.n273 0.004
R17146 VBN.n278 VBN.n274 0.004
R17147 VBN.n272 VBN.n271 0.004
R17148 VBN.n278 VBN.n272 0.004
R17149 VBN.n276 VBN.n275 0.004
R17150 VBN.n190 VBN.n189 0.004
R17151 VBN.n189 VBN.n188 0.004
R17152 VBN.n184 VBN.n183 0.004
R17153 VBN.n188 VBN.n184 0.004
R17154 VBN.n182 VBN.n181 0.004
R17155 VBN.n188 VBN.n182 0.004
R17156 VBN.n186 VBN.n185 0.004
R17157 VBN.n199 VBN.n198 0.004
R17158 VBN.n25 VBN.n24 0.004
R17159 VBN.n24 VBN.n23 0.004
R17160 VBN.n16 VBN.n15 0.004
R17161 VBN.n19 VBN.n18 0.004
R17162 VBN.n22 VBN.n21 0.004
R17163 VBN.n23 VBN.n22 0.004
R17164 VBN.n76 VBN.n75 0.004
R17165 VBN.n258 VBN.n257 0.004
R17166 VBN.n126 VBN.n125 0.004
R17167 VBN.n277 VBN.n276 0.002
R17168 VBN.n278 VBN.n277 0.002
R17169 VBN.n187 VBN.n186 0.002
R17170 VBN.n188 VBN.n187 0.002
R17171 VBN.n20 VBN.n19 0.002
R17172 VBN.n17 VBN.n16 0.002
R17173 VBN.n23 VBN.n17 0.002
R17174 VBN.n23 VBN.n20 0.002
R17175 VBN.n284 VBN.n283 0.002
R17176 VBN.n142 VBN.n141 0.002
R17177 VBN.n283 VBN.n142 0.002
R17178 VBN.n286 VBN.n284 0.002
R17179 p_bais.n12 p_bais.t19 308.184
R17180 p_bais.n0 p_bais.t7 308.183
R17181 p_bais.n4 p_bais.t16 307.987
R17182 p_bais.n16 p_bais.t18 307.987
R17183 p_bais.n14 p_bais.t20 307.987
R17184 p_bais.n12 p_bais.t21 307.987
R17185 p_bais.n3 p_bais.t9 307.986
R17186 p_bais.n2 p_bais.t13 307.986
R17187 p_bais.n1 p_bais.t8 307.986
R17188 p_bais.n0 p_bais.t10 307.986
R17189 p_bais.n15 p_bais.t15 307.986
R17190 p_bais.n13 p_bais.t17 307.986
R17191 p_bais.n7 p_bais.t11 307.161
R17192 p_bais.n100 p_bais.t6 200.105
R17193 p_bais.n51 p_bais.t5 199.973
R17194 p_bais.n49 p_bais.t12 199.786
R17195 p_bais.n104 p_bais.t14 199.786
R17196 p_bais.n357 p_bais.n356 175.251
R17197 p_bais.n293 p_bais.n292 175.251
R17198 p_bais.n144 p_bais.n143 175.251
R17199 p_bais.n356 p_bais.t2 122.709
R17200 p_bais.n292 p_bais.t4 122.709
R17201 p_bais.n143 p_bais.t3 122.709
R17202 p_bais.n923 p_bais.n922 13.176
R17203 p_bais.n562 p_bais.n561 13.176
R17204 p_bais.n957 p_bais.n956 9.3
R17205 p_bais.n1083 p_bais.n1082 9.3
R17206 p_bais.n1086 p_bais.n1085 9.3
R17207 p_bais.n1094 p_bais.n1093 9.3
R17208 p_bais.n1133 p_bais.n1132 9.3
R17209 p_bais.n1144 p_bais.n1143 9.3
R17210 p_bais.n1135 p_bais.n1134 9.3
R17211 p_bais.n1123 p_bais.n1122 9.3
R17212 p_bais.n1125 p_bais.n1124 9.3
R17213 p_bais.n1097 p_bais.n1096 9.3
R17214 p_bais.n1073 p_bais.n1072 9.3
R17215 p_bais.n928 p_bais.n927 9.3
R17216 p_bais.n959 p_bais.n958 9.3
R17217 p_bais.n844 p_bais.n843 9.3
R17218 p_bais.n832 p_bais.n831 9.3
R17219 p_bais.n830 p_bais.n829 9.3
R17220 p_bais.n596 p_bais.n595 9.3
R17221 p_bais.n722 p_bais.n721 9.3
R17222 p_bais.n725 p_bais.n724 9.3
R17223 p_bais.n733 p_bais.n732 9.3
R17224 p_bais.n772 p_bais.n771 9.3
R17225 p_bais.n783 p_bais.n782 9.3
R17226 p_bais.n774 p_bais.n773 9.3
R17227 p_bais.n762 p_bais.n761 9.3
R17228 p_bais.n764 p_bais.n763 9.3
R17229 p_bais.n736 p_bais.n735 9.3
R17230 p_bais.n712 p_bais.n711 9.3
R17231 p_bais.n567 p_bais.n566 9.3
R17232 p_bais.n598 p_bais.n597 9.3
R17233 p_bais.n483 p_bais.n482 9.3
R17234 p_bais.n471 p_bais.n470 9.3
R17235 p_bais.n469 p_bais.n468 9.3
R17236 p_bais.n179 p_bais.n178 9.3
R17237 p_bais.n340 p_bais.n339 9.013
R17238 p_bais.n253 p_bais.n252 9.013
R17239 p_bais.n402 p_bais.n401 9.013
R17240 p_bais.n327 p_bais.n326 9.013
R17241 p_bais.n139 p_bais.n138 9.013
R17242 p_bais.n210 p_bais.n209 9.013
R17243 p_bais.n854 p_bais.n853 8.454
R17244 p_bais.n493 p_bais.n492 8.454
R17245 p_bais.n1155 p_bais.n1154 8.454
R17246 p_bais.n794 p_bais.n793 8.454
R17247 p_bais.n358 p_bais.n357 6.413
R17248 p_bais.n294 p_bais.n293 6.413
R17249 p_bais.n145 p_bais.n144 6.413
R17250 p_bais.n1085 p_bais.n1084 5.458
R17251 p_bais.n724 p_bais.n723 5.458
R17252 p_bais.n956 p_bais.n955 5.081
R17253 p_bais.n595 p_bais.n594 5.081
R17254 p_bais.n822 p_bais.n821 4.65
R17255 p_bais.n949 p_bais.n948 4.65
R17256 p_bais.n461 p_bais.n460 4.65
R17257 p_bais.n588 p_bais.n587 4.65
R17258 p_bais.n837 p_bais.n836 4.5
R17259 p_bais.n1113 p_bais.n1112 4.5
R17260 p_bais.n1107 p_bais.n1064 4.5
R17261 p_bais.n1119 p_bais.n1060 4.5
R17262 p_bais.n1129 p_bais.n1128 4.5
R17263 p_bais.n1148 p_bais.n1147 4.5
R17264 p_bais.n1137 p_bais.n1057 4.5
R17265 p_bais.n1103 p_bais.n1102 4.5
R17266 p_bais.n1090 p_bais.n1066 4.5
R17267 p_bais.n1080 p_bais.n1079 4.5
R17268 p_bais.n1070 p_bais.n1068 4.5
R17269 p_bais.n925 p_bais.n924 4.5
R17270 p_bais.n962 p_bais.n961 4.5
R17271 p_bais.n943 p_bais.n934 4.5
R17272 p_bais.n891 p_bais.n888 4.5
R17273 p_bais.n939 p_bais.n938 4.5
R17274 p_bais.n818 p_bais.n817 4.5
R17275 p_bais.n848 p_bais.n847 4.5
R17276 p_bais.n476 p_bais.n475 4.5
R17277 p_bais.n752 p_bais.n751 4.5
R17278 p_bais.n746 p_bais.n703 4.5
R17279 p_bais.n758 p_bais.n699 4.5
R17280 p_bais.n768 p_bais.n767 4.5
R17281 p_bais.n787 p_bais.n786 4.5
R17282 p_bais.n776 p_bais.n696 4.5
R17283 p_bais.n742 p_bais.n741 4.5
R17284 p_bais.n729 p_bais.n705 4.5
R17285 p_bais.n719 p_bais.n718 4.5
R17286 p_bais.n709 p_bais.n707 4.5
R17287 p_bais.n564 p_bais.n563 4.5
R17288 p_bais.n601 p_bais.n600 4.5
R17289 p_bais.n582 p_bais.n573 4.5
R17290 p_bais.n530 p_bais.n527 4.5
R17291 p_bais.n578 p_bais.n577 4.5
R17292 p_bais.n457 p_bais.n456 4.5
R17293 p_bais.n487 p_bais.n486 4.5
R17294 p_bais.n361 p_bais.n360 4.5
R17295 p_bais.n435 p_bais.n432 4.5
R17296 p_bais.n371 p_bais.n370 4.5
R17297 p_bais.n389 p_bais.n387 4.5
R17298 p_bais.n428 p_bais.n425 4.5
R17299 p_bais.n417 p_bais.n414 4.5
R17300 p_bais.n297 p_bais.n296 4.5
R17301 p_bais.n279 p_bais.n260 4.5
R17302 p_bais.n284 p_bais.n256 4.5
R17303 p_bais.n281 p_bais.n258 4.5
R17304 p_bais.n276 p_bais.n264 4.5
R17305 p_bais.n271 p_bais.n268 4.5
R17306 p_bais.n165 p_bais.n164 4.5
R17307 p_bais.n156 p_bais.n155 4.5
R17308 p_bais.n148 p_bais.n147 4.5
R17309 p_bais.n161 p_bais.n160 4.5
R17310 p_bais.n171 p_bais.n170 4.5
R17311 p_bais.n182 p_bais.n181 4.5
R17312 p_bais.n1060 p_bais.n1058 4.325
R17313 p_bais.n699 p_bais.n697 4.325
R17314 p_bais.n1153 p_bais.t1 4.289
R17315 p_bais.n792 p_bais.t0 4.289
R17316 p_bais.n403 p_bais.n402 3.992
R17317 p_bais.n329 p_bais.n327 3.992
R17318 p_bais.n1064 p_bais.n1061 3.95
R17319 p_bais.n703 p_bais.n700 3.95
R17320 p_bais.n817 p_bais.n816 3.948
R17321 p_bais.n456 p_bais.n455 3.948
R17322 p_bais.n341 p_bais.n340 3.882
R17323 p_bais.n212 p_bais.n210 3.882
R17324 p_bais.n1165 p_bais.n125 3.588
R17325 p_bais.n938 p_bais.n937 3.573
R17326 p_bais.n577 p_bais.n576 3.573
R17327 p_bais.n1163 p_bais.n1162 3.044
R17328 p_bais.n1163 p_bais.n801 3.044
R17329 p_bais.n951 p_bais.n932 3.033
R17330 p_bais.n826 p_bais.n825 3.033
R17331 p_bais.n590 p_bais.n571 3.033
R17332 p_bais.n465 p_bais.n464 3.033
R17333 p_bais.n186 p_bais.n139 2.797
R17334 p_bais.n357 p_bais.n355 2.787
R17335 p_bais.n293 p_bais.n291 2.787
R17336 p_bais.n301 p_bais.n253 2.742
R17337 p_bais.n358 p_bais.n354 2.695
R17338 p_bais.n294 p_bais.n290 2.695
R17339 p_bais.n179 p_bais.n177 2.695
R17340 p_bais.n387 p_bais.n386 2.656
R17341 p_bais.n137 p_bais.n136 2.535
R17342 p_bais.n251 p_bais.n250 2.415
R17343 p_bais.n1063 p_bais.n1062 2.258
R17344 p_bais.n936 p_bais.n935 2.258
R17345 p_bais.n702 p_bais.n701 2.258
R17346 p_bais.n575 p_bais.n574 2.258
R17347 p_bais.n119 p_bais.n118 2.25
R17348 p_bais.n62 p_bais.n61 2.25
R17349 p_bais.n369 p_bais.n368 2.082
R17350 p_bais.n424 p_bais.n423 2.082
R17351 p_bais.n359 p_bais.n358 2.082
R17352 p_bais.n413 p_bais.n412 2.082
R17353 p_bais.n255 p_bais.n254 2.082
R17354 p_bais.n263 p_bais.n262 2.082
R17355 p_bais.n295 p_bais.n294 2.082
R17356 p_bais.n267 p_bais.n266 2.082
R17357 p_bais.n146 p_bais.n145 2.082
R17358 p_bais.n154 p_bais.n153 2.082
R17359 p_bais.n169 p_bais.n168 2.082
R17360 p_bais.n180 p_bais.n179 2.082
R17361 p_bais.n1111 p_bais.n1110 1.882
R17362 p_bais.n1112 p_bais.n1111 1.882
R17363 p_bais.n887 p_bais.n886 1.882
R17364 p_bais.n750 p_bais.n749 1.882
R17365 p_bais.n751 p_bais.n750 1.882
R17366 p_bais.n526 p_bais.n525 1.882
R17367 p_bais.n1154 p_bais.n1153 1.844
R17368 p_bais.n793 p_bais.n792 1.844
R17369 p_bais.n1164 p_bais.n440 1.637
R17370 p_bais.n938 p_bais.n936 1.505
R17371 p_bais.n888 p_bais.n887 1.505
R17372 p_bais.n577 p_bais.n575 1.505
R17373 p_bais.n527 p_bais.n526 1.505
R17374 p_bais.n436 p_bais.n435 1.5
R17375 p_bais.n372 p_bais.n371 1.5
R17376 p_bais.n390 p_bais.n389 1.5
R17377 p_bais.n429 p_bais.n428 1.5
R17378 p_bais.n362 p_bais.n361 1.5
R17379 p_bais.n418 p_bais.n417 1.5
R17380 p_bais.n405 p_bais.n404 1.5
R17381 p_bais.n345 p_bais.n344 1.5
R17382 p_bais.n331 p_bais.n330 1.5
R17383 p_bais.n216 p_bais.n215 1.5
R17384 p_bais.n359 p_bais.n353 1.449
R17385 p_bais.n295 p_bais.n289 1.449
R17386 p_bais.n146 p_bais.n142 1.449
R17387 p_bais.n20 p_bais.n11 1.364
R17388 p_bais.n340 p_bais.n338 1.328
R17389 p_bais.n413 p_bais.n411 1.328
R17390 p_bais.n253 p_bais.n251 1.328
R17391 p_bais.n267 p_bais.n265 1.328
R17392 p_bais.n210 p_bais.n208 1.328
R17393 p_bais.n180 p_bais.n176 1.328
R17394 p_bais p_bais.n27 1.217
R17395 p_bais.n387 p_bais.n376 1.207
R17396 p_bais.n425 p_bais.n424 1.207
R17397 p_bais.n402 p_bais.n400 1.207
R17398 p_bais.n258 p_bais.n257 1.207
R17399 p_bais.n264 p_bais.n263 1.207
R17400 p_bais.n327 p_bais.n325 1.207
R17401 p_bais.n160 p_bais.n159 1.207
R17402 p_bais.n170 p_bais.n169 1.207
R17403 p_bais.n139 p_bais.n137 1.207
R17404 p_bais.n914 p_bais.n913 1.137
R17405 p_bais.n992 p_bais.n991 1.137
R17406 p_bais.n999 p_bais.n998 1.137
R17407 p_bais.n1003 p_bais.n1002 1.137
R17408 p_bais.n1010 p_bais.n1009 1.137
R17409 p_bais.n1028 p_bais.n1027 1.137
R17410 p_bais.n1045 p_bais.n1044 1.137
R17411 p_bais.n1052 p_bais.n1051 1.137
R17412 p_bais.n1041 p_bais.n1040 1.137
R17413 p_bais.n1034 p_bais.n1033 1.137
R17414 p_bais.n1020 p_bais.n1019 1.137
R17415 p_bais.n984 p_bais.n983 1.137
R17416 p_bais.n975 p_bais.n974 1.137
R17417 p_bais.n966 p_bais.n965 1.137
R17418 p_bais.n903 p_bais.n902 1.137
R17419 p_bais.n910 p_bais.n909 1.137
R17420 p_bais.n895 p_bais.n894 1.137
R17421 p_bais.n880 p_bais.n879 1.137
R17422 p_bais.n864 p_bais.n863 1.137
R17423 p_bais.n871 p_bais.n870 1.137
R17424 p_bais.n1162 p_bais.n1161 1.137
R17425 p_bais.n553 p_bais.n552 1.137
R17426 p_bais.n631 p_bais.n630 1.137
R17427 p_bais.n638 p_bais.n637 1.137
R17428 p_bais.n642 p_bais.n641 1.137
R17429 p_bais.n649 p_bais.n648 1.137
R17430 p_bais.n667 p_bais.n666 1.137
R17431 p_bais.n684 p_bais.n683 1.137
R17432 p_bais.n691 p_bais.n690 1.137
R17433 p_bais.n680 p_bais.n679 1.137
R17434 p_bais.n673 p_bais.n672 1.137
R17435 p_bais.n659 p_bais.n658 1.137
R17436 p_bais.n623 p_bais.n622 1.137
R17437 p_bais.n614 p_bais.n613 1.137
R17438 p_bais.n605 p_bais.n604 1.137
R17439 p_bais.n542 p_bais.n541 1.137
R17440 p_bais.n549 p_bais.n548 1.137
R17441 p_bais.n534 p_bais.n533 1.137
R17442 p_bais.n519 p_bais.n518 1.137
R17443 p_bais.n503 p_bais.n502 1.137
R17444 p_bais.n510 p_bais.n509 1.137
R17445 p_bais.n801 p_bais.n800 1.137
R17446 p_bais.n26 p_bais.n22 1.135
R17447 p_bais.n1057 p_bais.n1056 1.129
R17448 p_bais.n1064 p_bais.n1063 1.129
R17449 p_bais.n1102 p_bais.n1101 1.129
R17450 p_bais.n696 p_bais.n695 1.129
R17451 p_bais.n703 p_bais.n702 1.129
R17452 p_bais.n741 p_bais.n740 1.129
R17453 p_bais.n892 p_bais.n891 1.125
R17454 p_bais.n531 p_bais.n530 1.125
R17455 p_bais.n370 p_bais.n369 1.086
R17456 p_bais.n432 p_bais.n431 1.086
R17457 p_bais.n256 p_bais.n255 1.086
R17458 p_bais.n260 p_bais.n259 1.086
R17459 p_bais.n155 p_bais.n154 1.086
R17460 p_bais.n164 p_bais.n163 1.086
R17461 p_bais.n965 p_bais.n962 1.042
R17462 p_bais.n604 p_bais.n601 1.042
R17463 p_bais.n856 p_bais.n855 0.869
R17464 p_bais.n495 p_bais.n494 0.869
R17465 p_bais.n1147 p_bais.n1146 0.752
R17466 p_bais.n961 p_bais.n960 0.752
R17467 p_bais.n934 p_bais.n933 0.752
R17468 p_bais.n817 p_bais.n815 0.752
R17469 p_bais.n836 p_bais.n835 0.752
R17470 p_bais.n847 p_bais.n846 0.752
R17471 p_bais.n786 p_bais.n785 0.752
R17472 p_bais.n600 p_bais.n599 0.752
R17473 p_bais.n573 p_bais.n572 0.752
R17474 p_bais.n456 p_bais.n454 0.752
R17475 p_bais.n475 p_bais.n474 0.752
R17476 p_bais.n486 p_bais.n485 0.752
R17477 p_bais.n855 p_bais.n854 0.728
R17478 p_bais.n494 p_bais.n493 0.728
R17479 p_bais.n1161 p_bais.n1155 0.725
R17480 p_bais.n800 p_bais.n794 0.725
R17481 p_bais.n414 p_bais.n413 0.724
R17482 p_bais.n268 p_bais.n267 0.724
R17483 p_bais.n181 p_bais.n180 0.724
R17484 p_bais.n187 p_bais.n186 0.722
R17485 p_bais.n302 p_bais.n301 0.722
R17486 p_bais.n31 p_bais.n30 0.695
R17487 p_bais.n89 p_bais.n88 0.693
R17488 p_bais p_bais.n1165 0.618
R17489 p_bais.n360 p_bais.n359 0.603
R17490 p_bais.n296 p_bais.n295 0.603
R17491 p_bais.n147 p_bais.n146 0.603
R17492 p_bais.n43 p_bais.n42 0.559
R17493 p_bais.n122 p_bais.n121 0.559
R17494 p_bais.n73 p_bais.n72 0.559
R17495 p_bais.n91 p_bais.n85 0.559
R17496 p_bais.n423 p_bais.n422 0.557
R17497 p_bais.n262 p_bais.n261 0.557
R17498 p_bais.n1164 p_bais.n1163 0.478
R17499 p_bais.n1128 p_bais.n1127 0.376
R17500 p_bais.n1060 p_bais.n1059 0.376
R17501 p_bais.n1066 p_bais.n1065 0.376
R17502 p_bais.n1079 p_bais.n1078 0.376
R17503 p_bais.n1068 p_bais.n1067 0.376
R17504 p_bais.n924 p_bais.n923 0.376
R17505 p_bais.n767 p_bais.n766 0.376
R17506 p_bais.n699 p_bais.n698 0.376
R17507 p_bais.n705 p_bais.n704 0.376
R17508 p_bais.n718 p_bais.n717 0.376
R17509 p_bais.n707 p_bais.n706 0.376
R17510 p_bais.n563 p_bais.n562 0.376
R17511 p_bais.n1165 p_bais.n1164 0.241
R17512 p_bais.n1 p_bais.n0 0.197
R17513 p_bais.n2 p_bais.n1 0.197
R17514 p_bais.n3 p_bais.n2 0.197
R17515 p_bais.n16 p_bais.n15 0.197
R17516 p_bais.n15 p_bais.n14 0.197
R17517 p_bais.n14 p_bais.n13 0.197
R17518 p_bais.n13 p_bais.n12 0.197
R17519 p_bais.n4 p_bais.n3 0.196
R17520 p_bais.n927 p_bais.n926 0.189
R17521 p_bais.n566 p_bais.n565 0.189
R17522 p_bais.n1072 p_bais.n1071 0.188
R17523 p_bais.n711 p_bais.n710 0.188
R17524 p_bais.n17 p_bais.n16 0.188
R17525 p_bais.n5 p_bais.n4 0.184
R17526 p_bais.n948 p_bais.n947 0.166
R17527 p_bais.n587 p_bais.n586 0.166
R17528 p_bais.n1096 p_bais.n1095 0.166
R17529 p_bais.n735 p_bais.n734 0.166
R17530 p_bais.n825 p_bais.n824 0.133
R17531 p_bais.n464 p_bais.n463 0.133
R17532 p_bais.n1127 p_bais.n1126 0.132
R17533 p_bais.n766 p_bais.n765 0.132
R17534 p_bais.n835 p_bais.n834 0.121
R17535 p_bais.n474 p_bais.n473 0.121
R17536 p_bais.n1056 p_bais.n1055 0.121
R17537 p_bais.n695 p_bais.n694 0.121
R17538 p_bais.n11 p_bais.n10 0.112
R17539 p_bais.n9 p_bais.n8 0.056
R17540 p_bais.n10 p_bais.n9 0.056
R17541 p_bais.n1033 p_bais.n1032 0.049
R17542 p_bais.n1028 p_bais.n1020 0.049
R17543 p_bais.n984 p_bais.n975 0.049
R17544 p_bais.n895 p_bais.n880 0.049
R17545 p_bais.n672 p_bais.n671 0.049
R17546 p_bais.n667 p_bais.n659 0.049
R17547 p_bais.n623 p_bais.n614 0.049
R17548 p_bais.n534 p_bais.n519 0.049
R17549 p_bais.n300 p_bais.n299 0.048
R17550 p_bais.n287 p_bais.n286 0.048
R17551 p_bais.n274 p_bais.n273 0.048
R17552 p_bais.n151 p_bais.n150 0.048
R17553 p_bais.n174 p_bais.n173 0.048
R17554 p_bais.n185 p_bais.n184 0.048
R17555 p_bais.n1152 p_bais.n1151 0.047
R17556 p_bais.n1133 p_bais.n1131 0.047
R17557 p_bais.n1131 p_bais.n1130 0.047
R17558 p_bais.n1123 p_bais.n1121 0.047
R17559 p_bais.n1075 p_bais.n1074 0.047
R17560 p_bais.n930 p_bais.n929 0.047
R17561 p_bais.n822 p_bais.n820 0.047
R17562 p_bais.n827 p_bais.n826 0.047
R17563 p_bais.n830 p_bais.n828 0.047
R17564 p_bais.n852 p_bais.n851 0.047
R17565 p_bais.n990 p_bais.n989 0.047
R17566 p_bais.n791 p_bais.n790 0.047
R17567 p_bais.n772 p_bais.n770 0.047
R17568 p_bais.n770 p_bais.n769 0.047
R17569 p_bais.n762 p_bais.n760 0.047
R17570 p_bais.n714 p_bais.n713 0.047
R17571 p_bais.n569 p_bais.n568 0.047
R17572 p_bais.n461 p_bais.n459 0.047
R17573 p_bais.n466 p_bais.n465 0.047
R17574 p_bais.n469 p_bais.n467 0.047
R17575 p_bais.n491 p_bais.n490 0.047
R17576 p_bais.n629 p_bais.n628 0.047
R17577 p_bais.n81 p_bais.n80 0.046
R17578 p_bais.n96 p_bais.n95 0.046
R17579 p_bais.n68 p_bais.n67 0.046
R17580 p_bais.n37 p_bais.n36 0.046
R17581 p_bais.n1077 p_bais.n1076 0.045
R17582 p_bais.n931 p_bais.n930 0.045
R17583 p_bais.n716 p_bais.n715 0.045
R17584 p_bais.n570 p_bais.n569 0.045
R17585 p_bais.n280 p_bais.n279 0.044
R17586 p_bais.n165 p_bais.n162 0.044
R17587 p_bais.n1100 p_bais.n1099 0.043
R17588 p_bais.n891 p_bais.n885 0.043
R17589 p_bais.n983 p_bais.n982 0.043
R17590 p_bais.n893 p_bais.n892 0.043
R17591 p_bais.n878 p_bais.n877 0.043
R17592 p_bais.n739 p_bais.n738 0.043
R17593 p_bais.n530 p_bais.n524 0.043
R17594 p_bais.n622 p_bais.n621 0.043
R17595 p_bais.n532 p_bais.n531 0.043
R17596 p_bais.n517 p_bais.n516 0.043
R17597 p_bais.n107 p_bais.n106 0.043
R17598 p_bais.n114 p_bais.n113 0.043
R17599 p_bais.n47 p_bais.n46 0.043
R17600 p_bais.n57 p_bais.n56 0.043
R17601 p_bais.n87 p_bais.n86 0.043
R17602 p_bais.n78 p_bais.n77 0.043
R17603 p_bais.n93 p_bais.n92 0.043
R17604 p_bais.n65 p_bais.n64 0.043
R17605 p_bais.n34 p_bais.n33 0.043
R17606 p_bais.n29 p_bais.n28 0.043
R17607 p_bais.n1155 p_bais.n1152 0.043
R17608 p_bais.n794 p_bais.n791 0.043
R17609 p_bais.n389 p_bais.n388 0.042
R17610 p_bais.n281 p_bais.n280 0.042
R17611 p_bais.n162 p_bais.n161 0.042
R17612 p_bais.n1120 p_bais.n1119 0.041
R17613 p_bais.n1113 p_bais.n1109 0.041
R17614 p_bais.n921 p_bais.n920 0.041
R17615 p_bais.n945 p_bais.n944 0.041
R17616 p_bais.n842 p_bais.n841 0.041
R17617 p_bais.n1027 p_bais.n1026 0.041
R17618 p_bais.n901 p_bais.n900 0.041
R17619 p_bais.n759 p_bais.n758 0.041
R17620 p_bais.n752 p_bais.n748 0.041
R17621 p_bais.n560 p_bais.n559 0.041
R17622 p_bais.n584 p_bais.n583 0.041
R17623 p_bais.n481 p_bais.n480 0.041
R17624 p_bais.n666 p_bais.n665 0.041
R17625 p_bais.n540 p_bais.n539 0.041
R17626 p_bais.n854 p_bais.n852 0.041
R17627 p_bais.n493 p_bais.n491 0.041
R17628 p_bais.n1142 p_bais.n1141 0.039
R17629 p_bais.n1098 p_bais.n1097 0.039
R17630 p_bais.n949 p_bais.n946 0.039
R17631 p_bais.n819 p_bais.n818 0.039
R17632 p_bais.n879 p_bais.n874 0.039
R17633 p_bais.n781 p_bais.n780 0.039
R17634 p_bais.n737 p_bais.n736 0.039
R17635 p_bais.n588 p_bais.n585 0.039
R17636 p_bais.n458 p_bais.n457 0.039
R17637 p_bais.n518 p_bais.n513 0.039
R17638 p_bais.n1108 p_bais.n1107 0.037
R17639 p_bais.n747 p_bais.n746 0.037
R17640 p_bais.n72 p_bais.n63 0.036
R17641 p_bais.n85 p_bais.n76 0.036
R17642 p_bais.n371 p_bais.n367 0.036
R17643 p_bais.n285 p_bais.n284 0.036
R17644 p_bais.n156 p_bais.n152 0.036
R17645 p_bais.n121 p_bais.n120 0.035
R17646 p_bais.n42 p_bais.n41 0.035
R17647 p_bais.n809 p_bais.n808 0.035
R17648 p_bais.n448 p_bais.n447 0.035
R17649 p_bais.n120 p_bais.n119 0.035
R17650 p_bais.n63 p_bais.n62 0.035
R17651 p_bais.n1087 p_bais.n1086 0.034
R17652 p_bais.n919 p_bais.n918 0.034
R17653 p_bais.n1032 p_bais.n1031 0.034
R17654 p_bais.n1025 p_bais.n1024 0.034
R17655 p_bais.n981 p_bais.n980 0.034
R17656 p_bais.n970 p_bais.n969 0.034
R17657 p_bais.n892 p_bais.n883 0.034
R17658 p_bais.n877 p_bais.n876 0.034
R17659 p_bais.n726 p_bais.n725 0.034
R17660 p_bais.n558 p_bais.n557 0.034
R17661 p_bais.n671 p_bais.n670 0.034
R17662 p_bais.n664 p_bais.n663 0.034
R17663 p_bais.n620 p_bais.n619 0.034
R17664 p_bais.n609 p_bais.n608 0.034
R17665 p_bais.n531 p_bais.n522 0.034
R17666 p_bais.n516 p_bais.n515 0.034
R17667 p_bais.n428 p_bais.n427 0.034
R17668 p_bais.n276 p_bais.n275 0.034
R17669 p_bais.n172 p_bais.n171 0.034
R17670 p_bais.n82 p_bais.n81 0.034
R17671 p_bais.n97 p_bais.n96 0.034
R17672 p_bais.n69 p_bais.n68 0.034
R17673 p_bais.n38 p_bais.n37 0.034
R17674 p_bais.n230 p_bais.n229 0.033
R17675 p_bais.n335 p_bais.n334 0.033
R17676 p_bais.n438 p_bais.n335 0.033
R17677 p_bais.n1150 p_bais.n1149 0.032
R17678 p_bais.n957 p_bais.n954 0.032
R17679 p_bais.n850 p_bais.n849 0.032
R17680 p_bais.n988 p_bais.n987 0.032
R17681 p_bais.n789 p_bais.n788 0.032
R17682 p_bais.n596 p_bais.n593 0.032
R17683 p_bais.n489 p_bais.n488 0.032
R17684 p_bais.n627 p_bais.n626 0.032
R17685 p_bais.n438 p_bais.n230 0.032
R17686 p_bais.n110 p_bais.n109 0.032
R17687 p_bais.n117 p_bais.n116 0.032
R17688 p_bais.n50 p_bais.n49 0.032
R17689 p_bais.n60 p_bais.n59 0.032
R17690 p_bais.n72 p_bais.n71 0.031
R17691 p_bais.n85 p_bais.n84 0.031
R17692 p_bais.n1053 p_bais.n1052 0.031
R17693 p_bais.n1034 p_bais.n1030 0.031
R17694 p_bais.n1011 p_bais.n1010 0.031
R17695 p_bais.n992 p_bais.n986 0.031
R17696 p_bais.n967 p_bais.n966 0.031
R17697 p_bais.n903 p_bais.n897 0.031
R17698 p_bais.n872 p_bais.n871 0.031
R17699 p_bais.n857 p_bais.n856 0.031
R17700 p_bais.n692 p_bais.n691 0.031
R17701 p_bais.n673 p_bais.n669 0.031
R17702 p_bais.n650 p_bais.n649 0.031
R17703 p_bais.n631 p_bais.n625 0.031
R17704 p_bais.n606 p_bais.n605 0.031
R17705 p_bais.n542 p_bais.n536 0.031
R17706 p_bais.n511 p_bais.n510 0.031
R17707 p_bais.n496 p_bais.n495 0.031
R17708 p_bais.n42 p_bais.n40 0.031
R17709 p_bais.n121 p_bais.n99 0.031
R17710 p_bais.n1129 p_bais.n1125 0.03
R17711 p_bais.n1073 p_bais.n1070 0.03
R17712 p_bais.n928 p_bais.n925 0.03
R17713 p_bais.n823 p_bais.n822 0.03
R17714 p_bais.n840 p_bais.n839 0.03
R17715 p_bais.n972 p_bais.n971 0.03
R17716 p_bais.n768 p_bais.n764 0.03
R17717 p_bais.n712 p_bais.n709 0.03
R17718 p_bais.n567 p_bais.n564 0.03
R17719 p_bais.n462 p_bais.n461 0.03
R17720 p_bais.n479 p_bais.n478 0.03
R17721 p_bais.n611 p_bais.n610 0.03
R17722 p_bais.n301 p_bais.n300 0.028
R17723 p_bais.n1140 p_bais.n1139 0.028
R17724 p_bais.n1083 p_bais.n1081 0.028
R17725 p_bais.n962 p_bais.n959 0.028
R17726 p_bais.n952 p_bais.n951 0.028
R17727 p_bais.n1043 p_bais.n1042 0.028
R17728 p_bais.n1018 p_bais.n1017 0.028
R17729 p_bais.n1016 p_bais.n1015 0.028
R17730 p_bais.n977 p_bais.n976 0.028
R17731 p_bais.n779 p_bais.n778 0.028
R17732 p_bais.n722 p_bais.n720 0.028
R17733 p_bais.n601 p_bais.n598 0.028
R17734 p_bais.n591 p_bais.n590 0.028
R17735 p_bais.n682 p_bais.n681 0.028
R17736 p_bais.n657 p_bais.n656 0.028
R17737 p_bais.n655 p_bais.n654 0.028
R17738 p_bais.n616 p_bais.n615 0.028
R17739 p_bais.n361 p_bais.n350 0.028
R17740 p_bais.n298 p_bais.n297 0.028
R17741 p_bais.n148 p_bais.n141 0.028
R17742 p_bais.n83 p_bais.n82 0.028
R17743 p_bais.n98 p_bais.n97 0.028
R17744 p_bais.n70 p_bais.n69 0.028
R17745 p_bais.n39 p_bais.n38 0.028
R17746 p_bais.n855 p_bais.n812 0.027
R17747 p_bais.n494 p_bais.n451 0.027
R17748 p_bais.n1045 p_bais.n1041 0.027
R17749 p_bais.n1003 p_bais.n999 0.027
R17750 p_bais.n914 p_bais.n910 0.027
R17751 p_bais.n864 p_bais.n860 0.027
R17752 p_bais.n684 p_bais.n680 0.027
R17753 p_bais.n642 p_bais.n638 0.027
R17754 p_bais.n553 p_bais.n549 0.027
R17755 p_bais.n503 p_bais.n499 0.027
R17756 p_bais.n186 p_bais.n185 0.027
R17757 p_bais.n1090 p_bais.n1089 0.026
R17758 p_bais.n1158 p_bais.n1157 0.026
R17759 p_bais.n1001 p_bais.n1000 0.026
R17760 p_bais.n899 p_bais.n898 0.026
R17761 p_bais.n882 p_bais.n881 0.026
R17762 p_bais.n729 p_bais.n728 0.026
R17763 p_bais.n797 p_bais.n796 0.026
R17764 p_bais.n640 p_bais.n639 0.026
R17765 p_bais.n538 p_bais.n537 0.026
R17766 p_bais.n521 p_bais.n520 0.026
R17767 p_bais.n417 p_bais.n416 0.026
R17768 p_bais.n271 p_bais.n270 0.026
R17769 p_bais.n183 p_bais.n182 0.026
R17770 p_bais.n8 p_bais.n7 0.025
R17771 p_bais.n950 p_bais.n949 0.024
R17772 p_bais.n1051 p_bais.n1050 0.024
R17773 p_bais.n1040 p_bais.n1039 0.024
R17774 p_bais.n1009 p_bais.n1008 0.024
R17775 p_bais.n998 p_bais.n997 0.024
R17776 p_bais.n965 p_bais.n964 0.024
R17777 p_bais.n909 p_bais.n908 0.024
R17778 p_bais.n804 p_bais.n803 0.024
R17779 p_bais.n811 p_bais.n810 0.024
R17780 p_bais.n589 p_bais.n588 0.024
R17781 p_bais.n690 p_bais.n689 0.024
R17782 p_bais.n679 p_bais.n678 0.024
R17783 p_bais.n648 p_bais.n647 0.024
R17784 p_bais.n637 p_bais.n636 0.024
R17785 p_bais.n604 p_bais.n603 0.024
R17786 p_bais.n548 p_bais.n547 0.024
R17787 p_bais.n443 p_bais.n442 0.024
R17788 p_bais.n450 p_bais.n449 0.024
R17789 p_bais.n352 p_bais.n351 0.023
R17790 p_bais.n416 p_bais.n415 0.023
R17791 p_bais.n288 p_bais.n287 0.023
R17792 p_bais.n270 p_bais.n269 0.023
R17793 p_bais.n150 p_bais.n149 0.023
R17794 p_bais.n184 p_bais.n183 0.023
R17795 p_bais.n1094 p_bais.n1092 0.022
R17796 p_bais.n1089 p_bais.n1088 0.022
R17797 p_bais.n1160 p_bais.n1159 0.022
R17798 p_bais.n869 p_bais.n868 0.022
R17799 p_bais.n807 p_bais.n806 0.022
R17800 p_bais.n812 p_bais.n811 0.022
R17801 p_bais.n733 p_bais.n731 0.022
R17802 p_bais.n728 p_bais.n727 0.022
R17803 p_bais.n799 p_bais.n798 0.022
R17804 p_bais.n508 p_bais.n507 0.022
R17805 p_bais.n446 p_bais.n445 0.022
R17806 p_bais.n451 p_bais.n450 0.022
R17807 p_bais.n343 p_bais.n342 0.021
R17808 p_bais.n350 p_bais.n349 0.021
R17809 p_bais.n410 p_bais.n409 0.021
R17810 p_bais.n299 p_bais.n298 0.021
R17811 p_bais.n273 p_bais.n272 0.021
R17812 p_bais.n214 p_bais.n213 0.021
R17813 p_bais.n141 p_bais.n140 0.021
R17814 p_bais.n175 p_bais.n174 0.021
R17815 p_bais.n102 p_bais.n101 0.021
R17816 p_bais.n112 p_bais.n111 0.021
R17817 p_bais.n45 p_bais.n44 0.021
R17818 p_bais.n55 p_bais.n54 0.021
R17819 p_bais.n53 p_bais.n52 0.021
R17820 p_bais.n1105 p_bais.n1104 0.02
R17821 p_bais.n953 p_bais.n952 0.02
R17822 p_bais.n942 p_bais.n941 0.02
R17823 p_bais.n1159 p_bais.n1158 0.02
R17824 p_bais.n912 p_bais.n911 0.02
R17825 p_bais.n744 p_bais.n743 0.02
R17826 p_bais.n592 p_bais.n591 0.02
R17827 p_bais.n581 p_bais.n580 0.02
R17828 p_bais.n798 p_bais.n797 0.02
R17829 p_bais.n551 p_bais.n550 0.02
R17830 p_bais.n84 p_bais.n83 0.02
R17831 p_bais.n99 p_bais.n98 0.02
R17832 p_bais.n71 p_bais.n70 0.02
R17833 p_bais.n40 p_bais.n39 0.02
R17834 p_bais.n389 p_bais.n375 0.019
R17835 p_bais.n399 p_bais.n398 0.019
R17836 p_bais.n282 p_bais.n281 0.019
R17837 p_bais.n277 p_bais.n276 0.019
R17838 p_bais.n324 p_bais.n323 0.019
R17839 p_bais.n161 p_bais.n158 0.019
R17840 p_bais.n171 p_bais.n167 0.019
R17841 p_bais.n862 p_bais.n861 0.018
R17842 p_bais.n501 p_bais.n500 0.018
R17843 p_bais.n303 p_bais.n302 0.018
R17844 p_bais.n1117 p_bais.n1116 0.017
R17845 p_bais.n837 p_bais.n833 0.017
R17846 p_bais.n863 p_bais.n862 0.017
R17847 p_bais.n756 p_bais.n755 0.017
R17848 p_bais.n476 p_bais.n472 0.017
R17849 p_bais.n502 p_bais.n501 0.017
R17850 p_bais.n435 p_bais.n434 0.017
R17851 p_bais.n284 p_bais.n283 0.017
R17852 p_bais.n279 p_bais.n278 0.017
R17853 p_bais.n157 p_bais.n156 0.017
R17854 p_bais.n166 p_bais.n165 0.017
R17855 p_bais.n103 p_bais.n102 0.017
R17856 p_bais.n104 p_bais.n103 0.017
R17857 p_bais.n118 p_bais.n110 0.017
R17858 p_bais.n118 p_bais.n117 0.017
R17859 p_bais.n61 p_bais.n50 0.017
R17860 p_bais.n61 p_bais.n60 0.017
R17861 p_bais.n54 p_bais.n53 0.017
R17862 p_bais.n1054 p_bais.n1053 0.016
R17863 p_bais.n1030 p_bais.n1029 0.016
R17864 p_bais.n1012 p_bais.n1011 0.016
R17865 p_bais.n986 p_bais.n985 0.016
R17866 p_bais.n968 p_bais.n967 0.016
R17867 p_bais.n897 p_bais.n896 0.016
R17868 p_bais.n873 p_bais.n872 0.016
R17869 p_bais.n693 p_bais.n692 0.016
R17870 p_bais.n669 p_bais.n668 0.016
R17871 p_bais.n651 p_bais.n650 0.016
R17872 p_bais.n625 p_bais.n624 0.016
R17873 p_bais.n607 p_bais.n606 0.016
R17874 p_bais.n536 p_bais.n535 0.016
R17875 p_bais.n512 p_bais.n511 0.016
R17876 p_bais.n188 p_bais.n187 0.016
R17877 p_bais.n212 p_bais.n211 0.015
R17878 p_bais.n1145 p_bais.n1144 0.015
R17879 p_bais.n1139 p_bais.n1138 0.015
R17880 p_bais.n1137 p_bais.n1136 0.015
R17881 p_bais.n954 p_bais.n953 0.015
R17882 p_bais.n839 p_bais.n838 0.015
R17883 p_bais.n845 p_bais.n844 0.015
R17884 p_bais.n1050 p_bais.n1049 0.015
R17885 p_bais.n1040 p_bais.n1037 0.015
R17886 p_bais.n1039 p_bais.n1038 0.015
R17887 p_bais.n1017 p_bais.n1016 0.015
R17888 p_bais.n1008 p_bais.n1007 0.015
R17889 p_bais.n997 p_bais.n996 0.015
R17890 p_bais.n964 p_bais.n963 0.015
R17891 p_bais.n913 p_bais.n912 0.015
R17892 p_bais.n908 p_bais.n907 0.015
R17893 p_bais.n868 p_bais.n867 0.015
R17894 p_bais.n805 p_bais.n804 0.015
R17895 p_bais.n784 p_bais.n783 0.015
R17896 p_bais.n778 p_bais.n777 0.015
R17897 p_bais.n776 p_bais.n775 0.015
R17898 p_bais.n593 p_bais.n592 0.015
R17899 p_bais.n478 p_bais.n477 0.015
R17900 p_bais.n484 p_bais.n483 0.015
R17901 p_bais.n689 p_bais.n688 0.015
R17902 p_bais.n679 p_bais.n676 0.015
R17903 p_bais.n678 p_bais.n677 0.015
R17904 p_bais.n656 p_bais.n655 0.015
R17905 p_bais.n647 p_bais.n646 0.015
R17906 p_bais.n636 p_bais.n635 0.015
R17907 p_bais.n603 p_bais.n602 0.015
R17908 p_bais.n552 p_bais.n551 0.015
R17909 p_bais.n547 p_bais.n546 0.015
R17910 p_bais.n507 p_bais.n506 0.015
R17911 p_bais.n444 p_bais.n443 0.015
R17912 p_bais.n427 p_bais.n426 0.015
R17913 p_bais.n275 p_bais.n274 0.015
R17914 p_bais.n173 p_bais.n172 0.015
R17915 p_bais.n25 p_bais.n24 0.015
R17916 p_bais.n26 p_bais.n25 0.014
R17917 p_bais.n307 p_bais.n306 0.014
R17918 p_bais.n364 p_bais.n363 0.014
R17919 p_bais.n203 p_bais.n202 0.014
R17920 p_bais.n108 p_bais.n107 0.014
R17921 p_bais.n115 p_bais.n114 0.014
R17922 p_bais.n48 p_bais.n47 0.014
R17923 p_bais.n58 p_bais.n57 0.014
R17924 p_bais.n329 p_bais.n328 0.014
R17925 p_bais.n1148 p_bais.n1145 0.013
R17926 p_bais.n1088 p_bais.n1087 0.013
R17927 p_bais.n848 p_bais.n845 0.013
R17928 p_bais.n1051 p_bais.n1048 0.013
R17929 p_bais.n998 p_bais.n995 0.013
R17930 p_bais.n971 p_bais.n970 0.013
R17931 p_bais.n808 p_bais.n807 0.013
R17932 p_bais.n787 p_bais.n784 0.013
R17933 p_bais.n727 p_bais.n726 0.013
R17934 p_bais.n487 p_bais.n484 0.013
R17935 p_bais.n690 p_bais.n687 0.013
R17936 p_bais.n637 p_bais.n634 0.013
R17937 p_bais.n610 p_bais.n609 0.013
R17938 p_bais.n447 p_bais.n446 0.013
R17939 p_bais.n367 p_bais.n366 0.013
R17940 p_bais.n404 p_bais.n399 0.013
R17941 p_bais.n286 p_bais.n285 0.013
R17942 p_bais.n330 p_bais.n324 0.013
R17943 p_bais.n152 p_bais.n151 0.013
R17944 p_bais.n313 p_bais.n312 0.013
R17945 p_bais.n318 p_bais.n317 0.013
R17946 p_bais.n420 p_bais.n419 0.013
R17947 p_bais.n197 p_bais.n196 0.013
R17948 p_bais.n192 p_bais.n191 0.013
R17949 p_bais.n312 p_bais.n311 0.012
R17950 p_bais.n331 p_bais.n322 0.012
R17951 p_bais.n346 p_bais.n345 0.012
R17952 p_bais.n347 p_bais.n346 0.012
R17953 p_bais.n391 p_bais.n390 0.012
R17954 p_bais.n437 p_bais.n436 0.012
R17955 p_bais.n406 p_bais.n405 0.012
R17956 p_bais.n216 p_bais.n207 0.012
R17957 p_bais.n207 p_bais.n206 0.012
R17958 p_bais.n198 p_bais.n197 0.012
R17959 p_bais.n1136 p_bais.n1135 0.011
R17960 p_bais.n1106 p_bais.n1105 0.011
R17961 p_bais.n941 p_bais.n940 0.011
R17962 p_bais.n833 p_bais.n832 0.011
R17963 p_bais.n775 p_bais.n774 0.011
R17964 p_bais.n745 p_bais.n744 0.011
R17965 p_bais.n580 p_bais.n579 0.011
R17966 p_bais.n472 p_bais.n471 0.011
R17967 p_bais.n344 p_bais.n343 0.011
R17968 p_bais.n417 p_bais.n410 0.011
R17969 p_bais.n272 p_bais.n271 0.011
R17970 p_bais.n215 p_bais.n214 0.011
R17971 p_bais.n182 p_bais.n175 0.011
R17972 p_bais.n322 p_bais.n321 0.011
R17973 p_bais.n407 p_bais.n406 0.011
R17974 p_bais.n24 p_bais.n23 0.01
R17975 p_bais.n309 p_bais.n308 0.01
R17976 p_bais.n316 p_bais.n315 0.01
R17977 p_bais.n319 p_bais.n318 0.01
R17978 p_bais.n372 p_bais.n365 0.01
R17979 p_bais.n429 p_bais.n421 0.01
R17980 p_bais.n419 p_bais.n418 0.01
R17981 p_bais.n201 p_bais.n200 0.01
R17982 p_bais.n194 p_bais.n193 0.01
R17983 p_bais.n191 p_bais.n190 0.01
R17984 p_bais.n109 p_bais.n108 0.01
R17985 p_bais.n116 p_bais.n115 0.01
R17986 p_bais.n49 p_bais.n48 0.01
R17987 p_bais.n59 p_bais.n58 0.01
R17988 p_bais.n333 p_bais.n240 0.009
R17989 p_bais.n27 p_bais.n26 0.009
R17990 p_bais.n1144 p_bais.n1142 0.009
R17991 p_bais.n1116 p_bais.n1115 0.009
R17992 p_bais.n890 p_bais.n889 0.009
R17993 p_bais.n820 p_bais.n819 0.009
R17994 p_bais.n851 p_bais.n850 0.009
R17995 p_bais.n1161 p_bais.n1160 0.009
R17996 p_bais.n1019 p_bais.n1018 0.009
R17997 p_bais.n1002 p_bais.n1001 0.009
R17998 p_bais.n894 p_bais.n882 0.009
R17999 p_bais.n879 p_bais.n878 0.009
R18000 p_bais.n810 p_bais.n809 0.009
R18001 p_bais.n1052 p_bais.n1047 0.009
R18002 p_bais.n1046 p_bais.n1045 0.009
R18003 p_bais.n1041 p_bais.n1036 0.009
R18004 p_bais.n1035 p_bais.n1034 0.009
R18005 p_bais.n1010 p_bais.n1005 0.009
R18006 p_bais.n1004 p_bais.n1003 0.009
R18007 p_bais.n999 p_bais.n994 0.009
R18008 p_bais.n993 p_bais.n992 0.009
R18009 p_bais.n966 p_bais.n916 0.009
R18010 p_bais.n915 p_bais.n914 0.009
R18011 p_bais.n910 p_bais.n905 0.009
R18012 p_bais.n904 p_bais.n903 0.009
R18013 p_bais.n871 p_bais.n866 0.009
R18014 p_bais.n865 p_bais.n864 0.009
R18015 p_bais.n860 p_bais.n859 0.009
R18016 p_bais.n858 p_bais.n857 0.009
R18017 p_bais.n783 p_bais.n781 0.009
R18018 p_bais.n755 p_bais.n754 0.009
R18019 p_bais.n529 p_bais.n528 0.009
R18020 p_bais.n459 p_bais.n458 0.009
R18021 p_bais.n490 p_bais.n489 0.009
R18022 p_bais.n800 p_bais.n799 0.009
R18023 p_bais.n658 p_bais.n657 0.009
R18024 p_bais.n641 p_bais.n640 0.009
R18025 p_bais.n533 p_bais.n521 0.009
R18026 p_bais.n518 p_bais.n517 0.009
R18027 p_bais.n449 p_bais.n448 0.009
R18028 p_bais.n691 p_bais.n686 0.009
R18029 p_bais.n685 p_bais.n684 0.009
R18030 p_bais.n680 p_bais.n675 0.009
R18031 p_bais.n674 p_bais.n673 0.009
R18032 p_bais.n649 p_bais.n644 0.009
R18033 p_bais.n643 p_bais.n642 0.009
R18034 p_bais.n638 p_bais.n633 0.009
R18035 p_bais.n632 p_bais.n631 0.009
R18036 p_bais.n605 p_bais.n555 0.009
R18037 p_bais.n554 p_bais.n553 0.009
R18038 p_bais.n549 p_bais.n544 0.009
R18039 p_bais.n543 p_bais.n542 0.009
R18040 p_bais.n510 p_bais.n505 0.009
R18041 p_bais.n504 p_bais.n503 0.009
R18042 p_bais.n499 p_bais.n498 0.009
R18043 p_bais.n497 p_bais.n496 0.009
R18044 p_bais.n361 p_bais.n352 0.009
R18045 p_bais.n297 p_bais.n288 0.009
R18046 p_bais.n149 p_bais.n148 0.009
R18047 p_bais.n306 p_bais.n305 0.009
R18048 p_bais.n363 p_bais.n362 0.009
R18049 p_bais.n204 p_bais.n203 0.009
R18050 p_bais.n228 p_bais.n227 0.009
R18051 p_bais.n305 p_bais.n304 0.008
R18052 p_bais.n315 p_bais.n314 0.008
R18053 p_bais.n320 p_bais.n319 0.008
R18054 p_bais.n362 p_bais.n348 0.008
R18055 p_bais.n430 p_bais.n429 0.008
R18056 p_bais.n418 p_bais.n408 0.008
R18057 p_bais.n205 p_bais.n204 0.008
R18058 p_bais.n195 p_bais.n194 0.008
R18059 p_bais.n190 p_bais.n189 0.008
R18060 p_bais.n36 p_bais.n35 0.008
R18061 p_bais.n67 p_bais.n66 0.008
R18062 p_bais.n95 p_bais.n94 0.008
R18063 p_bais.n80 p_bais.n79 0.008
R18064 p_bais.n1151 p_bais.n1150 0.007
R18065 p_bais.n1141 p_bais.n1140 0.007
R18066 p_bais.n1121 p_bais.n1120 0.007
R18067 p_bais.n1115 p_bais.n1114 0.007
R18068 p_bais.n1092 p_bais.n1091 0.007
R18069 p_bais.n920 p_bais.n919 0.007
R18070 p_bais.n929 p_bais.n928 0.007
R18071 p_bais.n951 p_bais.n950 0.007
R18072 p_bais.n946 p_bais.n945 0.007
R18073 p_bais.n944 p_bais.n943 0.007
R18074 p_bais.n940 p_bais.n939 0.007
R18075 p_bais.n891 p_bais.n890 0.007
R18076 p_bais.n844 p_bais.n842 0.007
R18077 p_bais.n1157 p_bais.n1156 0.007
R18078 p_bais.n1044 p_bais.n1043 0.007
R18079 p_bais.n1027 p_bais.n1022 0.007
R18080 p_bais.n1026 p_bais.n1025 0.007
R18081 p_bais.n978 p_bais.n977 0.007
R18082 p_bais.n980 p_bais.n979 0.007
R18083 p_bais.n973 p_bais.n972 0.007
R18084 p_bais.n909 p_bais.n906 0.007
R18085 p_bais.n902 p_bais.n901 0.007
R18086 p_bais.n900 p_bais.n899 0.007
R18087 p_bais.n790 p_bais.n789 0.007
R18088 p_bais.n780 p_bais.n779 0.007
R18089 p_bais.n760 p_bais.n759 0.007
R18090 p_bais.n754 p_bais.n753 0.007
R18091 p_bais.n731 p_bais.n730 0.007
R18092 p_bais.n559 p_bais.n558 0.007
R18093 p_bais.n568 p_bais.n567 0.007
R18094 p_bais.n590 p_bais.n589 0.007
R18095 p_bais.n585 p_bais.n584 0.007
R18096 p_bais.n583 p_bais.n582 0.007
R18097 p_bais.n579 p_bais.n578 0.007
R18098 p_bais.n530 p_bais.n529 0.007
R18099 p_bais.n483 p_bais.n481 0.007
R18100 p_bais.n796 p_bais.n795 0.007
R18101 p_bais.n683 p_bais.n682 0.007
R18102 p_bais.n666 p_bais.n661 0.007
R18103 p_bais.n665 p_bais.n664 0.007
R18104 p_bais.n617 p_bais.n616 0.007
R18105 p_bais.n619 p_bais.n618 0.007
R18106 p_bais.n612 p_bais.n611 0.007
R18107 p_bais.n548 p_bais.n545 0.007
R18108 p_bais.n541 p_bais.n540 0.007
R18109 p_bais.n539 p_bais.n538 0.007
R18110 p_bais.n375 p_bais.n374 0.007
R18111 p_bais.n434 p_bais.n433 0.007
R18112 p_bais.n227 p_bais.n226 0.007
R18113 p_bais.n226 p_bais.n225 0.007
R18114 p_bais.n225 p_bais.n224 0.007
R18115 p_bais.n224 p_bais.n223 0.007
R18116 p_bais.n223 p_bais.n222 0.007
R18117 p_bais.n222 p_bais.n221 0.007
R18118 p_bais.n221 p_bais.n220 0.007
R18119 p_bais.n220 p_bais.n219 0.007
R18120 p_bais.n219 p_bais.n218 0.007
R18121 p_bais.n232 p_bais.n231 0.007
R18122 p_bais.n233 p_bais.n232 0.007
R18123 p_bais.n234 p_bais.n233 0.007
R18124 p_bais.n235 p_bais.n234 0.007
R18125 p_bais.n236 p_bais.n235 0.007
R18126 p_bais.n237 p_bais.n236 0.007
R18127 p_bais.n238 p_bais.n237 0.007
R18128 p_bais.n239 p_bais.n238 0.007
R18129 p_bais.n240 p_bais.n239 0.007
R18130 p_bais.n283 p_bais.n282 0.007
R18131 p_bais.n278 p_bais.n277 0.007
R18132 p_bais.n158 p_bais.n157 0.007
R18133 p_bais.n167 p_bais.n166 0.007
R18134 p_bais.n310 p_bais.n309 0.007
R18135 p_bais.n373 p_bais.n372 0.007
R18136 p_bais.n200 p_bais.n199 0.007
R18137 p_bais.n215 p_bais.n212 0.007
R18138 p_bais.n344 p_bais.n341 0.007
R18139 p_bais.n404 p_bais.n403 0.006
R18140 p_bais.n330 p_bais.n329 0.006
R18141 p_bais.n304 p_bais.n303 0.006
R18142 p_bais.n321 p_bais.n320 0.006
R18143 p_bais.n345 p_bais.n337 0.006
R18144 p_bais.n348 p_bais.n347 0.006
R18145 p_bais.n408 p_bais.n407 0.006
R18146 p_bais.n217 p_bais.n216 0.006
R18147 p_bais.n206 p_bais.n205 0.006
R18148 p_bais.n189 p_bais.n188 0.006
R18149 p_bais.n333 p_bais.n332 0.005
R18150 p_bais.n1138 p_bais.n1137 0.005
R18151 p_bais.n1135 p_bais.n1133 0.005
R18152 p_bais.n1118 p_bais.n1117 0.005
R18153 p_bais.n1109 p_bais.n1108 0.005
R18154 p_bais.n1107 p_bais.n1106 0.005
R18155 p_bais.n1104 p_bais.n1103 0.005
R18156 p_bais.n1103 p_bais.n1100 0.005
R18157 p_bais.n1099 p_bais.n1098 0.005
R18158 p_bais.n1074 p_bais.n1073 0.005
R18159 p_bais.n918 p_bais.n917 0.005
R18160 p_bais.n885 p_bais.n884 0.005
R18161 p_bais.n814 p_bais.n813 0.005
R18162 p_bais.n841 p_bais.n840 0.005
R18163 p_bais.n1019 p_bais.n1013 0.005
R18164 p_bais.n1015 p_bais.n1014 0.005
R18165 p_bais.n1009 p_bais.n1006 0.005
R18166 p_bais.n982 p_bais.n981 0.005
R18167 p_bais.n894 p_bais.n893 0.005
R18168 p_bais.n803 p_bais.n802 0.005
R18169 p_bais.n1047 p_bais.n1046 0.005
R18170 p_bais.n1036 p_bais.n1035 0.005
R18171 p_bais.n1005 p_bais.n1004 0.005
R18172 p_bais.n994 p_bais.n993 0.005
R18173 p_bais.n916 p_bais.n915 0.005
R18174 p_bais.n905 p_bais.n904 0.005
R18175 p_bais.n866 p_bais.n865 0.005
R18176 p_bais.n859 p_bais.n858 0.005
R18177 p_bais.n777 p_bais.n776 0.005
R18178 p_bais.n774 p_bais.n772 0.005
R18179 p_bais.n757 p_bais.n756 0.005
R18180 p_bais.n748 p_bais.n747 0.005
R18181 p_bais.n746 p_bais.n745 0.005
R18182 p_bais.n743 p_bais.n742 0.005
R18183 p_bais.n742 p_bais.n739 0.005
R18184 p_bais.n738 p_bais.n737 0.005
R18185 p_bais.n713 p_bais.n712 0.005
R18186 p_bais.n557 p_bais.n556 0.005
R18187 p_bais.n524 p_bais.n523 0.005
R18188 p_bais.n453 p_bais.n452 0.005
R18189 p_bais.n480 p_bais.n479 0.005
R18190 p_bais.n658 p_bais.n652 0.005
R18191 p_bais.n654 p_bais.n653 0.005
R18192 p_bais.n648 p_bais.n645 0.005
R18193 p_bais.n621 p_bais.n620 0.005
R18194 p_bais.n533 p_bais.n532 0.005
R18195 p_bais.n442 p_bais.n441 0.005
R18196 p_bais.n686 p_bais.n685 0.005
R18197 p_bais.n675 p_bais.n674 0.005
R18198 p_bais.n644 p_bais.n643 0.005
R18199 p_bais.n633 p_bais.n632 0.005
R18200 p_bais.n555 p_bais.n554 0.005
R18201 p_bais.n544 p_bais.n543 0.005
R18202 p_bais.n505 p_bais.n504 0.005
R18203 p_bais.n498 p_bais.n497 0.005
R18204 p_bais.n311 p_bais.n310 0.005
R18205 p_bais.n314 p_bais.n313 0.005
R18206 p_bais.n332 p_bais.n331 0.005
R18207 p_bais.n390 p_bais.n373 0.005
R18208 p_bais.n436 p_bais.n430 0.005
R18209 p_bais.n405 p_bais.n397 0.005
R18210 p_bais.n199 p_bais.n198 0.005
R18211 p_bais.n196 p_bais.n195 0.005
R18212 p_bais.n88 p_bais.n87 0.005
R18213 p_bais.n79 p_bais.n78 0.005
R18214 p_bais.n94 p_bais.n93 0.005
R18215 p_bais.n66 p_bais.n65 0.005
R18216 p_bais.n35 p_bais.n34 0.005
R18217 p_bais.n30 p_bais.n29 0.005
R18218 p_bais.n18 p_bais.n17 0.005
R18219 p_bais.n19 p_bais.n18 0.005
R18220 p_bais.n22 p_bais.n6 0.005
R18221 p_bais.n6 p_bais.n5 0.005
R18222 p_bais.n228 p_bais.n217 0.005
R18223 p_bais.n397 p_bais.n396 0.004
R18224 p_bais.n378 p_bais.n377 0.004
R18225 p_bais.n386 p_bais.n378 0.004
R18226 p_bais.n382 p_bais.n381 0.004
R18227 p_bais.n386 p_bais.n382 0.004
R18228 p_bais.n380 p_bais.n379 0.004
R18229 p_bais.n386 p_bais.n380 0.004
R18230 p_bais.n384 p_bais.n383 0.004
R18231 p_bais.n250 p_bais.n249 0.004
R18232 p_bais.n249 p_bais.n248 0.004
R18233 p_bais.n244 p_bais.n243 0.004
R18234 p_bais.n248 p_bais.n244 0.004
R18235 p_bais.n242 p_bais.n241 0.004
R18236 p_bais.n248 p_bais.n242 0.004
R18237 p_bais.n246 p_bais.n245 0.004
R18238 p_bais.n136 p_bais.n135 0.004
R18239 p_bais.n135 p_bais.n134 0.004
R18240 p_bais.n133 p_bais.n132 0.004
R18241 p_bais.n134 p_bais.n133 0.004
R18242 p_bais.n130 p_bais.n129 0.004
R18243 p_bais.n127 p_bais.n126 0.004
R18244 p_bais.n308 p_bais.n307 0.004
R18245 p_bais.n317 p_bais.n316 0.004
R18246 p_bais.n365 p_bais.n364 0.004
R18247 p_bais.n421 p_bais.n420 0.004
R18248 p_bais.n202 p_bais.n201 0.004
R18249 p_bais.n193 p_bais.n192 0.004
R18250 p_bais.n105 p_bais.n104 0.004
R18251 p_bais.n337 p_bais.n336 0.004
R18252 p_bais.n334 p_bais.n333 0.003
R18253 p_bais.n1149 p_bais.n1148 0.003
R18254 p_bais.n962 p_bais.n931 0.003
R18255 p_bais.n959 p_bais.n957 0.003
R18256 p_bais.n943 p_bais.n942 0.003
R18257 p_bais.n818 p_bais.n814 0.003
R18258 p_bais.n832 p_bais.n830 0.003
R18259 p_bais.n838 p_bais.n837 0.003
R18260 p_bais.n849 p_bais.n848 0.003
R18261 p_bais.n1162 p_bais.n1054 0.003
R18262 p_bais.n1029 p_bais.n1028 0.003
R18263 p_bais.n1020 p_bais.n1012 0.003
R18264 p_bais.n985 p_bais.n984 0.003
R18265 p_bais.n975 p_bais.n968 0.003
R18266 p_bais.n896 p_bais.n895 0.003
R18267 p_bais.n880 p_bais.n873 0.003
R18268 p_bais.n788 p_bais.n787 0.003
R18269 p_bais.n601 p_bais.n570 0.003
R18270 p_bais.n598 p_bais.n596 0.003
R18271 p_bais.n582 p_bais.n581 0.003
R18272 p_bais.n457 p_bais.n453 0.003
R18273 p_bais.n471 p_bais.n469 0.003
R18274 p_bais.n477 p_bais.n476 0.003
R18275 p_bais.n488 p_bais.n487 0.003
R18276 p_bais.n801 p_bais.n693 0.003
R18277 p_bais.n668 p_bais.n667 0.003
R18278 p_bais.n659 p_bais.n651 0.003
R18279 p_bais.n624 p_bais.n623 0.003
R18280 p_bais.n614 p_bais.n607 0.003
R18281 p_bais.n535 p_bais.n534 0.003
R18282 p_bais.n519 p_bais.n512 0.003
R18283 p_bais.n229 p_bais.n228 0.003
R18284 p_bais.n385 p_bais.n384 0.002
R18285 p_bais.n386 p_bais.n385 0.002
R18286 p_bais.n247 p_bais.n246 0.002
R18287 p_bais.n248 p_bais.n247 0.002
R18288 p_bais.n131 p_bais.n130 0.002
R18289 p_bais.n128 p_bais.n127 0.002
R18290 p_bais.n134 p_bais.n131 0.002
R18291 p_bais.n134 p_bais.n128 0.002
R18292 p_bais.n439 p_bais.n438 0.002
R18293 p_bais.n101 p_bais.n100 0.002
R18294 p_bais.n106 p_bais.n105 0.002
R18295 p_bais.n113 p_bais.n112 0.002
R18296 p_bais.n46 p_bais.n45 0.002
R18297 p_bais.n56 p_bais.n55 0.002
R18298 p_bais.n52 p_bais.n51 0.002
R18299 p_bais.n91 p_bais.n90 0.002
R18300 p_bais.n122 p_bais.n91 0.002
R18301 p_bais.n123 p_bais.n122 0.002
R18302 p_bais.n125 p_bais.n124 0.002
R18303 p_bais.n74 p_bais.n73 0.002
R18304 p_bais.n73 p_bais.n43 0.002
R18305 p_bais.n43 p_bais.n32 0.002
R18306 p_bais.n394 p_bais.n393 0.001
R18307 p_bais.n393 p_bais.n392 0.001
R18308 p_bais.n395 p_bais.n394 0.001
R18309 p_bais.n395 p_bais.n391 0.001
R18310 p_bais.n21 p_bais.n20 0.001
R18311 p_bais.n1130 p_bais.n1129 0.001
R18312 p_bais.n1125 p_bais.n1123 0.001
R18313 p_bais.n1119 p_bais.n1118 0.001
R18314 p_bais.n1114 p_bais.n1113 0.001
R18315 p_bais.n1097 p_bais.n1094 0.001
R18316 p_bais.n1091 p_bais.n1090 0.001
R18317 p_bais.n1086 p_bais.n1083 0.001
R18318 p_bais.n1081 p_bais.n1080 0.001
R18319 p_bais.n1080 p_bais.n1077 0.001
R18320 p_bais.n1076 p_bais.n1075 0.001
R18321 p_bais.n1070 p_bais.n1069 0.001
R18322 p_bais.n925 p_bais.n921 0.001
R18323 p_bais.n826 p_bais.n823 0.001
R18324 p_bais.n828 p_bais.n827 0.001
R18325 p_bais.n1022 p_bais.n1021 0.001
R18326 p_bais.n1024 p_bais.n1023 0.001
R18327 p_bais.n991 p_bais.n990 0.001
R18328 p_bais.n989 p_bais.n988 0.001
R18329 p_bais.n983 p_bais.n978 0.001
R18330 p_bais.n974 p_bais.n973 0.001
R18331 p_bais.n876 p_bais.n875 0.001
R18332 p_bais.n870 p_bais.n869 0.001
R18333 p_bais.n806 p_bais.n805 0.001
R18334 p_bais.n769 p_bais.n768 0.001
R18335 p_bais.n764 p_bais.n762 0.001
R18336 p_bais.n758 p_bais.n757 0.001
R18337 p_bais.n753 p_bais.n752 0.001
R18338 p_bais.n736 p_bais.n733 0.001
R18339 p_bais.n730 p_bais.n729 0.001
R18340 p_bais.n725 p_bais.n722 0.001
R18341 p_bais.n720 p_bais.n719 0.001
R18342 p_bais.n719 p_bais.n716 0.001
R18343 p_bais.n715 p_bais.n714 0.001
R18344 p_bais.n709 p_bais.n708 0.001
R18345 p_bais.n564 p_bais.n560 0.001
R18346 p_bais.n465 p_bais.n462 0.001
R18347 p_bais.n467 p_bais.n466 0.001
R18348 p_bais.n661 p_bais.n660 0.001
R18349 p_bais.n663 p_bais.n662 0.001
R18350 p_bais.n630 p_bais.n629 0.001
R18351 p_bais.n628 p_bais.n627 0.001
R18352 p_bais.n622 p_bais.n617 0.001
R18353 p_bais.n613 p_bais.n612 0.001
R18354 p_bais.n515 p_bais.n514 0.001
R18355 p_bais.n509 p_bais.n508 0.001
R18356 p_bais.n445 p_bais.n444 0.001
R18357 p_bais.n440 p_bais.n439 0.001
R18358 p_bais.n438 p_bais.n437 0.001
R18359 p_bais.n90 p_bais.n89 0.001
R18360 p_bais.n124 p_bais.n123 0.001
R18361 p_bais.n125 p_bais.n75 0.001
R18362 p_bais.n75 p_bais.n74 0.001
R18363 p_bais.n32 p_bais.n31 0.001
R18364 p_bais.n22 p_bais.n21 0.001
R18365 p_bais.n20 p_bais.n19 0.001
R18366 p_bais.n437 p_bais.n395 0.001
R18367 net1_ota.n465 net1_ota.t0 39.189
R18368 net1_ota.n504 net1_ota.t3 17.4
R18369 net1_ota.n63 net1_ota.n62 9.3
R18370 net1_ota.n159 net1_ota.n158 9.3
R18371 net1_ota.n295 net1_ota.n294 9.3
R18372 net1_ota.n391 net1_ota.n390 9.3
R18373 net1_ota.n180 net1_ota.n179 8.886
R18374 net1_ota.n416 net1_ota.n415 8.886
R18375 net1_ota.n505 net1_ota.n504 8.5
R18376 net1_ota.n469 net1_ota.n468 8.282
R18377 net1_ota.n179 net1_ota.t1 7.141
R18378 net1_ota.n415 net1_ota.t2 7.141
R18379 net1_ota.n9 net1_ota.n8 7.033
R18380 net1_ota.n241 net1_ota.n240 7.033
R18381 net1_ota.n218 net1_ota.n217 7.03
R18382 net1_ota.n450 net1_ota.n449 7.03
R18383 net1_ota.n465 net1_ota.n464 6.101
R18384 net1_ota.n470 net1_ota.n469 4.5
R18385 net1_ota.n500 net1_ota.n499 4.5
R18386 net1_ota.n507 net1_ota.n506 4.5
R18387 net1_ota.n476 net1_ota.n475 4.5
R18388 net1_ota.n46 net1_ota.n45 4.5
R18389 net1_ota.n162 net1_ota.n154 4.5
R18390 net1_ota.n187 net1_ota.n182 4.5
R18391 net1_ota.n141 net1_ota.n140 4.5
R18392 net1_ota.n115 net1_ota.n113 4.5
R18393 net1_ota.n126 net1_ota.n121 4.5
R18394 net1_ota.n105 net1_ota.n102 4.5
R18395 net1_ota.n84 net1_ota.n83 4.5
R18396 net1_ota.n95 net1_ota.n90 4.5
R18397 net1_ota.n69 net1_ota.n68 4.5
R18398 net1_ota.n35 net1_ota.n34 4.5
R18399 net1_ota.n206 net1_ota.n205 4.5
R18400 net1_ota.n278 net1_ota.n277 4.5
R18401 net1_ota.n394 net1_ota.n386 4.5
R18402 net1_ota.n373 net1_ota.n372 4.5
R18403 net1_ota.n347 net1_ota.n345 4.5
R18404 net1_ota.n358 net1_ota.n353 4.5
R18405 net1_ota.n337 net1_ota.n334 4.5
R18406 net1_ota.n316 net1_ota.n315 4.5
R18407 net1_ota.n327 net1_ota.n322 4.5
R18408 net1_ota.n301 net1_ota.n300 4.5
R18409 net1_ota.n260 net1_ota.n259 4.5
R18410 net1_ota.n419 net1_ota.n418 4.5
R18411 net1_ota.n438 net1_ota.n437 4.5
R18412 net1_ota.n506 net1_ota.n503 4.141
R18413 net1_ota.n182 net1_ota.n178 4.141
R18414 net1_ota.n121 net1_ota.n120 4.141
R18415 net1_ota.n83 net1_ota.n82 4.141
R18416 net1_ota.n34 net1_ota.n33 4.141
R18417 net1_ota.n418 net1_ota.n414 4.141
R18418 net1_ota.n353 net1_ota.n352 4.141
R18419 net1_ota.n315 net1_ota.n314 4.141
R18420 net1_ota.n259 net1_ota.n258 4.141
R18421 net1_ota.n475 net1_ota.n474 3.764
R18422 net1_ota.n469 net1_ota.n467 3.764
R18423 net1_ota.n140 net1_ota.n139 3.764
R18424 net1_ota.n68 net1_ota.n67 3.764
R18425 net1_ota.n372 net1_ota.n371 3.764
R18426 net1_ota.n300 net1_ota.n299 3.764
R18427 net1_ota.n499 net1_ota.n498 3.388
R18428 net1_ota.n205 net1_ota.n202 3.388
R18429 net1_ota.n154 net1_ota.n151 3.388
R18430 net1_ota.n90 net1_ota.n88 3.388
R18431 net1_ota.n45 net1_ota.n44 3.388
R18432 net1_ota.n437 net1_ota.n434 3.388
R18433 net1_ota.n386 net1_ota.n383 3.388
R18434 net1_ota.n322 net1_ota.n320 3.388
R18435 net1_ota.n277 net1_ota.n276 3.388
R18436 net1_ota.n205 net1_ota.n204 3.011
R18437 net1_ota.n154 net1_ota.n153 3.011
R18438 net1_ota.n158 net1_ota.n157 3.011
R18439 net1_ota.n113 net1_ota.n111 3.011
R18440 net1_ota.n90 net1_ota.n89 3.011
R18441 net1_ota.n45 net1_ota.n43 3.011
R18442 net1_ota.n437 net1_ota.n436 3.011
R18443 net1_ota.n386 net1_ota.n385 3.011
R18444 net1_ota.n390 net1_ota.n389 3.011
R18445 net1_ota.n345 net1_ota.n343 3.011
R18446 net1_ota.n322 net1_ota.n321 3.011
R18447 net1_ota.n277 net1_ota.n275 3.011
R18448 net1_ota.n475 net1_ota.n473 2.635
R18449 net1_ota.n140 net1_ota.n137 2.635
R18450 net1_ota.n102 net1_ota.n101 2.635
R18451 net1_ota.n62 net1_ota.n61 2.635
R18452 net1_ota.n68 net1_ota.n66 2.635
R18453 net1_ota.n372 net1_ota.n369 2.635
R18454 net1_ota.n334 net1_ota.n333 2.635
R18455 net1_ota.n294 net1_ota.n293 2.635
R18456 net1_ota.n300 net1_ota.n298 2.635
R18457 net1_ota.n506 net1_ota.n505 2.258
R18458 net1_ota.n182 net1_ota.n181 2.258
R18459 net1_ota.n34 net1_ota.n32 2.258
R18460 net1_ota.n418 net1_ota.n417 2.258
R18461 net1_ota.n259 net1_ota.n257 2.258
R18462 net1_ota net1_ota.n510 2.24
R18463 net1_ota net1_ota.n465 1.603
R18464 net1_ota.n53 net1_ota.n9 1.508
R18465 net1_ota.n285 net1_ota.n241 1.508
R18466 net1_ota.n113 net1_ota.n112 1.505
R18467 net1_ota.n345 net1_ota.n344 1.505
R18468 net1_ota.n47 net1_ota.n46 1.5
R18469 net1_ota.n224 net1_ota.n223 1.5
R18470 net1_ota.n188 net1_ota.n187 1.5
R18471 net1_ota.n163 net1_ota.n162 1.5
R18472 net1_ota.n142 net1_ota.n141 1.5
R18473 net1_ota.n116 net1_ota.n115 1.5
R18474 net1_ota.n127 net1_ota.n126 1.5
R18475 net1_ota.n106 net1_ota.n105 1.5
R18476 net1_ota.n85 net1_ota.n84 1.5
R18477 net1_ota.n96 net1_ota.n95 1.5
R18478 net1_ota.n70 net1_ota.n69 1.5
R18479 net1_ota.n207 net1_ota.n206 1.5
R18480 net1_ota.n279 net1_ota.n278 1.5
R18481 net1_ota.n456 net1_ota.n455 1.5
R18482 net1_ota.n395 net1_ota.n394 1.5
R18483 net1_ota.n374 net1_ota.n373 1.5
R18484 net1_ota.n348 net1_ota.n347 1.5
R18485 net1_ota.n359 net1_ota.n358 1.5
R18486 net1_ota.n338 net1_ota.n337 1.5
R18487 net1_ota.n317 net1_ota.n316 1.5
R18488 net1_ota.n328 net1_ota.n327 1.5
R18489 net1_ota.n302 net1_ota.n301 1.5
R18490 net1_ota.n261 net1_ota.n260 1.5
R18491 net1_ota.n420 net1_ota.n419 1.5
R18492 net1_ota.n439 net1_ota.n438 1.5
R18493 net1_ota.n464 net1_ota.n463 1.426
R18494 net1_ota.n509 net1_ota.n508 1.384
R18495 net1_ota.n478 net1_ota.n477 1.384
R18496 net1_ota.n464 net1_ota.n231 1.169
R18497 net1_ota.n479 net1_ota.n478 1.146
R18498 net1_ota.n510 net1_ota.n509 1.137
R18499 net1_ota.n489 net1_ota.n488 1.137
R18500 net1_ota.n485 net1_ota.n484 1.137
R18501 net1_ota.n72 net1_ota.n71 1.137
R18502 net1_ota.n79 net1_ota.n78 1.137
R18503 net1_ota.n171 net1_ota.n170 1.137
R18504 net1_ota.n229 net1_ota.n228 1.137
R18505 net1_ota.n192 net1_ota.n191 1.137
R18506 net1_ota.n146 net1_ota.n145 1.137
R18507 net1_ota.n167 net1_ota.n166 1.137
R18508 net1_ota.n129 net1_ota.n128 1.137
R18509 net1_ota.n110 net1_ota.n109 1.137
R18510 net1_ota.n213 net1_ota.n212 1.137
R18511 net1_ota.n445 net1_ota.n444 1.137
R18512 net1_ota.n304 net1_ota.n303 1.137
R18513 net1_ota.n311 net1_ota.n310 1.137
R18514 net1_ota.n403 net1_ota.n402 1.137
R18515 net1_ota.n461 net1_ota.n460 1.137
R18516 net1_ota.n378 net1_ota.n377 1.137
R18517 net1_ota.n399 net1_ota.n398 1.137
R18518 net1_ota.n361 net1_ota.n360 1.137
R18519 net1_ota.n342 net1_ota.n341 1.137
R18520 net1_ota.n424 net1_ota.n423 1.137
R18521 net1_ota.n102 net1_ota.n100 1.129
R18522 net1_ota.n334 net1_ota.n332 1.129
R18523 net1_ota.n54 net1_ota.n53 0.72
R18524 net1_ota.n286 net1_ota.n285 0.72
R18525 net1_ota.n217 net1_ota.n216 0.155
R18526 net1_ota.n8 net1_ota.n7 0.155
R18527 net1_ota.n449 net1_ota.n448 0.155
R18528 net1_ota.n240 net1_ota.n239 0.155
R18529 net1_ota.n204 net1_ota.n203 0.144
R18530 net1_ota.n436 net1_ota.n435 0.144
R18531 net1_ota.n43 net1_ota.n42 0.144
R18532 net1_ota.n275 net1_ota.n274 0.144
R18533 net1_ota.n181 net1_ota.n180 0.133
R18534 net1_ota.n417 net1_ota.n416 0.133
R18535 net1_ota.n32 net1_ota.n31 0.132
R18536 net1_ota.n257 net1_ota.n256 0.132
R18537 net1_ota.n185 net1_ota.n184 0.056
R18538 net1_ota.n412 net1_ota.n411 0.056
R18539 net1_ota.n39 net1_ota.n38 0.047
R18540 net1_ota.n271 net1_ota.n270 0.047
R18541 net1_ota.n188 net1_ota.n174 0.045
R18542 net1_ota.n144 net1_ota.n143 0.045
R18543 net1_ota.n128 net1_ota.n127 0.045
R18544 net1_ota.n420 net1_ota.n406 0.045
R18545 net1_ota.n376 net1_ota.n375 0.045
R18546 net1_ota.n360 net1_ota.n359 0.045
R18547 net1_ota.n159 net1_ota.n156 0.043
R18548 net1_ota.n109 net1_ota.n85 0.043
R18549 net1_ota.n391 net1_ota.n388 0.043
R18550 net1_ota.n341 net1_ota.n317 0.043
R18551 net1_ota.n207 net1_ota.n195 0.041
R18552 net1_ota.n18 net1_ota.n17 0.041
R18553 net1_ota.n439 net1_ota.n427 0.041
R18554 net1_ota.n262 net1_ota.n261 0.041
R18555 net1_ota.n115 net1_ota.n114 0.039
R18556 net1_ota.n228 net1_ota.n227 0.039
R18557 net1_ota.n48 net1_ota.n47 0.039
R18558 net1_ota.n347 net1_ota.n346 0.039
R18559 net1_ota.n460 net1_ota.n459 0.039
R18560 net1_ota.n280 net1_ota.n279 0.039
R18561 net1_ota.n105 net1_ota.n99 0.037
R18562 net1_ota.n28 net1_ota.n27 0.037
R18563 net1_ota.n52 net1_ota.n51 0.037
R18564 net1_ota.n229 net1_ota.n213 0.037
R18565 net1_ota.n129 net1_ota.n110 0.037
R18566 net1_ota.n337 net1_ota.n331 0.037
R18567 net1_ota.n253 net1_ota.n252 0.037
R18568 net1_ota.n284 net1_ota.n283 0.037
R18569 net1_ota.n461 net1_ota.n445 0.037
R18570 net1_ota.n361 net1_ota.n342 0.037
R18571 net1_ota.n496 net1_ota.n495 0.035
R18572 net1_ota.n497 net1_ota.n496 0.035
R18573 net1_ota.n488 net1_ota.n486 0.035
R18574 net1_ota.n93 net1_ota.n92 0.034
R18575 net1_ota.n3 net1_ota.n2 0.034
R18576 net1_ota.n226 net1_ota.n225 0.034
R18577 net1_ota.n119 net1_ota.n118 0.034
R18578 net1_ota.n50 net1_ota.n49 0.034
R18579 net1_ota.n325 net1_ota.n324 0.034
R18580 net1_ota.n235 net1_ota.n234 0.034
R18581 net1_ota.n458 net1_ota.n457 0.034
R18582 net1_ota.n351 net1_ota.n350 0.034
R18583 net1_ota.n282 net1_ota.n281 0.034
R18584 net1_ota.n215 net1_ota.n214 0.032
R18585 net1_ota.n107 net1_ota.n106 0.032
R18586 net1_ota.n97 net1_ota.n96 0.032
R18587 net1_ota.n447 net1_ota.n446 0.032
R18588 net1_ota.n339 net1_ota.n338 0.032
R18589 net1_ota.n329 net1_ota.n328 0.032
R18590 net1_ota.n5 net1_ota.n4 0.03
R18591 net1_ota.n209 net1_ota.n208 0.03
R18592 net1_ota.n142 net1_ota.n132 0.03
R18593 net1_ota.n117 net1_ota.n116 0.03
R18594 net1_ota.n237 net1_ota.n236 0.03
R18595 net1_ota.n441 net1_ota.n440 0.03
R18596 net1_ota.n374 net1_ota.n364 0.03
R18597 net1_ota.n349 net1_ota.n348 0.03
R18598 net1_ota.n221 net1_ota.n220 0.028
R18599 net1_ota.n20 net1_ota.n19 0.028
R18600 net1_ota.n453 net1_ota.n452 0.028
R18601 net1_ota.n264 net1_ota.n263 0.028
R18602 net1_ota.n489 net1_ota.n485 0.027
R18603 net1_ota.n26 net1_ota.n25 0.026
R18604 net1_ota.n40 net1_ota.n39 0.026
R18605 net1_ota.n211 net1_ota.n210 0.026
R18606 net1_ota.n11 net1_ota.n10 0.026
R18607 net1_ota.n251 net1_ota.n250 0.026
R18608 net1_ota.n272 net1_ota.n271 0.026
R18609 net1_ota.n443 net1_ota.n442 0.026
R18610 net1_ota.n243 net1_ota.n242 0.026
R18611 net1_ota.n198 net1_ota.n197 0.024
R18612 net1_ota.n200 net1_ota.n199 0.024
R18613 net1_ota.n177 net1_ota.n176 0.024
R18614 net1_ota.n191 net1_ota.n190 0.024
R18615 net1_ota.n169 net1_ota.n168 0.024
R18616 net1_ota.n166 net1_ota.n165 0.024
R18617 net1_ota.n78 net1_ota.n77 0.024
R18618 net1_ota.n13 net1_ota.n12 0.024
R18619 net1_ota.n16 net1_ota.n15 0.024
R18620 net1_ota.n22 net1_ota.n21 0.024
R18621 net1_ota.n430 net1_ota.n429 0.024
R18622 net1_ota.n432 net1_ota.n431 0.024
R18623 net1_ota.n409 net1_ota.n408 0.024
R18624 net1_ota.n423 net1_ota.n422 0.024
R18625 net1_ota.n401 net1_ota.n400 0.024
R18626 net1_ota.n398 net1_ota.n397 0.024
R18627 net1_ota.n310 net1_ota.n309 0.024
R18628 net1_ota.n245 net1_ota.n244 0.024
R18629 net1_ota.n248 net1_ota.n247 0.024
R18630 net1_ota.n266 net1_ota.n265 0.024
R18631 net1_ota.n153 net1_ota.n152 0.024
R18632 net1_ota.n66 net1_ota.n65 0.024
R18633 net1_ota.n385 net1_ota.n384 0.024
R18634 net1_ota.n298 net1_ota.n297 0.024
R18635 net1_ota.n193 net1_ota.n192 0.023
R18636 net1_ota.n146 net1_ota.n131 0.023
R18637 net1_ota.n80 net1_ota.n79 0.023
R18638 net1_ota.n57 net1_ota.n56 0.023
R18639 net1_ota.n425 net1_ota.n424 0.023
R18640 net1_ota.n378 net1_ota.n363 0.023
R18641 net1_ota.n312 net1_ota.n311 0.023
R18642 net1_ota.n289 net1_ota.n288 0.023
R18643 net1_ota.n29 net1_ota.n28 0.022
R18644 net1_ota.n1 net1_ota.n0 0.022
R18645 net1_ota.n254 net1_ota.n253 0.022
R18646 net1_ota.n233 net1_ota.n232 0.022
R18647 net1_ota.n507 net1_ota.n502 0.02
R18648 net1_ota.n187 net1_ota.n177 0.02
R18649 net1_ota.n36 net1_ota.n35 0.02
R18650 net1_ota.n37 net1_ota.n36 0.02
R18651 net1_ota.n171 net1_ota.n167 0.02
R18652 net1_ota.n72 net1_ota.n60 0.02
R18653 net1_ota.n419 net1_ota.n409 0.02
R18654 net1_ota.n269 net1_ota.n268 0.02
R18655 net1_ota.n403 net1_ota.n399 0.02
R18656 net1_ota.n304 net1_ota.n292 0.02
R18657 net1_ota.n476 net1_ota.n472 0.018
R18658 net1_ota.n471 net1_ota.n470 0.018
R18659 net1_ota.n483 net1_ota.n482 0.018
R18660 net1_ota.n141 net1_ota.n136 0.018
R18661 net1_ota.n64 net1_ota.n63 0.018
R18662 net1_ota.n21 net1_ota.n20 0.018
R18663 net1_ota.n373 net1_ota.n368 0.018
R18664 net1_ota.n296 net1_ota.n295 0.018
R18665 net1_ota.n265 net1_ota.n264 0.018
R18666 net1_ota.n501 net1_ota.n500 0.017
R18667 net1_ota.n206 net1_ota.n198 0.017
R18668 net1_ota.n162 net1_ota.n150 0.017
R18669 net1_ota.n160 net1_ota.n159 0.017
R18670 net1_ota.n125 net1_ota.n124 0.017
R18671 net1_ota.n210 net1_ota.n209 0.017
R18672 net1_ota.n438 net1_ota.n430 0.017
R18673 net1_ota.n394 net1_ota.n382 0.017
R18674 net1_ota.n392 net1_ota.n391 0.017
R18675 net1_ota.n357 net1_ota.n356 0.017
R18676 net1_ota.n442 net1_ota.n441 0.017
R18677 net1_ota.n478 net1_ota.n466 0.015
R18678 net1_ota.n482 net1_ota.n481 0.015
R18679 net1_ota.n493 net1_ota.n492 0.015
R18680 net1_ota.n123 net1_ota.n122 0.015
R18681 net1_ota.n190 net1_ota.n189 0.015
R18682 net1_ota.n165 net1_ota.n164 0.015
R18683 net1_ota.n77 net1_ota.n76 0.015
R18684 net1_ota.n355 net1_ota.n354 0.015
R18685 net1_ota.n422 net1_ota.n421 0.015
R18686 net1_ota.n397 net1_ota.n396 0.015
R18687 net1_ota.n309 net1_ota.n308 0.015
R18688 net1_ota.n477 net1_ota.n476 0.013
R18689 net1_ota.n509 net1_ota.n494 0.013
R18690 net1_ota.n105 net1_ota.n104 0.013
R18691 net1_ota.n104 net1_ota.n103 0.013
R18692 net1_ota.n94 net1_ota.n93 0.013
R18693 net1_ota.n69 net1_ota.n64 0.013
R18694 net1_ota.n71 net1_ota.n70 0.013
R18695 net1_ota.n14 net1_ota.n13 0.013
R18696 net1_ota.n337 net1_ota.n336 0.013
R18697 net1_ota.n336 net1_ota.n335 0.013
R18698 net1_ota.n326 net1_ota.n325 0.013
R18699 net1_ota.n301 net1_ota.n296 0.013
R18700 net1_ota.n303 net1_ota.n302 0.013
R18701 net1_ota.n246 net1_ota.n245 0.013
R18702 net1_ota.n139 net1_ota.n138 0.012
R18703 net1_ota.n88 net1_ota.n87 0.012
R18704 net1_ota.n371 net1_ota.n370 0.012
R18705 net1_ota.n320 net1_ota.n319 0.012
R18706 net1_ota.n231 net1_ota.n230 0.012
R18707 net1_ota.n194 net1_ota.n193 0.012
R18708 net1_ota.n131 net1_ota.n130 0.012
R18709 net1_ota.n81 net1_ota.n80 0.012
R18710 net1_ota.n56 net1_ota.n55 0.012
R18711 net1_ota.n463 net1_ota.n462 0.012
R18712 net1_ota.n426 net1_ota.n425 0.012
R18713 net1_ota.n363 net1_ota.n362 0.012
R18714 net1_ota.n313 net1_ota.n312 0.012
R18715 net1_ota.n288 net1_ota.n287 0.012
R18716 net1_ota.n508 net1_ota.n507 0.011
R18717 net1_ota.n494 net1_ota.n493 0.011
R18718 net1_ota.n222 net1_ota.n221 0.011
R18719 net1_ota.n201 net1_ota.n200 0.011
R18720 net1_ota.n184 net1_ota.n183 0.011
R18721 net1_ota.n162 net1_ota.n161 0.011
R18722 net1_ota.n4 net1_ota.n3 0.011
R18723 net1_ota.n9 net1_ota.n6 0.011
R18724 net1_ota.n170 net1_ota.n169 0.011
R18725 net1_ota.n166 net1_ota.n163 0.011
R18726 net1_ota.n106 net1_ota.n97 0.011
R18727 net1_ota.n51 net1_ota.n50 0.011
R18728 net1_ota.n454 net1_ota.n453 0.011
R18729 net1_ota.n433 net1_ota.n432 0.011
R18730 net1_ota.n411 net1_ota.n410 0.011
R18731 net1_ota.n394 net1_ota.n393 0.011
R18732 net1_ota.n236 net1_ota.n235 0.011
R18733 net1_ota.n241 net1_ota.n238 0.011
R18734 net1_ota.n402 net1_ota.n401 0.011
R18735 net1_ota.n398 net1_ota.n395 0.011
R18736 net1_ota.n338 net1_ota.n329 0.011
R18737 net1_ota.n283 net1_ota.n282 0.011
R18738 net1_ota.n485 net1_ota.n480 0.009
R18739 net1_ota.n490 net1_ota.n489 0.009
R18740 net1_ota.n510 net1_ota.n491 0.009
R18741 net1_ota.n220 net1_ota.n219 0.009
R18742 net1_ota.n134 net1_ota.n133 0.009
R18743 net1_ota.n136 net1_ota.n135 0.009
R18744 net1_ota.n27 net1_ota.n26 0.009
R18745 net1_ota.n227 net1_ota.n226 0.009
R18746 net1_ota.n212 net1_ota.n211 0.009
R18747 net1_ota.n128 net1_ota.n117 0.009
R18748 net1_ota.n12 net1_ota.n11 0.009
R18749 net1_ota.n23 net1_ota.n22 0.009
R18750 net1_ota.n452 net1_ota.n451 0.009
R18751 net1_ota.n366 net1_ota.n365 0.009
R18752 net1_ota.n368 net1_ota.n367 0.009
R18753 net1_ota.n252 net1_ota.n251 0.009
R18754 net1_ota.n459 net1_ota.n458 0.009
R18755 net1_ota.n444 net1_ota.n443 0.009
R18756 net1_ota.n360 net1_ota.n349 0.009
R18757 net1_ota.n244 net1_ota.n243 0.009
R18758 net1_ota.n267 net1_ota.n266 0.009
R18759 net1_ota.n500 net1_ota.n497 0.007
R18760 net1_ota.n488 net1_ota.n487 0.007
R18761 net1_ota.n223 net1_ota.n222 0.007
R18762 net1_ota.n186 net1_ota.n185 0.007
R18763 net1_ota.n150 net1_ota.n149 0.007
R18764 net1_ota.n35 net1_ota.n30 0.007
R18765 net1_ota.n41 net1_ota.n40 0.007
R18766 net1_ota.n46 net1_ota.n41 0.007
R18767 net1_ota.n6 net1_ota.n5 0.007
R18768 net1_ota.n228 net1_ota.n224 0.007
R18769 net1_ota.n17 net1_ota.n16 0.007
R18770 net1_ota.n47 net1_ota.n23 0.007
R18771 net1_ota.n192 net1_ota.n173 0.007
R18772 net1_ota.n172 net1_ota.n171 0.007
R18773 net1_ota.n167 net1_ota.n148 0.007
R18774 net1_ota.n147 net1_ota.n146 0.007
R18775 net1_ota.n79 net1_ota.n74 0.007
R18776 net1_ota.n73 net1_ota.n72 0.007
R18777 net1_ota.n60 net1_ota.n59 0.007
R18778 net1_ota.n58 net1_ota.n57 0.007
R18779 net1_ota.n455 net1_ota.n454 0.007
R18780 net1_ota.n413 net1_ota.n412 0.007
R18781 net1_ota.n382 net1_ota.n381 0.007
R18782 net1_ota.n260 net1_ota.n255 0.007
R18783 net1_ota.n273 net1_ota.n272 0.007
R18784 net1_ota.n278 net1_ota.n273 0.007
R18785 net1_ota.n238 net1_ota.n237 0.007
R18786 net1_ota.n460 net1_ota.n456 0.007
R18787 net1_ota.n261 net1_ota.n248 0.007
R18788 net1_ota.n279 net1_ota.n267 0.007
R18789 net1_ota.n424 net1_ota.n405 0.007
R18790 net1_ota.n404 net1_ota.n403 0.007
R18791 net1_ota.n399 net1_ota.n380 0.007
R18792 net1_ota.n379 net1_ota.n378 0.007
R18793 net1_ota.n311 net1_ota.n306 0.007
R18794 net1_ota.n305 net1_ota.n304 0.007
R18795 net1_ota.n292 net1_ota.n291 0.007
R18796 net1_ota.n290 net1_ota.n289 0.007
R18797 net1_ota.n472 net1_ota.n471 0.005
R18798 net1_ota.n502 net1_ota.n501 0.005
R18799 net1_ota.n484 net1_ota.n483 0.005
R18800 net1_ota.n480 net1_ota.n479 0.005
R18801 net1_ota.n491 net1_ota.n490 0.005
R18802 net1_ota.n38 net1_ota.n37 0.005
R18803 net1_ota.n108 net1_ota.n107 0.005
R18804 net1_ota.n19 net1_ota.n18 0.005
R18805 net1_ota.n270 net1_ota.n269 0.005
R18806 net1_ota.n340 net1_ota.n339 0.005
R18807 net1_ota.n263 net1_ota.n262 0.005
R18808 net1_ota.n53 net1_ota.n52 0.004
R18809 net1_ota.n285 net1_ota.n284 0.004
R18810 net1_ota.n223 net1_ota.n218 0.004
R18811 net1_ota.n455 net1_ota.n450 0.004
R18812 net1_ota.n173 net1_ota.n172 0.004
R18813 net1_ota.n148 net1_ota.n147 0.004
R18814 net1_ota.n74 net1_ota.n73 0.004
R18815 net1_ota.n59 net1_ota.n58 0.004
R18816 net1_ota.n405 net1_ota.n404 0.004
R18817 net1_ota.n380 net1_ota.n379 0.004
R18818 net1_ota.n306 net1_ota.n305 0.004
R18819 net1_ota.n291 net1_ota.n290 0.004
R18820 net1_ota.n197 net1_ota.n196 0.003
R18821 net1_ota.n206 net1_ota.n201 0.003
R18822 net1_ota.n176 net1_ota.n175 0.003
R18823 net1_ota.n187 net1_ota.n186 0.003
R18824 net1_ota.n161 net1_ota.n160 0.003
R18825 net1_ota.n156 net1_ota.n155 0.003
R18826 net1_ota.n141 net1_ota.n134 0.003
R18827 net1_ota.n126 net1_ota.n125 0.003
R18828 net1_ota.n99 net1_ota.n98 0.003
R18829 net1_ota.n25 net1_ota.n24 0.003
R18830 net1_ota.n30 net1_ota.n29 0.003
R18831 net1_ota.n212 net1_ota.n207 0.003
R18832 net1_ota.n191 net1_ota.n188 0.003
R18833 net1_ota.n145 net1_ota.n144 0.003
R18834 net1_ota.n143 net1_ota.n142 0.003
R18835 net1_ota.n127 net1_ota.n119 0.003
R18836 net1_ota.n109 net1_ota.n108 0.003
R18837 net1_ota.n429 net1_ota.n428 0.003
R18838 net1_ota.n438 net1_ota.n433 0.003
R18839 net1_ota.n408 net1_ota.n407 0.003
R18840 net1_ota.n419 net1_ota.n413 0.003
R18841 net1_ota.n393 net1_ota.n392 0.003
R18842 net1_ota.n388 net1_ota.n387 0.003
R18843 net1_ota.n373 net1_ota.n366 0.003
R18844 net1_ota.n358 net1_ota.n357 0.003
R18845 net1_ota.n331 net1_ota.n330 0.003
R18846 net1_ota.n250 net1_ota.n249 0.003
R18847 net1_ota.n255 net1_ota.n254 0.003
R18848 net1_ota.n444 net1_ota.n439 0.003
R18849 net1_ota.n423 net1_ota.n420 0.003
R18850 net1_ota.n377 net1_ota.n376 0.003
R18851 net1_ota.n375 net1_ota.n374 0.003
R18852 net1_ota.n359 net1_ota.n351 0.003
R18853 net1_ota.n341 net1_ota.n340 0.003
R18854 net1_ota.n230 net1_ota.n229 0.002
R18855 net1_ota.n213 net1_ota.n194 0.002
R18856 net1_ota.n130 net1_ota.n129 0.002
R18857 net1_ota.n110 net1_ota.n81 0.002
R18858 net1_ota.n55 net1_ota.n54 0.002
R18859 net1_ota.n462 net1_ota.n461 0.002
R18860 net1_ota.n445 net1_ota.n426 0.002
R18861 net1_ota.n362 net1_ota.n361 0.002
R18862 net1_ota.n342 net1_ota.n313 0.002
R18863 net1_ota.n287 net1_ota.n286 0.002
R18864 net1_ota.n124 net1_ota.n123 0.001
R18865 net1_ota.n95 net1_ota.n94 0.001
R18866 net1_ota.n92 net1_ota.n91 0.001
R18867 net1_ota.n2 net1_ota.n1 0.001
R18868 net1_ota.n224 net1_ota.n215 0.001
R18869 net1_ota.n96 net1_ota.n86 0.001
R18870 net1_ota.n78 net1_ota.n75 0.001
R18871 net1_ota.n15 net1_ota.n14 0.001
R18872 net1_ota.n49 net1_ota.n48 0.001
R18873 net1_ota.n356 net1_ota.n355 0.001
R18874 net1_ota.n327 net1_ota.n326 0.001
R18875 net1_ota.n324 net1_ota.n323 0.001
R18876 net1_ota.n234 net1_ota.n233 0.001
R18877 net1_ota.n456 net1_ota.n447 0.001
R18878 net1_ota.n328 net1_ota.n318 0.001
R18879 net1_ota.n310 net1_ota.n307 0.001
R18880 net1_ota.n247 net1_ota.n246 0.001
R18881 net1_ota.n281 net1_ota.n280 0.001
R18882 net4.n1358 net4.t2 124.695
R18883 net4.n1337 net4.t5 124.695
R18884 net4.n1316 net4.t17 124.695
R18885 net4.n1295 net4.t0 124.695
R18886 net4.n1275 net4.t16 124.695
R18887 net4.n1251 net4.t1 124.695
R18888 net4.n1231 net4.t19 124.695
R18889 net4.n1211 net4.t18 124.695
R18890 net4.n1191 net4.t3 124.695
R18891 net4.n1171 net4.t4 124.695
R18892 net4.n1079 net4.n1078 92.5
R18893 net4.n1130 net4.n1129 92.5
R18894 net4.n962 net4.n961 92.5
R18895 net4.n1013 net4.n1012 92.5
R18896 net4.n845 net4.n844 92.5
R18897 net4.n896 net4.n895 92.5
R18898 net4.n728 net4.n727 92.5
R18899 net4.n779 net4.n778 92.5
R18900 net4.n611 net4.n610 92.5
R18901 net4.n662 net4.n661 92.5
R18902 net4.n494 net4.n493 92.5
R18903 net4.n545 net4.n544 92.5
R18904 net4.n377 net4.n376 92.5
R18905 net4.n428 net4.n427 92.5
R18906 net4.n260 net4.n259 92.5
R18907 net4.n311 net4.n310 92.5
R18908 net4.n143 net4.n142 92.5
R18909 net4.n194 net4.n193 92.5
R18910 net4.n15 net4.n14 92.5
R18911 net4.n78 net4.n77 92.5
R18912 net4.n1357 net4.n1356 92.5
R18913 net4.n1336 net4.n1335 92.5
R18914 net4.n1315 net4.n1314 92.5
R18915 net4.n1294 net4.n1293 92.5
R18916 net4.n1274 net4.n1273 92.5
R18917 net4.n1250 net4.n1249 92.5
R18918 net4.n1230 net4.n1229 92.5
R18919 net4.n1210 net4.n1209 92.5
R18920 net4.n1190 net4.n1189 92.5
R18921 net4.n1170 net4.n1169 92.5
R18922 net4.n1078 net4.t12 70.344
R18923 net4.n961 net4.t8 70.344
R18924 net4.n844 net4.t7 70.344
R18925 net4.n727 net4.t10 70.344
R18926 net4.n610 net4.t15 70.344
R18927 net4.n493 net4.t13 70.344
R18928 net4.n376 net4.t9 70.344
R18929 net4.n259 net4.t11 70.344
R18930 net4.n142 net4.t14 70.344
R18931 net4.n14 net4.t6 70.344
R18932 net4.n1069 net4.n1068 31.034
R18933 net4.n1147 net4.n1146 31.034
R18934 net4.n952 net4.n951 31.034
R18935 net4.n1030 net4.n1029 31.034
R18936 net4.n835 net4.n834 31.034
R18937 net4.n913 net4.n912 31.034
R18938 net4.n718 net4.n717 31.034
R18939 net4.n796 net4.n795 31.034
R18940 net4.n601 net4.n600 31.034
R18941 net4.n679 net4.n678 31.034
R18942 net4.n484 net4.n483 31.034
R18943 net4.n562 net4.n561 31.034
R18944 net4.n367 net4.n366 31.034
R18945 net4.n445 net4.n444 31.034
R18946 net4.n250 net4.n249 31.034
R18947 net4.n328 net4.n327 31.034
R18948 net4.n133 net4.n132 31.034
R18949 net4.n211 net4.n210 31.034
R18950 net4.n28 net4.n27 31.034
R18951 net4.n95 net4.n94 31.034
R18952 net4.n1367 net4.n1366 31.034
R18953 net4.n1346 net4.n1345 31.034
R18954 net4.n1325 net4.n1324 31.034
R18955 net4.n1304 net4.n1303 31.034
R18956 net4.n1284 net4.n1283 31.034
R18957 net4.n1260 net4.n1259 31.034
R18958 net4.n1240 net4.n1239 31.034
R18959 net4.n1220 net4.n1219 31.034
R18960 net4.n1200 net4.n1199 31.034
R18961 net4.n1180 net4.n1179 31.034
R18962 net4.n1358 net4.n1357 15.431
R18963 net4.n1337 net4.n1336 15.431
R18964 net4.n1316 net4.n1315 15.431
R18965 net4.n1295 net4.n1294 15.431
R18966 net4.n1275 net4.n1274 15.431
R18967 net4.n1251 net4.n1250 15.431
R18968 net4.n1231 net4.n1230 15.431
R18969 net4.n1211 net4.n1210 15.431
R18970 net4.n1191 net4.n1190 15.431
R18971 net4.n1171 net4.n1170 15.431
R18972 net4.n1090 net4.n1089 9.3
R18973 net4.n1070 net4.n1069 9.3
R18974 net4.n1148 net4.n1147 9.3
R18975 net4.n1156 net4.n1155 9.3
R18976 net4.n973 net4.n972 9.3
R18977 net4.n953 net4.n952 9.3
R18978 net4.n1031 net4.n1030 9.3
R18979 net4.n1039 net4.n1038 9.3
R18980 net4.n856 net4.n855 9.3
R18981 net4.n836 net4.n835 9.3
R18982 net4.n914 net4.n913 9.3
R18983 net4.n922 net4.n921 9.3
R18984 net4.n739 net4.n738 9.3
R18985 net4.n719 net4.n718 9.3
R18986 net4.n797 net4.n796 9.3
R18987 net4.n805 net4.n804 9.3
R18988 net4.n622 net4.n621 9.3
R18989 net4.n602 net4.n601 9.3
R18990 net4.n680 net4.n679 9.3
R18991 net4.n688 net4.n687 9.3
R18992 net4.n505 net4.n504 9.3
R18993 net4.n485 net4.n484 9.3
R18994 net4.n563 net4.n562 9.3
R18995 net4.n571 net4.n570 9.3
R18996 net4.n388 net4.n387 9.3
R18997 net4.n368 net4.n367 9.3
R18998 net4.n446 net4.n445 9.3
R18999 net4.n454 net4.n453 9.3
R19000 net4.n271 net4.n270 9.3
R19001 net4.n251 net4.n250 9.3
R19002 net4.n329 net4.n328 9.3
R19003 net4.n337 net4.n336 9.3
R19004 net4.n154 net4.n153 9.3
R19005 net4.n134 net4.n133 9.3
R19006 net4.n212 net4.n211 9.3
R19007 net4.n220 net4.n219 9.3
R19008 net4.n38 net4.n37 9.3
R19009 net4.n104 net4.n103 9.3
R19010 net4.n96 net4.n95 9.3
R19011 net4.n29 net4.n28 9.3
R19012 net4.n1373 net4.n1372 9.3
R19013 net4.n1362 net4.n1361 9.3
R19014 net4.n1360 net4.n1359 9.3
R19015 net4.n1369 net4.n1368 9.3
R19016 net4.n1368 net4.n1367 9.3
R19017 net4.n1371 net4.n1370 9.3
R19018 net4.n1375 net4.n1374 9.3
R19019 net4.n1352 net4.n1351 9.3
R19020 net4.n1341 net4.n1340 9.3
R19021 net4.n1339 net4.n1338 9.3
R19022 net4.n1348 net4.n1347 9.3
R19023 net4.n1347 net4.n1346 9.3
R19024 net4.n1350 net4.n1349 9.3
R19025 net4.n1354 net4.n1353 9.3
R19026 net4.n1331 net4.n1330 9.3
R19027 net4.n1320 net4.n1319 9.3
R19028 net4.n1318 net4.n1317 9.3
R19029 net4.n1327 net4.n1326 9.3
R19030 net4.n1326 net4.n1325 9.3
R19031 net4.n1329 net4.n1328 9.3
R19032 net4.n1333 net4.n1332 9.3
R19033 net4.n1310 net4.n1309 9.3
R19034 net4.n1299 net4.n1298 9.3
R19035 net4.n1297 net4.n1296 9.3
R19036 net4.n1306 net4.n1305 9.3
R19037 net4.n1305 net4.n1304 9.3
R19038 net4.n1308 net4.n1307 9.3
R19039 net4.n1312 net4.n1311 9.3
R19040 net4.n1290 net4.n1289 9.3
R19041 net4.n1279 net4.n1278 9.3
R19042 net4.n1277 net4.n1276 9.3
R19043 net4.n1286 net4.n1285 9.3
R19044 net4.n1285 net4.n1284 9.3
R19045 net4.n1288 net4.n1287 9.3
R19046 net4.n1292 net4.n1291 9.3
R19047 net4.n1266 net4.n1265 9.3
R19048 net4.n1255 net4.n1254 9.3
R19049 net4.n1253 net4.n1252 9.3
R19050 net4.n1262 net4.n1261 9.3
R19051 net4.n1261 net4.n1260 9.3
R19052 net4.n1264 net4.n1263 9.3
R19053 net4.n1268 net4.n1267 9.3
R19054 net4.n1246 net4.n1245 9.3
R19055 net4.n1235 net4.n1234 9.3
R19056 net4.n1233 net4.n1232 9.3
R19057 net4.n1242 net4.n1241 9.3
R19058 net4.n1241 net4.n1240 9.3
R19059 net4.n1244 net4.n1243 9.3
R19060 net4.n1248 net4.n1247 9.3
R19061 net4.n1226 net4.n1225 9.3
R19062 net4.n1215 net4.n1214 9.3
R19063 net4.n1213 net4.n1212 9.3
R19064 net4.n1222 net4.n1221 9.3
R19065 net4.n1221 net4.n1220 9.3
R19066 net4.n1224 net4.n1223 9.3
R19067 net4.n1228 net4.n1227 9.3
R19068 net4.n1206 net4.n1205 9.3
R19069 net4.n1195 net4.n1194 9.3
R19070 net4.n1193 net4.n1192 9.3
R19071 net4.n1202 net4.n1201 9.3
R19072 net4.n1201 net4.n1200 9.3
R19073 net4.n1204 net4.n1203 9.3
R19074 net4.n1208 net4.n1207 9.3
R19075 net4.n1186 net4.n1185 9.3
R19076 net4.n1175 net4.n1174 9.3
R19077 net4.n1173 net4.n1172 9.3
R19078 net4.n1182 net4.n1181 9.3
R19079 net4.n1181 net4.n1180 9.3
R19080 net4.n1184 net4.n1183 9.3
R19081 net4.n1188 net4.n1187 9.3
R19082 net4.n1080 net4.n1079 8.282
R19083 net4.n1131 net4.n1130 8.282
R19084 net4.n963 net4.n962 8.282
R19085 net4.n1014 net4.n1013 8.282
R19086 net4.n846 net4.n845 8.282
R19087 net4.n897 net4.n896 8.282
R19088 net4.n729 net4.n728 8.282
R19089 net4.n780 net4.n779 8.282
R19090 net4.n612 net4.n611 8.282
R19091 net4.n663 net4.n662 8.282
R19092 net4.n495 net4.n494 8.282
R19093 net4.n546 net4.n545 8.282
R19094 net4.n378 net4.n377 8.282
R19095 net4.n429 net4.n428 8.282
R19096 net4.n261 net4.n260 8.282
R19097 net4.n312 net4.n311 8.282
R19098 net4.n144 net4.n143 8.282
R19099 net4.n195 net4.n194 8.282
R19100 net4.n16 net4.n15 8.282
R19101 net4.n79 net4.n78 8.282
R19102 net4.n1070 net4.n1066 5.647
R19103 net4.n1148 net4.n1144 5.647
R19104 net4.n953 net4.n949 5.647
R19105 net4.n1031 net4.n1027 5.647
R19106 net4.n836 net4.n832 5.647
R19107 net4.n914 net4.n910 5.647
R19108 net4.n719 net4.n715 5.647
R19109 net4.n797 net4.n793 5.647
R19110 net4.n602 net4.n598 5.647
R19111 net4.n680 net4.n676 5.647
R19112 net4.n485 net4.n481 5.647
R19113 net4.n563 net4.n559 5.647
R19114 net4.n368 net4.n364 5.647
R19115 net4.n446 net4.n442 5.647
R19116 net4.n251 net4.n247 5.647
R19117 net4.n329 net4.n325 5.647
R19118 net4.n134 net4.n130 5.647
R19119 net4.n212 net4.n208 5.647
R19120 net4.n29 net4.n25 5.647
R19121 net4.n96 net4.n92 5.647
R19122 net4.n1368 net4.n1364 5.647
R19123 net4.n1347 net4.n1343 5.647
R19124 net4.n1326 net4.n1322 5.647
R19125 net4.n1305 net4.n1301 5.647
R19126 net4.n1285 net4.n1281 5.647
R19127 net4.n1261 net4.n1257 5.647
R19128 net4.n1241 net4.n1237 5.647
R19129 net4.n1221 net4.n1217 5.647
R19130 net4.n1201 net4.n1197 5.647
R19131 net4.n1181 net4.n1177 5.647
R19132 net4.n1128 net4.n1127 4.65
R19133 net4.n1011 net4.n1010 4.65
R19134 net4.n894 net4.n893 4.65
R19135 net4.n777 net4.n776 4.65
R19136 net4.n660 net4.n659 4.65
R19137 net4.n543 net4.n542 4.65
R19138 net4.n426 net4.n425 4.65
R19139 net4.n309 net4.n308 4.65
R19140 net4.n192 net4.n191 4.65
R19141 net4.n76 net4.n75 4.65
R19142 net4.n1162 net4.n1160 4.5
R19143 net4.n1150 net4.n1149 4.5
R19144 net4.n1139 net4.n1138 4.5
R19145 net4.n1132 net4.n1131 4.5
R19146 net4.n1084 net4.n1072 4.5
R19147 net4.n1081 net4.n1080 4.5
R19148 net4.n1126 net4.n1125 4.5
R19149 net4.n1095 net4.n1094 4.5
R19150 net4.n1045 net4.n1043 4.5
R19151 net4.n1033 net4.n1032 4.5
R19152 net4.n1022 net4.n1021 4.5
R19153 net4.n1015 net4.n1014 4.5
R19154 net4.n967 net4.n955 4.5
R19155 net4.n964 net4.n963 4.5
R19156 net4.n1009 net4.n1008 4.5
R19157 net4.n978 net4.n977 4.5
R19158 net4.n928 net4.n926 4.5
R19159 net4.n916 net4.n915 4.5
R19160 net4.n905 net4.n904 4.5
R19161 net4.n898 net4.n897 4.5
R19162 net4.n850 net4.n838 4.5
R19163 net4.n847 net4.n846 4.5
R19164 net4.n892 net4.n891 4.5
R19165 net4.n861 net4.n860 4.5
R19166 net4.n811 net4.n809 4.5
R19167 net4.n799 net4.n798 4.5
R19168 net4.n788 net4.n787 4.5
R19169 net4.n781 net4.n780 4.5
R19170 net4.n733 net4.n721 4.5
R19171 net4.n730 net4.n729 4.5
R19172 net4.n775 net4.n774 4.5
R19173 net4.n744 net4.n743 4.5
R19174 net4.n694 net4.n692 4.5
R19175 net4.n682 net4.n681 4.5
R19176 net4.n671 net4.n670 4.5
R19177 net4.n664 net4.n663 4.5
R19178 net4.n616 net4.n604 4.5
R19179 net4.n613 net4.n612 4.5
R19180 net4.n658 net4.n657 4.5
R19181 net4.n627 net4.n626 4.5
R19182 net4.n577 net4.n575 4.5
R19183 net4.n565 net4.n564 4.5
R19184 net4.n554 net4.n553 4.5
R19185 net4.n547 net4.n546 4.5
R19186 net4.n499 net4.n487 4.5
R19187 net4.n496 net4.n495 4.5
R19188 net4.n541 net4.n540 4.5
R19189 net4.n510 net4.n509 4.5
R19190 net4.n460 net4.n458 4.5
R19191 net4.n448 net4.n447 4.5
R19192 net4.n437 net4.n436 4.5
R19193 net4.n430 net4.n429 4.5
R19194 net4.n382 net4.n370 4.5
R19195 net4.n379 net4.n378 4.5
R19196 net4.n424 net4.n423 4.5
R19197 net4.n393 net4.n392 4.5
R19198 net4.n343 net4.n341 4.5
R19199 net4.n331 net4.n330 4.5
R19200 net4.n320 net4.n319 4.5
R19201 net4.n313 net4.n312 4.5
R19202 net4.n265 net4.n253 4.5
R19203 net4.n262 net4.n261 4.5
R19204 net4.n307 net4.n306 4.5
R19205 net4.n276 net4.n275 4.5
R19206 net4.n226 net4.n224 4.5
R19207 net4.n214 net4.n213 4.5
R19208 net4.n203 net4.n202 4.5
R19209 net4.n196 net4.n195 4.5
R19210 net4.n148 net4.n136 4.5
R19211 net4.n145 net4.n144 4.5
R19212 net4.n190 net4.n189 4.5
R19213 net4.n159 net4.n158 4.5
R19214 net4.n80 net4.n79 4.5
R19215 net4.n87 net4.n86 4.5
R19216 net4.n21 net4.n16 4.5
R19217 net4.n98 net4.n97 4.5
R19218 net4.n74 net4.n73 4.5
R19219 net4.n32 net4.n31 4.5
R19220 net4.n110 net4.n108 4.5
R19221 net4.n43 net4.n42 4.5
R19222 net4.n1068 net4.n1067 4.137
R19223 net4.n1146 net4.n1145 4.137
R19224 net4.n951 net4.n950 4.137
R19225 net4.n1029 net4.n1028 4.137
R19226 net4.n834 net4.n833 4.137
R19227 net4.n912 net4.n911 4.137
R19228 net4.n717 net4.n716 4.137
R19229 net4.n795 net4.n794 4.137
R19230 net4.n600 net4.n599 4.137
R19231 net4.n678 net4.n677 4.137
R19232 net4.n483 net4.n482 4.137
R19233 net4.n561 net4.n560 4.137
R19234 net4.n366 net4.n365 4.137
R19235 net4.n444 net4.n443 4.137
R19236 net4.n249 net4.n248 4.137
R19237 net4.n327 net4.n326 4.137
R19238 net4.n132 net4.n131 4.137
R19239 net4.n210 net4.n209 4.137
R19240 net4.n27 net4.n26 4.137
R19241 net4.n94 net4.n93 4.137
R19242 net4.n1366 net4.n1365 4.137
R19243 net4.n1345 net4.n1344 4.137
R19244 net4.n1324 net4.n1323 4.137
R19245 net4.n1303 net4.n1302 4.137
R19246 net4.n1283 net4.n1282 4.137
R19247 net4.n1259 net4.n1258 4.137
R19248 net4.n1239 net4.n1238 4.137
R19249 net4.n1219 net4.n1218 4.137
R19250 net4.n1199 net4.n1198 4.137
R19251 net4.n1179 net4.n1178 4.137
R19252 net4.n1094 net4.n1092 3.764
R19253 net4.n1149 net4.n1142 3.764
R19254 net4.n977 net4.n975 3.764
R19255 net4.n1032 net4.n1025 3.764
R19256 net4.n860 net4.n858 3.764
R19257 net4.n915 net4.n908 3.764
R19258 net4.n743 net4.n741 3.764
R19259 net4.n798 net4.n791 3.764
R19260 net4.n626 net4.n624 3.764
R19261 net4.n681 net4.n674 3.764
R19262 net4.n509 net4.n507 3.764
R19263 net4.n564 net4.n557 3.764
R19264 net4.n392 net4.n390 3.764
R19265 net4.n447 net4.n440 3.764
R19266 net4.n275 net4.n273 3.764
R19267 net4.n330 net4.n323 3.764
R19268 net4.n158 net4.n156 3.764
R19269 net4.n213 net4.n206 3.764
R19270 net4.n42 net4.n40 3.764
R19271 net4.n97 net4.n90 3.764
R19272 net4.n1072 net4.n1071 3.388
R19273 net4.n1160 net4.n1159 3.388
R19274 net4.n955 net4.n954 3.388
R19275 net4.n1043 net4.n1042 3.388
R19276 net4.n838 net4.n837 3.388
R19277 net4.n926 net4.n925 3.388
R19278 net4.n721 net4.n720 3.388
R19279 net4.n809 net4.n808 3.388
R19280 net4.n604 net4.n603 3.388
R19281 net4.n692 net4.n691 3.388
R19282 net4.n487 net4.n486 3.388
R19283 net4.n575 net4.n574 3.388
R19284 net4.n370 net4.n369 3.388
R19285 net4.n458 net4.n457 3.388
R19286 net4.n253 net4.n252 3.388
R19287 net4.n341 net4.n340 3.388
R19288 net4.n136 net4.n135 3.388
R19289 net4.n224 net4.n223 3.388
R19290 net4.n31 net4.n30 3.388
R19291 net4.n108 net4.n107 3.388
R19292 net4.n1072 net4.n1070 3.011
R19293 net4.n1080 net4.n1077 3.011
R19294 net4.n1160 net4.n1158 3.011
R19295 net4.n955 net4.n953 3.011
R19296 net4.n963 net4.n960 3.011
R19297 net4.n1043 net4.n1041 3.011
R19298 net4.n838 net4.n836 3.011
R19299 net4.n846 net4.n843 3.011
R19300 net4.n926 net4.n924 3.011
R19301 net4.n721 net4.n719 3.011
R19302 net4.n729 net4.n726 3.011
R19303 net4.n809 net4.n807 3.011
R19304 net4.n604 net4.n602 3.011
R19305 net4.n612 net4.n609 3.011
R19306 net4.n692 net4.n690 3.011
R19307 net4.n487 net4.n485 3.011
R19308 net4.n495 net4.n492 3.011
R19309 net4.n575 net4.n573 3.011
R19310 net4.n370 net4.n368 3.011
R19311 net4.n378 net4.n375 3.011
R19312 net4.n458 net4.n456 3.011
R19313 net4.n253 net4.n251 3.011
R19314 net4.n261 net4.n258 3.011
R19315 net4.n341 net4.n339 3.011
R19316 net4.n136 net4.n134 3.011
R19317 net4.n144 net4.n141 3.011
R19318 net4.n224 net4.n222 3.011
R19319 net4.n31 net4.n29 3.011
R19320 net4.n16 net4.n13 3.011
R19321 net4.n108 net4.n106 3.011
R19322 net4.n1094 net4.n1093 2.635
R19323 net4.n1138 net4.n1137 2.635
R19324 net4.n1149 net4.n1148 2.635
R19325 net4.n977 net4.n976 2.635
R19326 net4.n1021 net4.n1020 2.635
R19327 net4.n1032 net4.n1031 2.635
R19328 net4.n860 net4.n859 2.635
R19329 net4.n904 net4.n903 2.635
R19330 net4.n915 net4.n914 2.635
R19331 net4.n743 net4.n742 2.635
R19332 net4.n787 net4.n786 2.635
R19333 net4.n798 net4.n797 2.635
R19334 net4.n626 net4.n625 2.635
R19335 net4.n670 net4.n669 2.635
R19336 net4.n681 net4.n680 2.635
R19337 net4.n509 net4.n508 2.635
R19338 net4.n553 net4.n552 2.635
R19339 net4.n564 net4.n563 2.635
R19340 net4.n392 net4.n391 2.635
R19341 net4.n436 net4.n435 2.635
R19342 net4.n447 net4.n446 2.635
R19343 net4.n275 net4.n274 2.635
R19344 net4.n319 net4.n318 2.635
R19345 net4.n330 net4.n329 2.635
R19346 net4.n158 net4.n157 2.635
R19347 net4.n202 net4.n201 2.635
R19348 net4.n213 net4.n212 2.635
R19349 net4.n42 net4.n41 2.635
R19350 net4.n86 net4.n85 2.635
R19351 net4.n97 net4.n96 2.635
R19352 net4.n1313 net4.n1292 2.04
R19353 net4.n1269 net4.n1268 2.04
R19354 net4.n1272 net4.n1188 1.826
R19355 net4.n1271 net4.n1208 1.826
R19356 net4.n1270 net4.n1228 1.826
R19357 net4.n1269 net4.n1248 1.826
R19358 net4.n1313 net4.n1312 1.826
R19359 net4.n1355 net4.n1354 1.826
R19360 net4.n1376 net4.n1375 1.824
R19361 net4.n1334 net4.n1333 1.824
R19362 net4.n1360 net4.n1358 1.57
R19363 net4.n1339 net4.n1337 1.57
R19364 net4.n1318 net4.n1316 1.57
R19365 net4.n1297 net4.n1295 1.57
R19366 net4.n1277 net4.n1275 1.57
R19367 net4.n1253 net4.n1251 1.57
R19368 net4.n1233 net4.n1231 1.57
R19369 net4.n1213 net4.n1211 1.57
R19370 net4.n1193 net4.n1191 1.57
R19371 net4.n1173 net4.n1171 1.57
R19372 net4.n1163 net4.n1162 1.5
R19373 net4.n1096 net4.n1095 1.5
R19374 net4.n1046 net4.n1045 1.5
R19375 net4.n979 net4.n978 1.5
R19376 net4.n929 net4.n928 1.5
R19377 net4.n862 net4.n861 1.5
R19378 net4.n812 net4.n811 1.5
R19379 net4.n745 net4.n744 1.5
R19380 net4.n695 net4.n694 1.5
R19381 net4.n628 net4.n627 1.5
R19382 net4.n578 net4.n577 1.5
R19383 net4.n511 net4.n510 1.5
R19384 net4.n461 net4.n460 1.5
R19385 net4.n394 net4.n393 1.5
R19386 net4.n344 net4.n343 1.5
R19387 net4.n277 net4.n276 1.5
R19388 net4.n227 net4.n226 1.5
R19389 net4.n160 net4.n159 1.5
R19390 net4.n111 net4.n110 1.5
R19391 net4.n44 net4.n43 1.5
R19392 net4 net4.n1377 1.033
R19393 net4.n232 net4.n115 0.972
R19394 net4.n1051 net4.n1050 0.923
R19395 net4.n1168 net4.n1167 0.921
R19396 net4.n934 net4.n933 0.921
R19397 net4.n817 net4.n816 0.918
R19398 net4.n583 net4.n582 0.918
R19399 net4.n349 net4.n348 0.918
R19400 net4.n700 net4.n699 0.916
R19401 net4.n466 net4.n465 0.916
R19402 net4.n232 net4.n231 0.916
R19403 net4.n1166 net4.n1165 0.853
R19404 net4.n1049 net4.n1048 0.853
R19405 net4.n932 net4.n931 0.853
R19406 net4.n815 net4.n814 0.853
R19407 net4.n698 net4.n697 0.853
R19408 net4.n581 net4.n580 0.853
R19409 net4.n464 net4.n463 0.853
R19410 net4.n347 net4.n346 0.853
R19411 net4.n230 net4.n229 0.853
R19412 net4.n114 net4.n113 0.853
R19413 net4.n1066 net4.n1065 0.752
R19414 net4.n1144 net4.n1143 0.752
R19415 net4.n949 net4.n948 0.752
R19416 net4.n1027 net4.n1026 0.752
R19417 net4.n832 net4.n831 0.752
R19418 net4.n910 net4.n909 0.752
R19419 net4.n715 net4.n714 0.752
R19420 net4.n793 net4.n792 0.752
R19421 net4.n598 net4.n597 0.752
R19422 net4.n676 net4.n675 0.752
R19423 net4.n481 net4.n480 0.752
R19424 net4.n559 net4.n558 0.752
R19425 net4.n364 net4.n363 0.752
R19426 net4.n442 net4.n441 0.752
R19427 net4.n247 net4.n246 0.752
R19428 net4.n325 net4.n324 0.752
R19429 net4.n130 net4.n129 0.752
R19430 net4.n208 net4.n207 0.752
R19431 net4.n25 net4.n24 0.752
R19432 net4.n92 net4.n91 0.752
R19433 net4.n1364 net4.n1363 0.752
R19434 net4.n1343 net4.n1342 0.752
R19435 net4.n1322 net4.n1321 0.752
R19436 net4.n1301 net4.n1300 0.752
R19437 net4.n1281 net4.n1280 0.752
R19438 net4.n1257 net4.n1256 0.752
R19439 net4.n1237 net4.n1236 0.752
R19440 net4.n1217 net4.n1216 0.752
R19441 net4.n1197 net4.n1196 0.752
R19442 net4.n1177 net4.n1176 0.752
R19443 net4.n46 net4.n45 0.704
R19444 net4.n1098 net4.n1097 0.702
R19445 net4.n981 net4.n980 0.702
R19446 net4.n864 net4.n863 0.702
R19447 net4.n747 net4.n746 0.702
R19448 net4.n630 net4.n629 0.702
R19449 net4.n513 net4.n512 0.702
R19450 net4.n396 net4.n395 0.702
R19451 net4.n279 net4.n278 0.702
R19452 net4.n162 net4.n161 0.702
R19453 net4.n1334 net4.n1313 0.432
R19454 net4.n1355 net4.n1334 0.432
R19455 net4.n1271 net4.n1270 0.432
R19456 net4.n1270 net4.n1269 0.432
R19457 net4 net4.n1168 0.313
R19458 net4.n1377 net4.n1272 0.228
R19459 net4.n1376 net4.n1355 0.216
R19460 net4.n1272 net4.n1271 0.216
R19461 net4.n1377 net4.n1376 0.203
R19462 net4.n1371 net4.n1369 0.144
R19463 net4.n1350 net4.n1348 0.144
R19464 net4.n1329 net4.n1327 0.144
R19465 net4.n1308 net4.n1306 0.144
R19466 net4.n1288 net4.n1286 0.144
R19467 net4.n1264 net4.n1262 0.144
R19468 net4.n1244 net4.n1242 0.144
R19469 net4.n1224 net4.n1222 0.144
R19470 net4.n1204 net4.n1202 0.144
R19471 net4.n1184 net4.n1182 0.144
R19472 net4.n700 net4.n583 0.114
R19473 net4.n934 net4.n817 0.113
R19474 net4.n466 net4.n349 0.113
R19475 net4.n1168 net4.n1051 0.056
R19476 net4.n1051 net4.n934 0.056
R19477 net4.n817 net4.n700 0.056
R19478 net4.n583 net4.n466 0.056
R19479 net4.n349 net4.n232 0.056
R19480 net4.n1369 net4.n1362 0.04
R19481 net4.n1348 net4.n1341 0.04
R19482 net4.n1327 net4.n1320 0.04
R19483 net4.n1306 net4.n1299 0.04
R19484 net4.n1286 net4.n1279 0.04
R19485 net4.n1262 net4.n1255 0.04
R19486 net4.n1242 net4.n1235 0.04
R19487 net4.n1222 net4.n1215 0.04
R19488 net4.n1202 net4.n1195 0.04
R19489 net4.n1182 net4.n1175 0.04
R19490 net4.n1074 net4.n1073 0.035
R19491 net4.n1134 net4.n1133 0.035
R19492 net4.n1053 net4.n1052 0.035
R19493 net4.n1115 net4.n1114 0.035
R19494 net4.n957 net4.n956 0.035
R19495 net4.n1017 net4.n1016 0.035
R19496 net4.n936 net4.n935 0.035
R19497 net4.n998 net4.n997 0.035
R19498 net4.n840 net4.n839 0.035
R19499 net4.n900 net4.n899 0.035
R19500 net4.n819 net4.n818 0.035
R19501 net4.n881 net4.n880 0.035
R19502 net4.n723 net4.n722 0.035
R19503 net4.n783 net4.n782 0.035
R19504 net4.n702 net4.n701 0.035
R19505 net4.n764 net4.n763 0.035
R19506 net4.n606 net4.n605 0.035
R19507 net4.n666 net4.n665 0.035
R19508 net4.n585 net4.n584 0.035
R19509 net4.n647 net4.n646 0.035
R19510 net4.n489 net4.n488 0.035
R19511 net4.n549 net4.n548 0.035
R19512 net4.n468 net4.n467 0.035
R19513 net4.n530 net4.n529 0.035
R19514 net4.n372 net4.n371 0.035
R19515 net4.n432 net4.n431 0.035
R19516 net4.n351 net4.n350 0.035
R19517 net4.n413 net4.n412 0.035
R19518 net4.n255 net4.n254 0.035
R19519 net4.n315 net4.n314 0.035
R19520 net4.n234 net4.n233 0.035
R19521 net4.n296 net4.n295 0.035
R19522 net4.n138 net4.n137 0.035
R19523 net4.n198 net4.n197 0.035
R19524 net4.n117 net4.n116 0.035
R19525 net4.n179 net4.n178 0.035
R19526 net4.n18 net4.n17 0.035
R19527 net4.n82 net4.n81 0.035
R19528 net4.n1 net4.n0 0.035
R19529 net4.n63 net4.n62 0.035
R19530 net4.n1375 net4.n1373 0.035
R19531 net4.n1354 net4.n1352 0.035
R19532 net4.n1333 net4.n1331 0.035
R19533 net4.n1312 net4.n1310 0.035
R19534 net4.n1292 net4.n1290 0.035
R19535 net4.n1268 net4.n1266 0.035
R19536 net4.n1248 net4.n1246 0.035
R19537 net4.n1228 net4.n1226 0.035
R19538 net4.n1208 net4.n1206 0.035
R19539 net4.n1188 net4.n1186 0.035
R19540 net4.n1063 net4.n1062 0.034
R19541 net4.n1124 net4.n1123 0.034
R19542 net4.n946 net4.n945 0.034
R19543 net4.n1007 net4.n1006 0.034
R19544 net4.n829 net4.n828 0.034
R19545 net4.n890 net4.n889 0.034
R19546 net4.n712 net4.n711 0.034
R19547 net4.n773 net4.n772 0.034
R19548 net4.n595 net4.n594 0.034
R19549 net4.n656 net4.n655 0.034
R19550 net4.n478 net4.n477 0.034
R19551 net4.n539 net4.n538 0.034
R19552 net4.n361 net4.n360 0.034
R19553 net4.n422 net4.n421 0.034
R19554 net4.n244 net4.n243 0.034
R19555 net4.n305 net4.n304 0.034
R19556 net4.n127 net4.n126 0.034
R19557 net4.n188 net4.n187 0.034
R19558 net4.n11 net4.n10 0.034
R19559 net4.n72 net4.n71 0.034
R19560 net4.n1153 net4.n1152 0.032
R19561 net4.n1122 net4.n1121 0.032
R19562 net4.n1036 net4.n1035 0.032
R19563 net4.n1005 net4.n1004 0.032
R19564 net4.n919 net4.n918 0.032
R19565 net4.n888 net4.n887 0.032
R19566 net4.n802 net4.n801 0.032
R19567 net4.n771 net4.n770 0.032
R19568 net4.n685 net4.n684 0.032
R19569 net4.n654 net4.n653 0.032
R19570 net4.n568 net4.n567 0.032
R19571 net4.n537 net4.n536 0.032
R19572 net4.n451 net4.n450 0.032
R19573 net4.n420 net4.n419 0.032
R19574 net4.n334 net4.n333 0.032
R19575 net4.n303 net4.n302 0.032
R19576 net4.n217 net4.n216 0.032
R19577 net4.n186 net4.n185 0.032
R19578 net4.n101 net4.n100 0.032
R19579 net4.n70 net4.n69 0.032
R19580 net4.n1099 net4.n1098 0.031
R19581 net4.n1110 net4.n1109 0.031
R19582 net4.n982 net4.n981 0.031
R19583 net4.n993 net4.n992 0.031
R19584 net4.n865 net4.n864 0.031
R19585 net4.n876 net4.n875 0.031
R19586 net4.n748 net4.n747 0.031
R19587 net4.n759 net4.n758 0.031
R19588 net4.n631 net4.n630 0.031
R19589 net4.n642 net4.n641 0.031
R19590 net4.n514 net4.n513 0.031
R19591 net4.n525 net4.n524 0.031
R19592 net4.n397 net4.n396 0.031
R19593 net4.n408 net4.n407 0.031
R19594 net4.n280 net4.n279 0.031
R19595 net4.n291 net4.n290 0.031
R19596 net4.n163 net4.n162 0.031
R19597 net4.n174 net4.n173 0.031
R19598 net4.n47 net4.n46 0.031
R19599 net4.n58 net4.n57 0.031
R19600 net4.n1087 net4.n1086 0.03
R19601 net4.n1156 net4.n1154 0.03
R19602 net4.n1061 net4.n1060 0.03
R19603 net4.n1120 net4.n1119 0.03
R19604 net4.n970 net4.n969 0.03
R19605 net4.n1039 net4.n1037 0.03
R19606 net4.n944 net4.n943 0.03
R19607 net4.n1003 net4.n1002 0.03
R19608 net4.n853 net4.n852 0.03
R19609 net4.n922 net4.n920 0.03
R19610 net4.n827 net4.n826 0.03
R19611 net4.n886 net4.n885 0.03
R19612 net4.n736 net4.n735 0.03
R19613 net4.n805 net4.n803 0.03
R19614 net4.n710 net4.n709 0.03
R19615 net4.n769 net4.n768 0.03
R19616 net4.n619 net4.n618 0.03
R19617 net4.n688 net4.n686 0.03
R19618 net4.n593 net4.n592 0.03
R19619 net4.n652 net4.n651 0.03
R19620 net4.n502 net4.n501 0.03
R19621 net4.n571 net4.n569 0.03
R19622 net4.n476 net4.n475 0.03
R19623 net4.n535 net4.n534 0.03
R19624 net4.n385 net4.n384 0.03
R19625 net4.n454 net4.n452 0.03
R19626 net4.n359 net4.n358 0.03
R19627 net4.n418 net4.n417 0.03
R19628 net4.n268 net4.n267 0.03
R19629 net4.n337 net4.n335 0.03
R19630 net4.n242 net4.n241 0.03
R19631 net4.n301 net4.n300 0.03
R19632 net4.n151 net4.n150 0.03
R19633 net4.n220 net4.n218 0.03
R19634 net4.n125 net4.n124 0.03
R19635 net4.n184 net4.n183 0.03
R19636 net4.n35 net4.n34 0.03
R19637 net4.n104 net4.n102 0.03
R19638 net4.n9 net4.n8 0.03
R19639 net4.n68 net4.n67 0.03
R19640 net4.n1090 net4.n1088 0.028
R19641 net4.n1076 net4.n1075 0.028
R19642 net4.n1136 net4.n1135 0.028
R19643 net4.n1058 net4.n1057 0.028
R19644 net4.n1055 net4.n1054 0.028
R19645 net4.n1117 net4.n1116 0.028
R19646 net4.n1163 net4.n1124 0.028
R19647 net4.n973 net4.n971 0.028
R19648 net4.n959 net4.n958 0.028
R19649 net4.n1019 net4.n1018 0.028
R19650 net4.n941 net4.n940 0.028
R19651 net4.n938 net4.n937 0.028
R19652 net4.n1000 net4.n999 0.028
R19653 net4.n1046 net4.n1007 0.028
R19654 net4.n856 net4.n854 0.028
R19655 net4.n842 net4.n841 0.028
R19656 net4.n902 net4.n901 0.028
R19657 net4.n824 net4.n823 0.028
R19658 net4.n821 net4.n820 0.028
R19659 net4.n883 net4.n882 0.028
R19660 net4.n929 net4.n890 0.028
R19661 net4.n739 net4.n737 0.028
R19662 net4.n725 net4.n724 0.028
R19663 net4.n785 net4.n784 0.028
R19664 net4.n707 net4.n706 0.028
R19665 net4.n704 net4.n703 0.028
R19666 net4.n766 net4.n765 0.028
R19667 net4.n812 net4.n773 0.028
R19668 net4.n622 net4.n620 0.028
R19669 net4.n608 net4.n607 0.028
R19670 net4.n668 net4.n667 0.028
R19671 net4.n590 net4.n589 0.028
R19672 net4.n587 net4.n586 0.028
R19673 net4.n649 net4.n648 0.028
R19674 net4.n695 net4.n656 0.028
R19675 net4.n505 net4.n503 0.028
R19676 net4.n491 net4.n490 0.028
R19677 net4.n551 net4.n550 0.028
R19678 net4.n473 net4.n472 0.028
R19679 net4.n470 net4.n469 0.028
R19680 net4.n532 net4.n531 0.028
R19681 net4.n578 net4.n539 0.028
R19682 net4.n388 net4.n386 0.028
R19683 net4.n374 net4.n373 0.028
R19684 net4.n434 net4.n433 0.028
R19685 net4.n356 net4.n355 0.028
R19686 net4.n353 net4.n352 0.028
R19687 net4.n415 net4.n414 0.028
R19688 net4.n461 net4.n422 0.028
R19689 net4.n271 net4.n269 0.028
R19690 net4.n257 net4.n256 0.028
R19691 net4.n317 net4.n316 0.028
R19692 net4.n239 net4.n238 0.028
R19693 net4.n236 net4.n235 0.028
R19694 net4.n298 net4.n297 0.028
R19695 net4.n344 net4.n305 0.028
R19696 net4.n154 net4.n152 0.028
R19697 net4.n140 net4.n139 0.028
R19698 net4.n200 net4.n199 0.028
R19699 net4.n122 net4.n121 0.028
R19700 net4.n119 net4.n118 0.028
R19701 net4.n181 net4.n180 0.028
R19702 net4.n227 net4.n188 0.028
R19703 net4.n38 net4.n36 0.028
R19704 net4.n20 net4.n19 0.028
R19705 net4.n84 net4.n83 0.028
R19706 net4.n6 net4.n5 0.028
R19707 net4.n3 net4.n2 0.028
R19708 net4.n65 net4.n64 0.028
R19709 net4.n111 net4.n72 0.028
R19710 net4.n1097 net4.n1096 0.028
R19711 net4.n980 net4.n979 0.028
R19712 net4.n863 net4.n862 0.028
R19713 net4.n746 net4.n745 0.028
R19714 net4.n629 net4.n628 0.028
R19715 net4.n512 net4.n511 0.028
R19716 net4.n395 net4.n394 0.028
R19717 net4.n278 net4.n277 0.028
R19718 net4.n161 net4.n160 0.028
R19719 net4.n45 net4.n44 0.027
R19720 net4.n1103 net4.n1102 0.027
R19721 net4.n1106 net4.n1105 0.027
R19722 net4.n986 net4.n985 0.027
R19723 net4.n989 net4.n988 0.027
R19724 net4.n869 net4.n868 0.027
R19725 net4.n872 net4.n871 0.027
R19726 net4.n752 net4.n751 0.027
R19727 net4.n755 net4.n754 0.027
R19728 net4.n635 net4.n634 0.027
R19729 net4.n638 net4.n637 0.027
R19730 net4.n518 net4.n517 0.027
R19731 net4.n521 net4.n520 0.027
R19732 net4.n401 net4.n400 0.027
R19733 net4.n404 net4.n403 0.027
R19734 net4.n284 net4.n283 0.027
R19735 net4.n287 net4.n286 0.027
R19736 net4.n167 net4.n166 0.027
R19737 net4.n170 net4.n169 0.027
R19738 net4.n51 net4.n50 0.027
R19739 net4.n54 net4.n53 0.027
R19740 net4.n1096 net4.n1063 0.026
R19741 net4.n979 net4.n946 0.026
R19742 net4.n862 net4.n829 0.026
R19743 net4.n745 net4.n712 0.026
R19744 net4.n628 net4.n595 0.026
R19745 net4.n511 net4.n478 0.026
R19746 net4.n394 net4.n361 0.026
R19747 net4.n277 net4.n244 0.026
R19748 net4.n160 net4.n127 0.026
R19749 net4.n44 net4.n11 0.026
R19750 net4.n1132 net4.n1128 0.022
R19751 net4.n1113 net4.n1112 0.022
R19752 net4.n1165 net4.n1163 0.022
R19753 net4.n1015 net4.n1011 0.022
R19754 net4.n996 net4.n995 0.022
R19755 net4.n1048 net4.n1046 0.022
R19756 net4.n898 net4.n894 0.022
R19757 net4.n879 net4.n878 0.022
R19758 net4.n931 net4.n929 0.022
R19759 net4.n781 net4.n777 0.022
R19760 net4.n762 net4.n761 0.022
R19761 net4.n814 net4.n812 0.022
R19762 net4.n664 net4.n660 0.022
R19763 net4.n645 net4.n644 0.022
R19764 net4.n697 net4.n695 0.022
R19765 net4.n547 net4.n543 0.022
R19766 net4.n528 net4.n527 0.022
R19767 net4.n580 net4.n578 0.022
R19768 net4.n430 net4.n426 0.022
R19769 net4.n411 net4.n410 0.022
R19770 net4.n463 net4.n461 0.022
R19771 net4.n313 net4.n309 0.022
R19772 net4.n294 net4.n293 0.022
R19773 net4.n346 net4.n344 0.022
R19774 net4.n196 net4.n192 0.022
R19775 net4.n177 net4.n176 0.022
R19776 net4.n229 net4.n227 0.022
R19777 net4.n80 net4.n76 0.022
R19778 net4.n61 net4.n60 0.022
R19779 net4.n113 net4.n111 0.022
R19780 net4.n1128 net4.n1126 0.02
R19781 net4.n1112 net4.n1111 0.02
R19782 net4.n1011 net4.n1009 0.02
R19783 net4.n995 net4.n994 0.02
R19784 net4.n894 net4.n892 0.02
R19785 net4.n878 net4.n877 0.02
R19786 net4.n777 net4.n775 0.02
R19787 net4.n761 net4.n760 0.02
R19788 net4.n660 net4.n658 0.02
R19789 net4.n644 net4.n643 0.02
R19790 net4.n543 net4.n541 0.02
R19791 net4.n527 net4.n526 0.02
R19792 net4.n426 net4.n424 0.02
R19793 net4.n410 net4.n409 0.02
R19794 net4.n309 net4.n307 0.02
R19795 net4.n293 net4.n292 0.02
R19796 net4.n192 net4.n190 0.02
R19797 net4.n176 net4.n175 0.02
R19798 net4.n76 net4.n74 0.02
R19799 net4.n60 net4.n59 0.02
R19800 net4.n1166 net4.n1110 0.019
R19801 net4.n1167 net4.n1166 0.019
R19802 net4.n1049 net4.n993 0.019
R19803 net4.n1050 net4.n1049 0.019
R19804 net4.n932 net4.n876 0.019
R19805 net4.n933 net4.n932 0.019
R19806 net4.n815 net4.n759 0.019
R19807 net4.n816 net4.n815 0.019
R19808 net4.n698 net4.n642 0.019
R19809 net4.n699 net4.n698 0.019
R19810 net4.n581 net4.n525 0.019
R19811 net4.n582 net4.n581 0.019
R19812 net4.n464 net4.n408 0.019
R19813 net4.n465 net4.n464 0.019
R19814 net4.n347 net4.n291 0.019
R19815 net4.n348 net4.n347 0.019
R19816 net4.n230 net4.n174 0.019
R19817 net4.n231 net4.n230 0.019
R19818 net4.n114 net4.n58 0.019
R19819 net4.n115 net4.n114 0.019
R19820 net4.n1095 net4.n1064 0.018
R19821 net4.n1091 net4.n1090 0.018
R19822 net4.n1088 net4.n1087 0.018
R19823 net4.n1150 net4.n1141 0.018
R19824 net4.n1062 net4.n1061 0.018
R19825 net4.n978 net4.n947 0.018
R19826 net4.n974 net4.n973 0.018
R19827 net4.n971 net4.n970 0.018
R19828 net4.n1033 net4.n1024 0.018
R19829 net4.n945 net4.n944 0.018
R19830 net4.n861 net4.n830 0.018
R19831 net4.n857 net4.n856 0.018
R19832 net4.n854 net4.n853 0.018
R19833 net4.n916 net4.n907 0.018
R19834 net4.n828 net4.n827 0.018
R19835 net4.n744 net4.n713 0.018
R19836 net4.n740 net4.n739 0.018
R19837 net4.n737 net4.n736 0.018
R19838 net4.n799 net4.n790 0.018
R19839 net4.n711 net4.n710 0.018
R19840 net4.n627 net4.n596 0.018
R19841 net4.n623 net4.n622 0.018
R19842 net4.n620 net4.n619 0.018
R19843 net4.n682 net4.n673 0.018
R19844 net4.n594 net4.n593 0.018
R19845 net4.n510 net4.n479 0.018
R19846 net4.n506 net4.n505 0.018
R19847 net4.n503 net4.n502 0.018
R19848 net4.n565 net4.n556 0.018
R19849 net4.n477 net4.n476 0.018
R19850 net4.n393 net4.n362 0.018
R19851 net4.n389 net4.n388 0.018
R19852 net4.n386 net4.n385 0.018
R19853 net4.n448 net4.n439 0.018
R19854 net4.n360 net4.n359 0.018
R19855 net4.n276 net4.n245 0.018
R19856 net4.n272 net4.n271 0.018
R19857 net4.n269 net4.n268 0.018
R19858 net4.n331 net4.n322 0.018
R19859 net4.n243 net4.n242 0.018
R19860 net4.n159 net4.n128 0.018
R19861 net4.n155 net4.n154 0.018
R19862 net4.n152 net4.n151 0.018
R19863 net4.n214 net4.n205 0.018
R19864 net4.n126 net4.n125 0.018
R19865 net4.n43 net4.n12 0.018
R19866 net4.n39 net4.n38 0.018
R19867 net4.n36 net4.n35 0.018
R19868 net4.n98 net4.n89 0.018
R19869 net4.n10 net4.n9 0.018
R19870 net4.n1084 net4.n1083 0.017
R19871 net4.n1154 net4.n1153 0.017
R19872 net4.n1157 net4.n1156 0.017
R19873 net4.n1162 net4.n1161 0.017
R19874 net4.n1060 net4.n1059 0.017
R19875 net4.n1121 net4.n1120 0.017
R19876 net4.n1123 net4.n1122 0.017
R19877 net4.n967 net4.n966 0.017
R19878 net4.n1037 net4.n1036 0.017
R19879 net4.n1040 net4.n1039 0.017
R19880 net4.n1045 net4.n1044 0.017
R19881 net4.n943 net4.n942 0.017
R19882 net4.n1004 net4.n1003 0.017
R19883 net4.n1006 net4.n1005 0.017
R19884 net4.n850 net4.n849 0.017
R19885 net4.n920 net4.n919 0.017
R19886 net4.n923 net4.n922 0.017
R19887 net4.n928 net4.n927 0.017
R19888 net4.n826 net4.n825 0.017
R19889 net4.n887 net4.n886 0.017
R19890 net4.n889 net4.n888 0.017
R19891 net4.n733 net4.n732 0.017
R19892 net4.n803 net4.n802 0.017
R19893 net4.n806 net4.n805 0.017
R19894 net4.n811 net4.n810 0.017
R19895 net4.n709 net4.n708 0.017
R19896 net4.n770 net4.n769 0.017
R19897 net4.n772 net4.n771 0.017
R19898 net4.n616 net4.n615 0.017
R19899 net4.n686 net4.n685 0.017
R19900 net4.n689 net4.n688 0.017
R19901 net4.n694 net4.n693 0.017
R19902 net4.n592 net4.n591 0.017
R19903 net4.n653 net4.n652 0.017
R19904 net4.n655 net4.n654 0.017
R19905 net4.n499 net4.n498 0.017
R19906 net4.n569 net4.n568 0.017
R19907 net4.n572 net4.n571 0.017
R19908 net4.n577 net4.n576 0.017
R19909 net4.n475 net4.n474 0.017
R19910 net4.n536 net4.n535 0.017
R19911 net4.n538 net4.n537 0.017
R19912 net4.n382 net4.n381 0.017
R19913 net4.n452 net4.n451 0.017
R19914 net4.n455 net4.n454 0.017
R19915 net4.n460 net4.n459 0.017
R19916 net4.n358 net4.n357 0.017
R19917 net4.n419 net4.n418 0.017
R19918 net4.n421 net4.n420 0.017
R19919 net4.n265 net4.n264 0.017
R19920 net4.n335 net4.n334 0.017
R19921 net4.n338 net4.n337 0.017
R19922 net4.n343 net4.n342 0.017
R19923 net4.n241 net4.n240 0.017
R19924 net4.n302 net4.n301 0.017
R19925 net4.n304 net4.n303 0.017
R19926 net4.n148 net4.n147 0.017
R19927 net4.n218 net4.n217 0.017
R19928 net4.n221 net4.n220 0.017
R19929 net4.n226 net4.n225 0.017
R19930 net4.n124 net4.n123 0.017
R19931 net4.n185 net4.n184 0.017
R19932 net4.n187 net4.n186 0.017
R19933 net4.n32 net4.n23 0.017
R19934 net4.n102 net4.n101 0.017
R19935 net4.n105 net4.n104 0.017
R19936 net4.n110 net4.n109 0.017
R19937 net4.n8 net4.n7 0.017
R19938 net4.n69 net4.n68 0.017
R19939 net4.n71 net4.n70 0.017
R19940 net4.n1085 net4.n1084 0.015
R19941 net4.n1082 net4.n1081 0.015
R19942 net4.n1162 net4.n1157 0.015
R19943 net4.n1057 net4.n1056 0.015
R19944 net4.n968 net4.n967 0.015
R19945 net4.n965 net4.n964 0.015
R19946 net4.n1045 net4.n1040 0.015
R19947 net4.n940 net4.n939 0.015
R19948 net4.n851 net4.n850 0.015
R19949 net4.n848 net4.n847 0.015
R19950 net4.n928 net4.n923 0.015
R19951 net4.n823 net4.n822 0.015
R19952 net4.n734 net4.n733 0.015
R19953 net4.n731 net4.n730 0.015
R19954 net4.n811 net4.n806 0.015
R19955 net4.n706 net4.n705 0.015
R19956 net4.n617 net4.n616 0.015
R19957 net4.n614 net4.n613 0.015
R19958 net4.n694 net4.n689 0.015
R19959 net4.n589 net4.n588 0.015
R19960 net4.n500 net4.n499 0.015
R19961 net4.n497 net4.n496 0.015
R19962 net4.n577 net4.n572 0.015
R19963 net4.n472 net4.n471 0.015
R19964 net4.n383 net4.n382 0.015
R19965 net4.n380 net4.n379 0.015
R19966 net4.n460 net4.n455 0.015
R19967 net4.n355 net4.n354 0.015
R19968 net4.n266 net4.n265 0.015
R19969 net4.n263 net4.n262 0.015
R19970 net4.n343 net4.n338 0.015
R19971 net4.n238 net4.n237 0.015
R19972 net4.n149 net4.n148 0.015
R19973 net4.n146 net4.n145 0.015
R19974 net4.n226 net4.n221 0.015
R19975 net4.n121 net4.n120 0.015
R19976 net4.n33 net4.n32 0.015
R19977 net4.n22 net4.n21 0.015
R19978 net4.n110 net4.n105 0.015
R19979 net4.n5 net4.n4 0.015
R19980 net4.n1095 net4.n1091 0.013
R19981 net4.n1140 net4.n1139 0.013
R19982 net4.n1151 net4.n1150 0.013
R19983 net4.n1119 net4.n1118 0.013
R19984 net4.n978 net4.n974 0.013
R19985 net4.n1023 net4.n1022 0.013
R19986 net4.n1034 net4.n1033 0.013
R19987 net4.n1002 net4.n1001 0.013
R19988 net4.n861 net4.n857 0.013
R19989 net4.n906 net4.n905 0.013
R19990 net4.n917 net4.n916 0.013
R19991 net4.n885 net4.n884 0.013
R19992 net4.n744 net4.n740 0.013
R19993 net4.n789 net4.n788 0.013
R19994 net4.n800 net4.n799 0.013
R19995 net4.n768 net4.n767 0.013
R19996 net4.n627 net4.n623 0.013
R19997 net4.n672 net4.n671 0.013
R19998 net4.n683 net4.n682 0.013
R19999 net4.n651 net4.n650 0.013
R20000 net4.n510 net4.n506 0.013
R20001 net4.n555 net4.n554 0.013
R20002 net4.n566 net4.n565 0.013
R20003 net4.n534 net4.n533 0.013
R20004 net4.n393 net4.n389 0.013
R20005 net4.n438 net4.n437 0.013
R20006 net4.n449 net4.n448 0.013
R20007 net4.n417 net4.n416 0.013
R20008 net4.n276 net4.n272 0.013
R20009 net4.n321 net4.n320 0.013
R20010 net4.n332 net4.n331 0.013
R20011 net4.n300 net4.n299 0.013
R20012 net4.n159 net4.n155 0.013
R20013 net4.n204 net4.n203 0.013
R20014 net4.n215 net4.n214 0.013
R20015 net4.n183 net4.n182 0.013
R20016 net4.n43 net4.n39 0.013
R20017 net4.n88 net4.n87 0.013
R20018 net4.n99 net4.n98 0.013
R20019 net4.n67 net4.n66 0.013
R20020 net4.n1104 net4.n1103 0.012
R20021 net4.n1105 net4.n1104 0.012
R20022 net4.n987 net4.n986 0.012
R20023 net4.n988 net4.n987 0.012
R20024 net4.n870 net4.n869 0.012
R20025 net4.n871 net4.n870 0.012
R20026 net4.n753 net4.n752 0.012
R20027 net4.n754 net4.n753 0.012
R20028 net4.n636 net4.n635 0.012
R20029 net4.n637 net4.n636 0.012
R20030 net4.n519 net4.n518 0.012
R20031 net4.n520 net4.n519 0.012
R20032 net4.n402 net4.n401 0.012
R20033 net4.n403 net4.n402 0.012
R20034 net4.n285 net4.n284 0.012
R20035 net4.n286 net4.n285 0.012
R20036 net4.n168 net4.n167 0.012
R20037 net4.n169 net4.n168 0.012
R20038 net4.n52 net4.n51 0.012
R20039 net4.n53 net4.n52 0.012
R20040 net4.n1165 net4.n1164 0.012
R20041 net4.n1048 net4.n1047 0.012
R20042 net4.n931 net4.n930 0.012
R20043 net4.n814 net4.n813 0.012
R20044 net4.n697 net4.n696 0.012
R20045 net4.n580 net4.n579 0.012
R20046 net4.n463 net4.n462 0.012
R20047 net4.n346 net4.n345 0.012
R20048 net4.n229 net4.n228 0.012
R20049 net4.n113 net4.n112 0.012
R20050 net4.n1083 net4.n1082 0.011
R20051 net4.n1141 net4.n1140 0.011
R20052 net4.n1101 net4.n1100 0.011
R20053 net4.n1108 net4.n1107 0.011
R20054 net4.n966 net4.n965 0.011
R20055 net4.n1024 net4.n1023 0.011
R20056 net4.n984 net4.n983 0.011
R20057 net4.n991 net4.n990 0.011
R20058 net4.n849 net4.n848 0.011
R20059 net4.n907 net4.n906 0.011
R20060 net4.n867 net4.n866 0.011
R20061 net4.n874 net4.n873 0.011
R20062 net4.n732 net4.n731 0.011
R20063 net4.n790 net4.n789 0.011
R20064 net4.n750 net4.n749 0.011
R20065 net4.n757 net4.n756 0.011
R20066 net4.n615 net4.n614 0.011
R20067 net4.n673 net4.n672 0.011
R20068 net4.n633 net4.n632 0.011
R20069 net4.n640 net4.n639 0.011
R20070 net4.n498 net4.n497 0.011
R20071 net4.n556 net4.n555 0.011
R20072 net4.n516 net4.n515 0.011
R20073 net4.n523 net4.n522 0.011
R20074 net4.n381 net4.n380 0.011
R20075 net4.n439 net4.n438 0.011
R20076 net4.n399 net4.n398 0.011
R20077 net4.n406 net4.n405 0.011
R20078 net4.n264 net4.n263 0.011
R20079 net4.n322 net4.n321 0.011
R20080 net4.n282 net4.n281 0.011
R20081 net4.n289 net4.n288 0.011
R20082 net4.n147 net4.n146 0.011
R20083 net4.n205 net4.n204 0.011
R20084 net4.n165 net4.n164 0.011
R20085 net4.n172 net4.n171 0.011
R20086 net4.n23 net4.n22 0.011
R20087 net4.n89 net4.n88 0.011
R20088 net4.n49 net4.n48 0.011
R20089 net4.n56 net4.n55 0.011
R20090 net4.n1373 net4.n1371 0.01
R20091 net4.n1352 net4.n1350 0.01
R20092 net4.n1331 net4.n1329 0.01
R20093 net4.n1310 net4.n1308 0.01
R20094 net4.n1290 net4.n1288 0.01
R20095 net4.n1266 net4.n1264 0.01
R20096 net4.n1246 net4.n1244 0.01
R20097 net4.n1226 net4.n1224 0.01
R20098 net4.n1206 net4.n1204 0.01
R20099 net4.n1186 net4.n1184 0.01
R20100 net4.n1133 net4.n1132 0.009
R20101 net4.n1114 net4.n1113 0.009
R20102 net4.n1016 net4.n1015 0.009
R20103 net4.n997 net4.n996 0.009
R20104 net4.n899 net4.n898 0.009
R20105 net4.n880 net4.n879 0.009
R20106 net4.n782 net4.n781 0.009
R20107 net4.n763 net4.n762 0.009
R20108 net4.n665 net4.n664 0.009
R20109 net4.n646 net4.n645 0.009
R20110 net4.n548 net4.n547 0.009
R20111 net4.n529 net4.n528 0.009
R20112 net4.n431 net4.n430 0.009
R20113 net4.n412 net4.n411 0.009
R20114 net4.n314 net4.n313 0.009
R20115 net4.n295 net4.n294 0.009
R20116 net4.n197 net4.n196 0.009
R20117 net4.n178 net4.n177 0.009
R20118 net4.n81 net4.n80 0.009
R20119 net4.n62 net4.n61 0.009
R20120 net4.n1075 net4.n1074 0.007
R20121 net4.n1135 net4.n1134 0.007
R20122 net4.n1054 net4.n1053 0.007
R20123 net4.n1116 net4.n1115 0.007
R20124 net4.n958 net4.n957 0.007
R20125 net4.n1018 net4.n1017 0.007
R20126 net4.n937 net4.n936 0.007
R20127 net4.n999 net4.n998 0.007
R20128 net4.n841 net4.n840 0.007
R20129 net4.n901 net4.n900 0.007
R20130 net4.n820 net4.n819 0.007
R20131 net4.n882 net4.n881 0.007
R20132 net4.n724 net4.n723 0.007
R20133 net4.n784 net4.n783 0.007
R20134 net4.n703 net4.n702 0.007
R20135 net4.n765 net4.n764 0.007
R20136 net4.n607 net4.n606 0.007
R20137 net4.n667 net4.n666 0.007
R20138 net4.n586 net4.n585 0.007
R20139 net4.n648 net4.n647 0.007
R20140 net4.n490 net4.n489 0.007
R20141 net4.n550 net4.n549 0.007
R20142 net4.n469 net4.n468 0.007
R20143 net4.n531 net4.n530 0.007
R20144 net4.n373 net4.n372 0.007
R20145 net4.n433 net4.n432 0.007
R20146 net4.n352 net4.n351 0.007
R20147 net4.n414 net4.n413 0.007
R20148 net4.n256 net4.n255 0.007
R20149 net4.n316 net4.n315 0.007
R20150 net4.n235 net4.n234 0.007
R20151 net4.n297 net4.n296 0.007
R20152 net4.n139 net4.n138 0.007
R20153 net4.n199 net4.n198 0.007
R20154 net4.n118 net4.n117 0.007
R20155 net4.n180 net4.n179 0.007
R20156 net4.n19 net4.n18 0.007
R20157 net4.n83 net4.n82 0.007
R20158 net4.n2 net4.n1 0.007
R20159 net4.n64 net4.n63 0.007
R20160 net4.n1100 net4.n1099 0.006
R20161 net4.n1102 net4.n1101 0.006
R20162 net4.n1107 net4.n1106 0.006
R20163 net4.n1109 net4.n1108 0.006
R20164 net4.n983 net4.n982 0.006
R20165 net4.n985 net4.n984 0.006
R20166 net4.n990 net4.n989 0.006
R20167 net4.n992 net4.n991 0.006
R20168 net4.n866 net4.n865 0.006
R20169 net4.n868 net4.n867 0.006
R20170 net4.n873 net4.n872 0.006
R20171 net4.n875 net4.n874 0.006
R20172 net4.n749 net4.n748 0.006
R20173 net4.n751 net4.n750 0.006
R20174 net4.n756 net4.n755 0.006
R20175 net4.n758 net4.n757 0.006
R20176 net4.n632 net4.n631 0.006
R20177 net4.n634 net4.n633 0.006
R20178 net4.n639 net4.n638 0.006
R20179 net4.n641 net4.n640 0.006
R20180 net4.n515 net4.n514 0.006
R20181 net4.n517 net4.n516 0.006
R20182 net4.n522 net4.n521 0.006
R20183 net4.n524 net4.n523 0.006
R20184 net4.n398 net4.n397 0.006
R20185 net4.n400 net4.n399 0.006
R20186 net4.n405 net4.n404 0.006
R20187 net4.n407 net4.n406 0.006
R20188 net4.n281 net4.n280 0.006
R20189 net4.n283 net4.n282 0.006
R20190 net4.n288 net4.n287 0.006
R20191 net4.n290 net4.n289 0.006
R20192 net4.n164 net4.n163 0.006
R20193 net4.n166 net4.n165 0.006
R20194 net4.n171 net4.n170 0.006
R20195 net4.n173 net4.n172 0.006
R20196 net4.n48 net4.n47 0.006
R20197 net4.n50 net4.n49 0.006
R20198 net4.n55 net4.n54 0.006
R20199 net4.n57 net4.n56 0.006
R20200 net4.n1362 net4.n1360 0.005
R20201 net4.n1341 net4.n1339 0.005
R20202 net4.n1320 net4.n1318 0.005
R20203 net4.n1299 net4.n1297 0.005
R20204 net4.n1279 net4.n1277 0.005
R20205 net4.n1255 net4.n1253 0.005
R20206 net4.n1235 net4.n1233 0.005
R20207 net4.n1215 net4.n1213 0.005
R20208 net4.n1195 net4.n1193 0.005
R20209 net4.n1175 net4.n1173 0.005
R20210 net4.n1086 net4.n1085 0.003
R20211 net4.n1139 net4.n1136 0.003
R20212 net4.n1152 net4.n1151 0.003
R20213 net4.n1118 net4.n1117 0.003
R20214 net4.n969 net4.n968 0.003
R20215 net4.n1022 net4.n1019 0.003
R20216 net4.n1035 net4.n1034 0.003
R20217 net4.n1001 net4.n1000 0.003
R20218 net4.n852 net4.n851 0.003
R20219 net4.n905 net4.n902 0.003
R20220 net4.n918 net4.n917 0.003
R20221 net4.n884 net4.n883 0.003
R20222 net4.n735 net4.n734 0.003
R20223 net4.n788 net4.n785 0.003
R20224 net4.n801 net4.n800 0.003
R20225 net4.n767 net4.n766 0.003
R20226 net4.n618 net4.n617 0.003
R20227 net4.n671 net4.n668 0.003
R20228 net4.n684 net4.n683 0.003
R20229 net4.n650 net4.n649 0.003
R20230 net4.n501 net4.n500 0.003
R20231 net4.n554 net4.n551 0.003
R20232 net4.n567 net4.n566 0.003
R20233 net4.n533 net4.n532 0.003
R20234 net4.n384 net4.n383 0.003
R20235 net4.n437 net4.n434 0.003
R20236 net4.n450 net4.n449 0.003
R20237 net4.n416 net4.n415 0.003
R20238 net4.n267 net4.n266 0.003
R20239 net4.n320 net4.n317 0.003
R20240 net4.n333 net4.n332 0.003
R20241 net4.n299 net4.n298 0.003
R20242 net4.n150 net4.n149 0.003
R20243 net4.n203 net4.n200 0.003
R20244 net4.n216 net4.n215 0.003
R20245 net4.n182 net4.n181 0.003
R20246 net4.n34 net4.n33 0.003
R20247 net4.n87 net4.n84 0.003
R20248 net4.n100 net4.n99 0.003
R20249 net4.n66 net4.n65 0.003
R20250 net4.n1081 net4.n1076 0.001
R20251 net4.n1059 net4.n1058 0.001
R20252 net4.n1056 net4.n1055 0.001
R20253 net4.n964 net4.n959 0.001
R20254 net4.n942 net4.n941 0.001
R20255 net4.n939 net4.n938 0.001
R20256 net4.n847 net4.n842 0.001
R20257 net4.n825 net4.n824 0.001
R20258 net4.n822 net4.n821 0.001
R20259 net4.n730 net4.n725 0.001
R20260 net4.n708 net4.n707 0.001
R20261 net4.n705 net4.n704 0.001
R20262 net4.n613 net4.n608 0.001
R20263 net4.n591 net4.n590 0.001
R20264 net4.n588 net4.n587 0.001
R20265 net4.n496 net4.n491 0.001
R20266 net4.n474 net4.n473 0.001
R20267 net4.n471 net4.n470 0.001
R20268 net4.n379 net4.n374 0.001
R20269 net4.n357 net4.n356 0.001
R20270 net4.n354 net4.n353 0.001
R20271 net4.n262 net4.n257 0.001
R20272 net4.n240 net4.n239 0.001
R20273 net4.n237 net4.n236 0.001
R20274 net4.n145 net4.n140 0.001
R20275 net4.n123 net4.n122 0.001
R20276 net4.n120 net4.n119 0.001
R20277 net4.n21 net4.n20 0.001
R20278 net4.n7 net4.n6 0.001
R20279 net4.n4 net4.n3 0.001
R20280 net5.n29 net5.t4 124.695
R20281 net5.n70 net5.t2 124.695
R20282 net5.n9 net5.t3 124.695
R20283 net5.n92 net5.t5 124.695
R20284 net5.n196 net5.t7 124.695
R20285 net5.n175 net5.t6 124.695
R20286 net5.n154 net5.t8 124.695
R20287 net5.n133 net5.t10 124.695
R20288 net5.n113 net5.t9 124.695
R20289 net5.n49 net5.t1 124.695
R20290 net5.n28 net5.n27 92.5
R20291 net5.n69 net5.n68 92.5
R20292 net5.n8 net5.n7 92.5
R20293 net5.n91 net5.n90 92.5
R20294 net5.n195 net5.n194 92.5
R20295 net5.n174 net5.n173 92.5
R20296 net5.n153 net5.n152 92.5
R20297 net5.n132 net5.n131 92.5
R20298 net5.n112 net5.n111 92.5
R20299 net5.n48 net5.n47 92.5
R20300 net5.n38 net5.n37 31.034
R20301 net5.n79 net5.n78 31.034
R20302 net5.n18 net5.n17 31.034
R20303 net5.n101 net5.n100 31.034
R20304 net5.n205 net5.n204 31.034
R20305 net5.n184 net5.n183 31.034
R20306 net5.n163 net5.n162 31.034
R20307 net5.n142 net5.n141 31.034
R20308 net5.n122 net5.n121 31.034
R20309 net5.n58 net5.n57 31.034
R20310 net5.n29 net5.n28 15.431
R20311 net5.n70 net5.n69 15.431
R20312 net5.n9 net5.n8 15.431
R20313 net5.n92 net5.n91 15.431
R20314 net5.n196 net5.n195 15.431
R20315 net5.n175 net5.n174 15.431
R20316 net5.n154 net5.n153 15.431
R20317 net5.n133 net5.n132 15.431
R20318 net5.n113 net5.n112 15.431
R20319 net5.n49 net5.n48 15.431
R20320 net5.n44 net5.n43 9.3
R20321 net5.n33 net5.n32 9.3
R20322 net5.n31 net5.n30 9.3
R20323 net5.n40 net5.n39 9.3
R20324 net5.n39 net5.n38 9.3
R20325 net5.n42 net5.n41 9.3
R20326 net5.n46 net5.n45 9.3
R20327 net5.n85 net5.n84 9.3
R20328 net5.n74 net5.n73 9.3
R20329 net5.n72 net5.n71 9.3
R20330 net5.n81 net5.n80 9.3
R20331 net5.n80 net5.n79 9.3
R20332 net5.n83 net5.n82 9.3
R20333 net5.n87 net5.n86 9.3
R20334 net5.n24 net5.n23 9.3
R20335 net5.n13 net5.n12 9.3
R20336 net5.n11 net5.n10 9.3
R20337 net5.n20 net5.n19 9.3
R20338 net5.n19 net5.n18 9.3
R20339 net5.n22 net5.n21 9.3
R20340 net5.n26 net5.n25 9.3
R20341 net5.n107 net5.n106 9.3
R20342 net5.n96 net5.n95 9.3
R20343 net5.n94 net5.n93 9.3
R20344 net5.n103 net5.n102 9.3
R20345 net5.n102 net5.n101 9.3
R20346 net5.n105 net5.n104 9.3
R20347 net5.n109 net5.n108 9.3
R20348 net5.n211 net5.n210 9.3
R20349 net5.n200 net5.n199 9.3
R20350 net5.n198 net5.n197 9.3
R20351 net5.n207 net5.n206 9.3
R20352 net5.n206 net5.n205 9.3
R20353 net5.n209 net5.n208 9.3
R20354 net5.n213 net5.n212 9.3
R20355 net5.n190 net5.n189 9.3
R20356 net5.n179 net5.n178 9.3
R20357 net5.n177 net5.n176 9.3
R20358 net5.n186 net5.n185 9.3
R20359 net5.n185 net5.n184 9.3
R20360 net5.n188 net5.n187 9.3
R20361 net5.n192 net5.n191 9.3
R20362 net5.n169 net5.n168 9.3
R20363 net5.n158 net5.n157 9.3
R20364 net5.n156 net5.n155 9.3
R20365 net5.n165 net5.n164 9.3
R20366 net5.n164 net5.n163 9.3
R20367 net5.n167 net5.n166 9.3
R20368 net5.n171 net5.n170 9.3
R20369 net5.n148 net5.n147 9.3
R20370 net5.n137 net5.n136 9.3
R20371 net5.n135 net5.n134 9.3
R20372 net5.n144 net5.n143 9.3
R20373 net5.n143 net5.n142 9.3
R20374 net5.n146 net5.n145 9.3
R20375 net5.n150 net5.n149 9.3
R20376 net5.n128 net5.n127 9.3
R20377 net5.n117 net5.n116 9.3
R20378 net5.n115 net5.n114 9.3
R20379 net5.n124 net5.n123 9.3
R20380 net5.n123 net5.n122 9.3
R20381 net5.n126 net5.n125 9.3
R20382 net5.n130 net5.n129 9.3
R20383 net5.n62 net5.n61 9.3
R20384 net5.n53 net5.n52 9.3
R20385 net5.n51 net5.n50 9.3
R20386 net5.n60 net5.n59 9.3
R20387 net5.n59 net5.n58 9.3
R20388 net5.n64 net5.n63 9.3
R20389 net5.n66 net5.n65 9.3
R20390 net5.n2 net5.t0 7.863
R20391 net5.n0 net5.t11 7.863
R20392 net5.n39 net5.n35 5.647
R20393 net5.n80 net5.n76 5.647
R20394 net5.n19 net5.n15 5.647
R20395 net5.n102 net5.n98 5.647
R20396 net5.n206 net5.n202 5.647
R20397 net5.n185 net5.n181 5.647
R20398 net5.n164 net5.n160 5.647
R20399 net5.n143 net5.n139 5.647
R20400 net5.n123 net5.n119 5.647
R20401 net5.n59 net5.n55 5.647
R20402 net5.n37 net5.n36 4.137
R20403 net5.n78 net5.n77 4.137
R20404 net5.n17 net5.n16 4.137
R20405 net5.n100 net5.n99 4.137
R20406 net5.n204 net5.n203 4.137
R20407 net5.n183 net5.n182 4.137
R20408 net5.n162 net5.n161 4.137
R20409 net5.n141 net5.n140 4.137
R20410 net5.n121 net5.n120 4.137
R20411 net5.n57 net5.n56 4.137
R20412 net5.n67 net5.n66 2.043
R20413 net5.n151 net5.n130 2.041
R20414 net5.n151 net5.n150 1.826
R20415 net5.n193 net5.n192 1.826
R20416 net5.n89 net5.n26 1.826
R20417 net5.n67 net5.n46 1.826
R20418 net5.n88 net5.n87 1.824
R20419 net5.n110 net5.n109 1.824
R20420 net5.n214 net5.n213 1.824
R20421 net5.n172 net5.n171 1.824
R20422 net5 net5.n6 1.696
R20423 net5.n31 net5.n29 1.57
R20424 net5.n72 net5.n70 1.57
R20425 net5.n11 net5.n9 1.57
R20426 net5.n94 net5.n92 1.57
R20427 net5.n198 net5.n196 1.57
R20428 net5.n177 net5.n175 1.57
R20429 net5.n156 net5.n154 1.57
R20430 net5.n135 net5.n133 1.57
R20431 net5.n115 net5.n113 1.57
R20432 net5.n51 net5.n49 1.57
R20433 net5 net5.n215 1.05
R20434 net5.n6 net5.n4 0.82
R20435 net5.n35 net5.n34 0.752
R20436 net5.n76 net5.n75 0.752
R20437 net5.n15 net5.n14 0.752
R20438 net5.n98 net5.n97 0.752
R20439 net5.n202 net5.n201 0.752
R20440 net5.n181 net5.n180 0.752
R20441 net5.n160 net5.n159 0.752
R20442 net5.n139 net5.n138 0.752
R20443 net5.n119 net5.n118 0.752
R20444 net5.n55 net5.n54 0.752
R20445 net5.n193 net5.n172 0.434
R20446 net5.n89 net5.n88 0.434
R20447 net5.n215 net5.n110 0.225
R20448 net5.n172 net5.n151 0.217
R20449 net5.n214 net5.n193 0.217
R20450 net5.n110 net5.n89 0.217
R20451 net5.n88 net5.n67 0.217
R20452 net5.n215 net5.n214 0.208
R20453 net5.n42 net5.n40 0.144
R20454 net5.n83 net5.n81 0.144
R20455 net5.n22 net5.n20 0.144
R20456 net5.n105 net5.n103 0.144
R20457 net5.n209 net5.n207 0.144
R20458 net5.n188 net5.n186 0.144
R20459 net5.n167 net5.n165 0.144
R20460 net5.n146 net5.n144 0.144
R20461 net5.n126 net5.n124 0.144
R20462 net5.n62 net5.n60 0.144
R20463 net5.n4 net5.n3 0.113
R20464 net5.n4 net5.n1 0.111
R20465 net5.n40 net5.n33 0.04
R20466 net5.n81 net5.n74 0.04
R20467 net5.n20 net5.n13 0.04
R20468 net5.n103 net5.n96 0.04
R20469 net5.n207 net5.n200 0.04
R20470 net5.n186 net5.n179 0.04
R20471 net5.n165 net5.n158 0.04
R20472 net5.n144 net5.n137 0.04
R20473 net5.n124 net5.n117 0.04
R20474 net5.n60 net5.n53 0.04
R20475 net5.n46 net5.n44 0.035
R20476 net5.n87 net5.n85 0.035
R20477 net5.n26 net5.n24 0.035
R20478 net5.n109 net5.n107 0.035
R20479 net5.n213 net5.n211 0.035
R20480 net5.n192 net5.n190 0.035
R20481 net5.n171 net5.n169 0.035
R20482 net5.n150 net5.n148 0.035
R20483 net5.n130 net5.n128 0.035
R20484 net5.n66 net5.n64 0.035
R20485 net5.n1 net5.n0 0.017
R20486 net5.n3 net5.n2 0.014
R20487 net5.n44 net5.n42 0.01
R20488 net5.n85 net5.n83 0.01
R20489 net5.n24 net5.n22 0.01
R20490 net5.n107 net5.n105 0.01
R20491 net5.n211 net5.n209 0.01
R20492 net5.n190 net5.n188 0.01
R20493 net5.n169 net5.n167 0.01
R20494 net5.n148 net5.n146 0.01
R20495 net5.n128 net5.n126 0.01
R20496 net5.n64 net5.n62 0.01
R20497 net5.n33 net5.n31 0.005
R20498 net5.n74 net5.n72 0.005
R20499 net5.n13 net5.n11 0.005
R20500 net5.n96 net5.n94 0.005
R20501 net5.n200 net5.n198 0.005
R20502 net5.n179 net5.n177 0.005
R20503 net5.n158 net5.n156 0.005
R20504 net5.n137 net5.n135 0.005
R20505 net5.n117 net5.n115 0.005
R20506 net5.n53 net5.n51 0.005
R20507 net5.n6 net5.n5 0.002
R20508 GND.n587 GND.n586 21413.3
R20509 GND.n2579 GND.n2577 20223.5
R20510 GND.n2661 GND.n2660 18154.5
R20511 GND.n2408 GND.n2406 16072.6
R20512 GND.n2490 GND.n2489 14260.7
R20513 GND.n2 GND.n603 8883.81
R20514 GND.n603 GND.n602 8883.81
R20515 GND.n602 GND.n601 8883.81
R20516 GND.n601 GND.n600 8883.81
R20517 GND.n600 GND.n599 8883.81
R20518 GND.n599 GND.n598 8883.81
R20519 GND.n598 GND.n597 8883.81
R20520 GND.n597 GND.n596 8883.81
R20521 GND.n596 GND.n595 8883.81
R20522 GND.n595 GND.n594 8883.81
R20523 GND.n594 GND.n593 8883.81
R20524 GND.n585 GND.n584 8883.81
R20525 GND.n586 GND.n585 8883.81
R20526 GND.n1 GND.n254 8800
R20527 GND.n254 GND.n253 8800
R20528 GND.n253 GND.n252 8800
R20529 GND.n252 GND.n251 8800
R20530 GND.n251 GND.n250 8800
R20531 GND.n250 GND.n249 8800
R20532 GND.n249 GND.n248 8800
R20533 GND.n447 GND.n446 8800
R20534 GND.n448 GND.n447 8800
R20535 GND.n449 GND.n448 8800
R20536 GND.n450 GND.n449 8800
R20537 GND.n2489 GND.t27 6555.56
R20538 GND.n2660 GND.t22 6555.56
R20539 GND.n3009 GND.t19 -6114.59
R20540 GND.n3035 GND.t1 -5965.62
R20541 GND.n2 GND.t43 5500
R20542 GND.n603 GND.t2 5500
R20543 GND.n602 GND.t47 5500
R20544 GND.n601 GND.t45 5500
R20545 GND.n600 GND.t4 5500
R20546 GND.n599 GND.t14 5500
R20547 GND.n598 GND.t8 5500
R20548 GND.n597 GND.t41 5500
R20549 GND.n596 GND.t12 5500
R20550 GND.n595 GND.t10 5500
R20551 GND.n594 GND.t51 5500
R20552 GND.n593 GND.t53 5500
R20553 GND.n584 GND.t16 5500
R20554 GND.n585 GND.t55 5500
R20555 GND.n586 GND.t6 5500
R20556 GND.n1 GND.t35 5484.72
R20557 GND.n254 GND.t37 5484.72
R20558 GND.n253 GND.t34 5484.72
R20559 GND.n252 GND.t36 5484.72
R20560 GND.n251 GND.t32 5484.72
R20561 GND.n250 GND.t33 5484.72
R20562 GND.n249 GND.t29 5484.72
R20563 GND.n248 GND.t31 5484.72
R20564 GND.n446 GND.t25 5484.72
R20565 GND.n447 GND.t30 5484.72
R20566 GND.n448 GND.t24 5484.72
R20567 GND.n449 GND.t26 5484.72
R20568 GND.n450 GND.t23 5484.72
R20569 GND.t19 GND.n3008 -7929.71
R20570 GND.t1 GND.n3034 -7790.44
R20571 GND.t39 GND.n2515 2179.44
R20572 GND.n2511 GND.n2510 2179.44
R20573 GND.n2510 GND.n2509 2179.44
R20574 GND.n2505 GND.n2504 2179.44
R20575 GND.n451 GND.n450 1417.83
R20576 GND.n0 GND.t39 1211.98
R20577 GND.n2278 GND.t18 1113.92
R20578 GND.t18 GND.t38 742.616
R20579 GND.n3030 GND.n3029 664.15
R20580 GND.n3034 GND.n3033 664.15
R20581 GND.n3004 GND.n3003 657.943
R20582 GND.n3008 GND.n3007 657.943
R20583 GND.n2514 GND.n2511 616.822
R20584 GND.n2509 GND.n2506 616.822
R20585 GND.n591 GND.n590 585
R20586 GND.n626 GND.n625 585
R20587 GND.n640 GND.n639 585
R20588 GND.n654 GND.n653 585
R20589 GND.n668 GND.n667 585
R20590 GND.n678 GND.n677 585
R20591 GND.n692 GND.n691 585
R20592 GND.n706 GND.n705 585
R20593 GND.n720 GND.n719 585
R20594 GND.n734 GND.n733 585
R20595 GND.n581 GND.n580 585
R20596 GND.n612 GND.n611 585
R20597 GND.n443 GND.n442 585
R20598 GND.n543 GND.n542 585
R20599 GND.n561 GND.n560 585
R20600 GND.n505 GND.n504 585
R20601 GND.n486 GND.n485 585
R20602 GND.n461 GND.n460 585
R20603 GND.n272 GND.n271 585
R20604 GND.n294 GND.n293 585
R20605 GND.n260 GND.n259 585
R20606 GND.n320 GND.n319 585
R20607 GND.n246 GND.n245 585
R20608 GND.n525 GND.n524 585
R20609 GND.n3033 GND.n3032 585
R20610 GND.n3031 GND.n3030 585
R20611 GND.n3007 GND.n3006 585
R20612 GND.n3005 GND.n3004 585
R20613 GND.n2539 GND.n2538 585
R20614 GND.n2525 GND.n2524 585
R20615 GND.n2499 GND.n2498 585
R20616 GND.n2553 GND.n2552 585
R20617 GND.n2514 GND.n2513 585
R20618 GND.n2509 GND.n2508 585
R20619 GND.n2504 GND.n2503 585
R20620 GND.n2575 GND.n2574 585
R20621 GND.n2657 GND.n2656 585
R20622 GND.n2596 GND.n2595 585
R20623 GND.n2639 GND.n2638 585
R20624 GND.n2486 GND.n2485 585
R20625 GND.n2468 GND.n2467 585
R20626 GND.n2422 GND.n2421 585
R20627 GND.n2404 GND.n2403 585
R20628 GND.n2504 GND.n2501 534.579
R20629 GND.n2 GND.n604 460.952
R20630 GND.n587 GND.n583 460.952
R20631 GND.n1 GND.n255 460.952
R20632 GND.n451 GND.n445 460.952
R20633 GND.n615 GND.n614 377.142
R20634 GND.n737 GND.n736 377.142
R20635 GND.n323 GND.n322 377.142
R20636 GND.n564 GND.n563 377.142
R20637 GND.n629 GND.n628 293.333
R20638 GND.n723 GND.n722 293.333
R20639 GND.n263 GND.n262 293.333
R20640 GND.n546 GND.n545 293.333
R20641 GND.n3073 GND.n3072 226.441
R20642 GND.n3080 GND.n3079 226.441
R20643 GND.n3118 GND.n3117 226.441
R20644 GND.n3111 GND.n3110 226.441
R20645 GND.n643 GND.n642 209.523
R20646 GND.n709 GND.n708 209.523
R20647 GND.n297 GND.n296 209.523
R20648 GND.n528 GND.n527 209.523
R20649 GND.n3072 GND.t20 205.247
R20650 GND.n3117 GND.t57 205.247
R20651 GND.n2408 GND.n2407 162.962
R20652 GND.n2490 GND.n2488 162.962
R20653 GND.n2579 GND.n2578 162.962
R20654 GND.n2661 GND.n2659 162.962
R20655 GND.n0 GND.n2516 162.962
R20656 GND.n2556 GND.n2555 162.962
R20657 GND.n3032 GND.n3031 131.333
R20658 GND.n3006 GND.n3005 128.945
R20659 GND.n657 GND.n656 125.714
R20660 GND.n695 GND.n694 125.714
R20661 GND.n275 GND.n274 125.714
R20662 GND.n508 GND.n507 125.714
R20663 GND.n146 GND.n145 92.5
R20664 GND.n197 GND.n196 92.5
R20665 GND.n778 GND.n777 92.5
R20666 GND.n829 GND.n828 92.5
R20667 GND.n30 GND.n29 92.5
R20668 GND.n81 GND.n80 92.5
R20669 GND.n896 GND.n895 92.5
R20670 GND.n947 GND.n946 92.5
R20671 GND.n2182 GND.n2181 92.5
R20672 GND.n2233 GND.n2232 92.5
R20673 GND.n2065 GND.n2064 92.5
R20674 GND.n2116 GND.n2115 92.5
R20675 GND.n1948 GND.n1947 92.5
R20676 GND.n1999 GND.n1998 92.5
R20677 GND.n1831 GND.n1830 92.5
R20678 GND.n1882 GND.n1881 92.5
R20679 GND.n1714 GND.n1713 92.5
R20680 GND.n1765 GND.n1764 92.5
R20681 GND.n1597 GND.n1596 92.5
R20682 GND.n1648 GND.n1647 92.5
R20683 GND.n1480 GND.n1479 92.5
R20684 GND.n1531 GND.n1530 92.5
R20685 GND.n1363 GND.n1362 92.5
R20686 GND.n1414 GND.n1413 92.5
R20687 GND.n1246 GND.n1245 92.5
R20688 GND.n1297 GND.n1296 92.5
R20689 GND.n1129 GND.n1128 92.5
R20690 GND.n1180 GND.n1179 92.5
R20691 GND.n1013 GND.n1012 92.5
R20692 GND.n1064 GND.n1063 92.5
R20693 GND.n2515 GND.n2514 82.242
R20694 GND.n2506 GND.n2505 82.242
R20695 GND.n2425 GND.n2424 81.481
R20696 GND.n2471 GND.n2470 81.481
R20697 GND.n2599 GND.n2598 81.481
R20698 GND.n2642 GND.n2641 81.481
R20699 GND.n2528 GND.n2527 81.481
R20700 GND.n2542 GND.n2541 81.481
R20701 GND.n145 GND.t7 70.344
R20702 GND.n777 GND.t56 70.344
R20703 GND.n29 GND.t17 70.344
R20704 GND.n895 GND.t54 70.344
R20705 GND.n2181 GND.t52 70.344
R20706 GND.n2064 GND.t11 70.344
R20707 GND.n1947 GND.t13 70.344
R20708 GND.n1830 GND.t42 70.344
R20709 GND.n1713 GND.t9 70.344
R20710 GND.n1596 GND.t15 70.344
R20711 GND.n1479 GND.t5 70.344
R20712 GND.n1362 GND.t46 70.344
R20713 GND.n1245 GND.t48 70.344
R20714 GND.n1128 GND.t3 70.344
R20715 GND.n1012 GND.t44 70.344
R20716 GND.n669 GND.n668 59.471
R20717 GND.n679 GND.n678 59.471
R20718 GND.n462 GND.n461 59.471
R20719 GND.n487 GND.n486 59.471
R20720 GND.n3071 GND.n3070 58.37
R20721 GND.n3078 GND.n3077 58.37
R20722 GND.n3116 GND.n3115 58.37
R20723 GND.n3109 GND.n3108 58.37
R20724 GND.n2513 GND.n2512 53.727
R20725 GND.n2508 GND.n2507 53.727
R20726 GND.n2526 GND.n2525 52.767
R20727 GND.n2540 GND.n2539 52.767
R20728 GND.n2597 GND.n2596 52.767
R20729 GND.n2640 GND.n2639 52.767
R20730 GND.n2423 GND.n2422 52.767
R20731 GND.n2469 GND.n2468 52.767
R20732 GND.n655 GND.n654 52.037
R20733 GND.n693 GND.n692 52.037
R20734 GND.n273 GND.n272 52.037
R20735 GND.n506 GND.n505 52.037
R20736 GND.n2503 GND.n2502 46.563
R20737 GND.n2500 GND.n2499 45.732
R20738 GND.n2554 GND.n2553 45.732
R20739 GND.n2576 GND.n2575 45.732
R20740 GND.n2658 GND.n2657 45.732
R20741 GND.n2405 GND.n2404 45.732
R20742 GND.n2487 GND.n2486 45.732
R20743 GND.n641 GND.n640 44.603
R20744 GND.n707 GND.n706 44.603
R20745 GND.n295 GND.n294 44.603
R20746 GND.n526 GND.n525 44.603
R20747 GND.n671 GND.n670 41.904
R20748 GND.n681 GND.n680 41.904
R20749 GND.n464 GND.n463 41.904
R20750 GND.n489 GND.n488 41.904
R20751 GND.n2 GND.n592 40.886
R20752 GND.n588 GND.n582 40.886
R20753 GND.n1 GND.n247 40.886
R20754 GND.n452 GND.n444 40.886
R20755 GND.n2320 GND.n2319 38.803
R20756 GND.n2357 GND.n2356 38.803
R20757 GND.n627 GND.n626 37.169
R20758 GND.n721 GND.n720 37.169
R20759 GND.n261 GND.n260 37.169
R20760 GND.n544 GND.n543 37.169
R20761 GND.n616 GND.n613 33.452
R20762 GND.n738 GND.n735 33.452
R20763 GND.n324 GND.n321 33.452
R20764 GND.n565 GND.n562 33.452
R20765 GND.n136 GND.n135 31.034
R20766 GND.n214 GND.n213 31.034
R20767 GND.n768 GND.n767 31.034
R20768 GND.n846 GND.n845 31.034
R20769 GND.n20 GND.n19 31.034
R20770 GND.n98 GND.n97 31.034
R20771 GND.n886 GND.n885 31.034
R20772 GND.n964 GND.n963 31.034
R20773 GND.n2172 GND.n2171 31.034
R20774 GND.n2250 GND.n2249 31.034
R20775 GND.n2055 GND.n2054 31.034
R20776 GND.n2133 GND.n2132 31.034
R20777 GND.n1938 GND.n1937 31.034
R20778 GND.n2016 GND.n2015 31.034
R20779 GND.n1821 GND.n1820 31.034
R20780 GND.n1899 GND.n1898 31.034
R20781 GND.n1704 GND.n1703 31.034
R20782 GND.n1782 GND.n1781 31.034
R20783 GND.n1587 GND.n1586 31.034
R20784 GND.n1665 GND.n1664 31.034
R20785 GND.n1470 GND.n1469 31.034
R20786 GND.n1548 GND.n1547 31.034
R20787 GND.n1353 GND.n1352 31.034
R20788 GND.n1431 GND.n1430 31.034
R20789 GND.n1236 GND.n1235 31.034
R20790 GND.n1314 GND.n1313 31.034
R20791 GND.n1119 GND.n1118 31.034
R20792 GND.n1197 GND.n1196 31.034
R20793 GND.n1003 GND.n1002 31.034
R20794 GND.n1081 GND.n1080 31.034
R20795 GND.n2279 GND.n2277 29.848
R20796 GND.n613 GND.n612 29.735
R20797 GND.n735 GND.n734 29.735
R20798 GND.n321 GND.n320 29.735
R20799 GND.n562 GND.n561 29.735
R20800 GND.n2285 GND.n2284 27.976
R20801 GND.n3052 GND.n3051 27.617
R20802 GND.n2998 GND.t28 27.523
R20803 GND.n3026 GND.n3025 27.215
R20804 GND.n2295 GND.n2294 26.863
R20805 GND.n2382 GND.n2381 26.863
R20806 GND.n630 GND.n627 26.018
R20807 GND.n724 GND.n721 26.018
R20808 GND.n264 GND.n261 26.018
R20809 GND.n547 GND.n544 26.018
R20810 GND.n3057 GND.t21 23.416
R20811 GND.n3093 GND.t58 23.416
R20812 GND.n2383 GND.n2382 22.597
R20813 GND.n2296 GND.n2295 22.597
R20814 GND.n592 GND.n591 22.301
R20815 GND.n582 GND.n581 22.301
R20816 GND.n247 GND.n246 22.301
R20817 GND.n444 GND.n443 22.301
R20818 GND.n2333 GND.n2332 21.561
R20819 GND.n2344 GND.n2343 21.561
R20820 GND.n2345 GND.n2344 21.561
R20821 GND.n2332 GND.n2331 21.561
R20822 GND.n2392 GND.t49 21.289
R20823 GND.n2392 GND.t40 21.191
R20824 GND.n2284 GND.n2283 20.893
R20825 GND.n2696 GND.n2695 20.382
R20826 GND.n2560 GND.n2559 20.068
R20827 GND.n644 GND.n641 18.584
R20828 GND.n710 GND.n707 18.584
R20829 GND.n298 GND.n295 18.584
R20830 GND.n529 GND.n526 18.584
R20831 GND.n2310 GND.n2308 17.909
R20832 GND.n2372 GND.n2370 17.909
R20833 GND.n2308 GND.n2307 15.969
R20834 GND.n2369 GND.n2368 15.969
R20835 GND.n2370 GND.n2369 15.969
R20836 GND.n2307 GND.n2306 15.969
R20837 GND.n0 GND.n2500 14.071
R20838 GND.n2557 GND.n2554 14.071
R20839 GND.n2580 GND.n2576 14.071
R20840 GND.n2662 GND.n2658 14.071
R20841 GND.n2409 GND.n2405 14.071
R20842 GND.n2491 GND.n2487 14.071
R20843 GND.n2952 GND.t50 13.384
R20844 GND.n2358 GND.n2357 11.521
R20845 GND.n2321 GND.n2320 11.521
R20846 GND.n658 GND.n655 11.15
R20847 GND.n696 GND.n693 11.15
R20848 GND.n276 GND.n273 11.15
R20849 GND.n509 GND.n506 11.15
R20850 GND.n2276 GND.n2275 10.264
R20851 GND.n2277 GND.n2276 10.264
R20852 GND.n3053 GND.n2391 10.213
R20853 GND.n3074 GND.n3073 9.433
R20854 GND.n3081 GND.n3080 9.433
R20855 GND.n3119 GND.n3118 9.433
R20856 GND.n3112 GND.n3111 9.433
R20857 GND.n157 GND.n156 9.3
R20858 GND.n137 GND.n136 9.3
R20859 GND.n215 GND.n214 9.3
R20860 GND.n223 GND.n222 9.3
R20861 GND.n789 GND.n788 9.3
R20862 GND.n769 GND.n768 9.3
R20863 GND.n847 GND.n846 9.3
R20864 GND.n855 GND.n854 9.3
R20865 GND.n41 GND.n40 9.3
R20866 GND.n21 GND.n20 9.3
R20867 GND.n99 GND.n98 9.3
R20868 GND.n107 GND.n106 9.3
R20869 GND.n907 GND.n906 9.3
R20870 GND.n887 GND.n886 9.3
R20871 GND.n965 GND.n964 9.3
R20872 GND.n973 GND.n972 9.3
R20873 GND.n2193 GND.n2192 9.3
R20874 GND.n2173 GND.n2172 9.3
R20875 GND.n2251 GND.n2250 9.3
R20876 GND.n2259 GND.n2258 9.3
R20877 GND.n2076 GND.n2075 9.3
R20878 GND.n2056 GND.n2055 9.3
R20879 GND.n2134 GND.n2133 9.3
R20880 GND.n2142 GND.n2141 9.3
R20881 GND.n1959 GND.n1958 9.3
R20882 GND.n1939 GND.n1938 9.3
R20883 GND.n2017 GND.n2016 9.3
R20884 GND.n2025 GND.n2024 9.3
R20885 GND.n1842 GND.n1841 9.3
R20886 GND.n1822 GND.n1821 9.3
R20887 GND.n1900 GND.n1899 9.3
R20888 GND.n1908 GND.n1907 9.3
R20889 GND.n1725 GND.n1724 9.3
R20890 GND.n1705 GND.n1704 9.3
R20891 GND.n1783 GND.n1782 9.3
R20892 GND.n1791 GND.n1790 9.3
R20893 GND.n1608 GND.n1607 9.3
R20894 GND.n1588 GND.n1587 9.3
R20895 GND.n1666 GND.n1665 9.3
R20896 GND.n1674 GND.n1673 9.3
R20897 GND.n1491 GND.n1490 9.3
R20898 GND.n1471 GND.n1470 9.3
R20899 GND.n1549 GND.n1548 9.3
R20900 GND.n1557 GND.n1556 9.3
R20901 GND.n1374 GND.n1373 9.3
R20902 GND.n1354 GND.n1353 9.3
R20903 GND.n1432 GND.n1431 9.3
R20904 GND.n1440 GND.n1439 9.3
R20905 GND.n1257 GND.n1256 9.3
R20906 GND.n1237 GND.n1236 9.3
R20907 GND.n1315 GND.n1314 9.3
R20908 GND.n1323 GND.n1322 9.3
R20909 GND.n1140 GND.n1139 9.3
R20910 GND.n1120 GND.n1119 9.3
R20911 GND.n1198 GND.n1197 9.3
R20912 GND.n1206 GND.n1205 9.3
R20913 GND.n1024 GND.n1023 9.3
R20914 GND.n1004 GND.n1003 9.3
R20915 GND.n1082 GND.n1081 9.3
R20916 GND.n1090 GND.n1089 9.3
R20917 GND.n742 GND.n741 9.3
R20918 GND.n728 GND.n727 9.3
R20919 GND.n714 GND.n713 9.3
R20920 GND.n700 GND.n699 9.3
R20921 GND.n686 GND.n685 9.3
R20922 GND.n664 GND.n663 9.3
R20923 GND.n650 GND.n649 9.3
R20924 GND.n636 GND.n635 9.3
R20925 GND.n622 GND.n621 9.3
R20926 GND.n608 GND.n607 9.3
R20927 GND.n618 GND.n617 9.3
R20928 GND.n617 GND.n616 9.3
R20929 GND.n616 GND.n615 9.3
R20930 GND.n620 GND.n619 9.3
R20931 GND.n632 GND.n631 9.3
R20932 GND.n631 GND.n630 9.3
R20933 GND.n630 GND.n629 9.3
R20934 GND.n634 GND.n633 9.3
R20935 GND.n646 GND.n645 9.3
R20936 GND.n645 GND.n644 9.3
R20937 GND.n644 GND.n643 9.3
R20938 GND.n648 GND.n647 9.3
R20939 GND.n660 GND.n659 9.3
R20940 GND.n659 GND.n658 9.3
R20941 GND.n658 GND.n657 9.3
R20942 GND.n662 GND.n661 9.3
R20943 GND.n674 GND.n673 9.3
R20944 GND.n673 GND.n672 9.3
R20945 GND.n672 GND.n671 9.3
R20946 GND.n688 GND.n687 9.3
R20947 GND.n684 GND.n683 9.3
R20948 GND.n683 GND.n682 9.3
R20949 GND.n682 GND.n681 9.3
R20950 GND.n702 GND.n701 9.3
R20951 GND.n698 GND.n697 9.3
R20952 GND.n697 GND.n696 9.3
R20953 GND.n696 GND.n695 9.3
R20954 GND.n716 GND.n715 9.3
R20955 GND.n712 GND.n711 9.3
R20956 GND.n711 GND.n710 9.3
R20957 GND.n710 GND.n709 9.3
R20958 GND.n730 GND.n729 9.3
R20959 GND.n726 GND.n725 9.3
R20960 GND.n725 GND.n724 9.3
R20961 GND.n724 GND.n723 9.3
R20962 GND.n744 GND.n743 9.3
R20963 GND.n740 GND.n739 9.3
R20964 GND.n739 GND.n738 9.3
R20965 GND.n738 GND.n737 9.3
R20966 GND.n589 GND.n588 9.3
R20967 GND.n588 GND.n587 9.3
R20968 GND.n606 GND.n605 9.3
R20969 GND.n530 GND.n529 9.3
R20970 GND.n529 GND.n528 9.3
R20971 GND.n548 GND.n547 9.3
R20972 GND.n547 GND.n546 9.3
R20973 GND.n566 GND.n565 9.3
R20974 GND.n565 GND.n564 9.3
R20975 GND.n453 GND.n452 9.3
R20976 GND.n452 GND.n451 9.3
R20977 GND.n325 GND.n324 9.3
R20978 GND.n324 GND.n323 9.3
R20979 GND.n265 GND.n264 9.3
R20980 GND.n264 GND.n263 9.3
R20981 GND.n299 GND.n298 9.3
R20982 GND.n298 GND.n297 9.3
R20983 GND.n277 GND.n276 9.3
R20984 GND.n276 GND.n275 9.3
R20985 GND.n466 GND.n465 9.3
R20986 GND.n465 GND.n464 9.3
R20987 GND.n491 GND.n490 9.3
R20988 GND.n490 GND.n489 9.3
R20989 GND.n510 GND.n509 9.3
R20990 GND.n509 GND.n508 9.3
R20991 GND.n2759 GND.n2758 9.3
R20992 GND.n2861 GND.n2860 9.3
R20993 GND.n2388 GND.n2387 9.3
R20994 GND.n2376 GND.n2375 9.3
R20995 GND.n2363 GND.n2362 9.3
R20996 GND.n2351 GND.n2350 9.3
R20997 GND.n2328 GND.n2327 9.3
R20998 GND.n2316 GND.n2315 9.3
R20999 GND.n2303 GND.n2302 9.3
R21000 GND.n2291 GND.n2290 9.3
R21001 GND.n2390 GND.n2389 9.3
R21002 GND.n2378 GND.n2377 9.3
R21003 GND.n2365 GND.n2364 9.3
R21004 GND.n2353 GND.n2352 9.3
R21005 GND.n2289 GND.n2288 9.3
R21006 GND.n2299 GND.n2298 9.3
R21007 GND.n2298 GND.n2297 9.3
R21008 GND.n2301 GND.n2300 9.3
R21009 GND.n2312 GND.n2311 9.3
R21010 GND.n2311 GND.n2310 9.3
R21011 GND.n2314 GND.n2313 9.3
R21012 GND.n2324 GND.n2323 9.3
R21013 GND.n2323 GND.n2322 9.3
R21014 GND.n2326 GND.n2325 9.3
R21015 GND.n2337 GND.n2336 9.3
R21016 GND.n2336 GND.n2335 9.3
R21017 GND.n2349 GND.n2348 9.3
R21018 GND.n2348 GND.n2347 9.3
R21019 GND.n2361 GND.n2360 9.3
R21020 GND.n2360 GND.n2359 9.3
R21021 GND.n2374 GND.n2373 9.3
R21022 GND.n2373 GND.n2372 9.3
R21023 GND.n2386 GND.n2385 9.3
R21024 GND.n2385 GND.n2384 9.3
R21025 GND.n2280 GND.n2279 9.3
R21026 GND.n2279 GND.n2278 9.3
R21027 GND.n2287 GND.n2286 9.3
R21028 GND.n3036 GND.n3035 9.3
R21029 GND.n3043 GND.n3042 9.3
R21030 GND.n3010 GND.n3009 9.3
R21031 GND.n3022 GND.n3021 9.3
R21032 GND.n2692 GND.n2691 9.3
R21033 GND.n2677 GND.n2676 9.3
R21034 GND.n2672 GND.n2671 9.3
R21035 GND.n2675 GND.n2674 9.3
R21036 GND.n2682 GND.n2681 9.3
R21037 GND.n2681 GND.n2680 9.3
R21038 GND.n2694 GND.n2693 9.3
R21039 GND.n2690 GND.n2689 9.3
R21040 GND.n2689 GND.n2688 9.3
R21041 GND.n2565 GND.n2564 9.3
R21042 GND.n2564 GND.n2563 9.3
R21043 GND.n2644 GND.n2643 9.3
R21044 GND.n2643 GND.n2642 9.3
R21045 GND.n2601 GND.n2600 9.3
R21046 GND.n2600 GND.n2599 9.3
R21047 GND.n2663 GND.n2662 9.3
R21048 GND.n2662 GND.n2661 9.3
R21049 GND.n2581 GND.n2580 9.3
R21050 GND.n2580 GND.n2579 9.3
R21051 GND.n2410 GND.n2409 9.3
R21052 GND.n2409 GND.n2408 9.3
R21053 GND.n2427 GND.n2426 9.3
R21054 GND.n2426 GND.n2425 9.3
R21055 GND.n2473 GND.n2472 9.3
R21056 GND.n2472 GND.n2471 9.3
R21057 GND.n2492 GND.n2491 9.3
R21058 GND.n2491 GND.n2490 9.3
R21059 GND.n2521 GND.n2520 9.3
R21060 GND.n2547 GND.n2546 9.3
R21061 GND.n2558 GND.n2557 9.3
R21062 GND.n2557 GND.n2556 9.3
R21063 GND.n2549 GND.n2548 9.3
R21064 GND.n2519 GND.n2518 9.3
R21065 GND.n2531 GND.n2530 9.3
R21066 GND.n2530 GND.n2529 9.3
R21067 GND.n2529 GND.n2528 9.3
R21068 GND.n2545 GND.n2544 9.3
R21069 GND.n2544 GND.n2543 9.3
R21070 GND.n2543 GND.n2542 9.3
R21071 GND.n2825 GND.n2824 9.154
R21072 GND.n2339 GND.n2338 9.154
R21073 GND.n2684 GND.n2683 9.154
R21074 GND.n2618 GND.n2617 9.154
R21075 GND.n2617 GND.n2616 9.154
R21076 GND.n2447 GND.n2446 9.154
R21077 GND.n2446 GND.n2445 9.154
R21078 GND.n2534 GND.n2533 9.154
R21079 GND.n2533 GND.n2532 9.154
R21080 GND.n2953 GND.n2952 8.855
R21081 GND.n147 GND.n146 8.282
R21082 GND.n198 GND.n197 8.282
R21083 GND.n779 GND.n778 8.282
R21084 GND.n830 GND.n829 8.282
R21085 GND.n31 GND.n30 8.282
R21086 GND.n82 GND.n81 8.282
R21087 GND.n897 GND.n896 8.282
R21088 GND.n948 GND.n947 8.282
R21089 GND.n2183 GND.n2182 8.282
R21090 GND.n2234 GND.n2233 8.282
R21091 GND.n2066 GND.n2065 8.282
R21092 GND.n2117 GND.n2116 8.282
R21093 GND.n1949 GND.n1948 8.282
R21094 GND.n2000 GND.n1999 8.282
R21095 GND.n1832 GND.n1831 8.282
R21096 GND.n1883 GND.n1882 8.282
R21097 GND.n1715 GND.n1714 8.282
R21098 GND.n1766 GND.n1765 8.282
R21099 GND.n1598 GND.n1597 8.282
R21100 GND.n1649 GND.n1648 8.282
R21101 GND.n1481 GND.n1480 8.282
R21102 GND.n1532 GND.n1531 8.282
R21103 GND.n1364 GND.n1363 8.282
R21104 GND.n1415 GND.n1414 8.282
R21105 GND.n1247 GND.n1246 8.282
R21106 GND.n1298 GND.n1297 8.282
R21107 GND.n1130 GND.n1129 8.282
R21108 GND.n1181 GND.n1180 8.282
R21109 GND.n1014 GND.n1013 8.282
R21110 GND.n1065 GND.n1064 8.282
R21111 GND.n2824 GND.t0 7.141
R21112 GND.n2529 GND.n2526 7.035
R21113 GND.n2543 GND.n2540 7.035
R21114 GND.n2600 GND.n2597 7.035
R21115 GND.n2643 GND.n2640 7.035
R21116 GND.n2426 GND.n2423 7.035
R21117 GND.n2472 GND.n2469 7.035
R21118 GND.n2970 GND.n2969 7.03
R21119 GND.n2919 GND.n2918 7.029
R21120 GND.n2703 GND.n2702 7.029
R21121 GND.n2993 GND.n2992 6.681
R21122 GND.n577 GND.n576 6.436
R21123 GND.n2335 GND.n2333 5.969
R21124 GND.n2347 GND.n2345 5.969
R21125 GND.n137 GND.n133 5.647
R21126 GND.n215 GND.n211 5.647
R21127 GND.n769 GND.n765 5.647
R21128 GND.n847 GND.n843 5.647
R21129 GND.n21 GND.n17 5.647
R21130 GND.n99 GND.n95 5.647
R21131 GND.n887 GND.n883 5.647
R21132 GND.n965 GND.n961 5.647
R21133 GND.n2173 GND.n2169 5.647
R21134 GND.n2251 GND.n2247 5.647
R21135 GND.n2056 GND.n2052 5.647
R21136 GND.n2134 GND.n2130 5.647
R21137 GND.n1939 GND.n1935 5.647
R21138 GND.n2017 GND.n2013 5.647
R21139 GND.n1822 GND.n1818 5.647
R21140 GND.n1900 GND.n1896 5.647
R21141 GND.n1705 GND.n1701 5.647
R21142 GND.n1783 GND.n1779 5.647
R21143 GND.n1588 GND.n1584 5.647
R21144 GND.n1666 GND.n1662 5.647
R21145 GND.n1471 GND.n1467 5.647
R21146 GND.n1549 GND.n1545 5.647
R21147 GND.n1354 GND.n1350 5.647
R21148 GND.n1432 GND.n1428 5.647
R21149 GND.n1237 GND.n1233 5.647
R21150 GND.n1315 GND.n1311 5.647
R21151 GND.n1120 GND.n1116 5.647
R21152 GND.n1198 GND.n1194 5.647
R21153 GND.n1004 GND.n1000 5.647
R21154 GND.n1082 GND.n1078 5.647
R21155 GND.n3127 GND.n3090 5.223
R21156 GND.n2664 GND.n2663 5.122
R21157 GND.n2493 GND.n2492 5.122
R21158 GND.n2582 GND.n2581 4.903
R21159 GND.n2411 GND.n2410 4.903
R21160 GND.n195 GND.n194 4.65
R21161 GND.n827 GND.n826 4.65
R21162 GND.n79 GND.n78 4.65
R21163 GND.n945 GND.n944 4.65
R21164 GND.n2231 GND.n2230 4.65
R21165 GND.n2114 GND.n2113 4.65
R21166 GND.n1997 GND.n1996 4.65
R21167 GND.n1880 GND.n1879 4.65
R21168 GND.n1763 GND.n1762 4.65
R21169 GND.n1646 GND.n1645 4.65
R21170 GND.n1529 GND.n1528 4.65
R21171 GND.n1412 GND.n1411 4.65
R21172 GND.n1295 GND.n1294 4.65
R21173 GND.n1178 GND.n1177 4.65
R21174 GND.n1062 GND.n1061 4.65
R21175 GND.n2954 GND.n2953 4.65
R21176 GND.n2826 GND.n2825 4.65
R21177 GND.n2340 GND.n2339 4.65
R21178 GND.n2685 GND.n2684 4.65
R21179 GND.n2619 GND.n2618 4.65
R21180 GND.n2448 GND.n2447 4.65
R21181 GND.n2535 GND.n2534 4.65
R21182 GND.n229 GND.n227 4.5
R21183 GND.n217 GND.n216 4.5
R21184 GND.n206 GND.n205 4.5
R21185 GND.n199 GND.n198 4.5
R21186 GND.n151 GND.n139 4.5
R21187 GND.n148 GND.n147 4.5
R21188 GND.n193 GND.n192 4.5
R21189 GND.n162 GND.n161 4.5
R21190 GND.n861 GND.n859 4.5
R21191 GND.n849 GND.n848 4.5
R21192 GND.n838 GND.n837 4.5
R21193 GND.n831 GND.n830 4.5
R21194 GND.n783 GND.n771 4.5
R21195 GND.n780 GND.n779 4.5
R21196 GND.n825 GND.n824 4.5
R21197 GND.n794 GND.n793 4.5
R21198 GND.n113 GND.n111 4.5
R21199 GND.n101 GND.n100 4.5
R21200 GND.n90 GND.n89 4.5
R21201 GND.n83 GND.n82 4.5
R21202 GND.n35 GND.n23 4.5
R21203 GND.n32 GND.n31 4.5
R21204 GND.n77 GND.n76 4.5
R21205 GND.n46 GND.n45 4.5
R21206 GND.n979 GND.n977 4.5
R21207 GND.n967 GND.n966 4.5
R21208 GND.n956 GND.n955 4.5
R21209 GND.n949 GND.n948 4.5
R21210 GND.n901 GND.n889 4.5
R21211 GND.n898 GND.n897 4.5
R21212 GND.n943 GND.n942 4.5
R21213 GND.n912 GND.n911 4.5
R21214 GND.n2265 GND.n2263 4.5
R21215 GND.n2253 GND.n2252 4.5
R21216 GND.n2242 GND.n2241 4.5
R21217 GND.n2235 GND.n2234 4.5
R21218 GND.n2187 GND.n2175 4.5
R21219 GND.n2184 GND.n2183 4.5
R21220 GND.n2229 GND.n2228 4.5
R21221 GND.n2198 GND.n2197 4.5
R21222 GND.n2148 GND.n2146 4.5
R21223 GND.n2136 GND.n2135 4.5
R21224 GND.n2125 GND.n2124 4.5
R21225 GND.n2118 GND.n2117 4.5
R21226 GND.n2070 GND.n2058 4.5
R21227 GND.n2067 GND.n2066 4.5
R21228 GND.n2112 GND.n2111 4.5
R21229 GND.n2081 GND.n2080 4.5
R21230 GND.n2031 GND.n2029 4.5
R21231 GND.n2019 GND.n2018 4.5
R21232 GND.n2008 GND.n2007 4.5
R21233 GND.n2001 GND.n2000 4.5
R21234 GND.n1953 GND.n1941 4.5
R21235 GND.n1950 GND.n1949 4.5
R21236 GND.n1995 GND.n1994 4.5
R21237 GND.n1964 GND.n1963 4.5
R21238 GND.n1914 GND.n1912 4.5
R21239 GND.n1902 GND.n1901 4.5
R21240 GND.n1891 GND.n1890 4.5
R21241 GND.n1884 GND.n1883 4.5
R21242 GND.n1836 GND.n1824 4.5
R21243 GND.n1833 GND.n1832 4.5
R21244 GND.n1878 GND.n1877 4.5
R21245 GND.n1847 GND.n1846 4.5
R21246 GND.n1797 GND.n1795 4.5
R21247 GND.n1785 GND.n1784 4.5
R21248 GND.n1774 GND.n1773 4.5
R21249 GND.n1767 GND.n1766 4.5
R21250 GND.n1719 GND.n1707 4.5
R21251 GND.n1716 GND.n1715 4.5
R21252 GND.n1761 GND.n1760 4.5
R21253 GND.n1730 GND.n1729 4.5
R21254 GND.n1680 GND.n1678 4.5
R21255 GND.n1668 GND.n1667 4.5
R21256 GND.n1657 GND.n1656 4.5
R21257 GND.n1650 GND.n1649 4.5
R21258 GND.n1602 GND.n1590 4.5
R21259 GND.n1599 GND.n1598 4.5
R21260 GND.n1644 GND.n1643 4.5
R21261 GND.n1613 GND.n1612 4.5
R21262 GND.n1563 GND.n1561 4.5
R21263 GND.n1551 GND.n1550 4.5
R21264 GND.n1540 GND.n1539 4.5
R21265 GND.n1533 GND.n1532 4.5
R21266 GND.n1485 GND.n1473 4.5
R21267 GND.n1482 GND.n1481 4.5
R21268 GND.n1527 GND.n1526 4.5
R21269 GND.n1496 GND.n1495 4.5
R21270 GND.n1446 GND.n1444 4.5
R21271 GND.n1434 GND.n1433 4.5
R21272 GND.n1423 GND.n1422 4.5
R21273 GND.n1416 GND.n1415 4.5
R21274 GND.n1368 GND.n1356 4.5
R21275 GND.n1365 GND.n1364 4.5
R21276 GND.n1410 GND.n1409 4.5
R21277 GND.n1379 GND.n1378 4.5
R21278 GND.n1329 GND.n1327 4.5
R21279 GND.n1317 GND.n1316 4.5
R21280 GND.n1306 GND.n1305 4.5
R21281 GND.n1299 GND.n1298 4.5
R21282 GND.n1251 GND.n1239 4.5
R21283 GND.n1248 GND.n1247 4.5
R21284 GND.n1293 GND.n1292 4.5
R21285 GND.n1262 GND.n1261 4.5
R21286 GND.n1212 GND.n1210 4.5
R21287 GND.n1200 GND.n1199 4.5
R21288 GND.n1189 GND.n1188 4.5
R21289 GND.n1182 GND.n1181 4.5
R21290 GND.n1134 GND.n1122 4.5
R21291 GND.n1131 GND.n1130 4.5
R21292 GND.n1176 GND.n1175 4.5
R21293 GND.n1145 GND.n1144 4.5
R21294 GND.n1096 GND.n1094 4.5
R21295 GND.n1084 GND.n1083 4.5
R21296 GND.n1073 GND.n1072 4.5
R21297 GND.n1066 GND.n1065 4.5
R21298 GND.n1018 GND.n1006 4.5
R21299 GND.n1015 GND.n1014 4.5
R21300 GND.n1060 GND.n1059 4.5
R21301 GND.n1029 GND.n1028 4.5
R21302 GND.n327 GND.n326 4.5
R21303 GND.n569 GND.n568 4.5
R21304 GND.n551 GND.n550 4.5
R21305 GND.n494 GND.n493 4.5
R21306 GND.n301 GND.n300 4.5
R21307 GND.n308 GND.n266 4.5
R21308 GND.n281 GND.n278 4.5
R21309 GND.n468 GND.n467 4.5
R21310 GND.n474 GND.n473 4.5
R21311 GND.n482 GND.n481 4.5
R21312 GND.n513 GND.n512 4.5
R21313 GND.n533 GND.n532 4.5
R21314 GND.n2964 GND.n2963 4.5
R21315 GND.n2987 GND.n2986 4.5
R21316 GND.n2951 GND.n2950 4.5
R21317 GND.n2956 GND.n2955 4.5
R21318 GND.n2725 GND.n2720 4.5
R21319 GND.n2864 GND.n2856 4.5
R21320 GND.n2888 GND.n2882 4.5
R21321 GND.n2843 GND.n2842 4.5
R21322 GND.n2813 GND.n2810 4.5
R21323 GND.n2828 GND.n2822 4.5
R21324 GND.n2802 GND.n2799 4.5
R21325 GND.n2818 GND.n2817 4.5
R21326 GND.n2792 GND.n2787 4.5
R21327 GND.n2770 GND.n2769 4.5
R21328 GND.n2744 GND.n2740 4.5
R21329 GND.n2907 GND.n2906 4.5
R21330 GND.n3039 GND.n3038 4.5
R21331 GND.n3046 GND.n3045 4.5
R21332 GND.n3013 GND.n3012 4.5
R21333 GND.n3023 GND.n3018 4.5
R21334 GND.n2614 GND.n2613 4.5
R21335 GND.n2632 GND.n2631 4.5
R21336 GND.n2621 GND.n2620 4.5
R21337 GND.n2647 GND.n2646 4.5
R21338 GND.n2609 GND.n2608 4.5
R21339 GND.n2603 GND.n2602 4.5
R21340 GND.n2450 GND.n2449 4.5
R21341 GND.n2443 GND.n2442 4.5
R21342 GND.n2461 GND.n2460 4.5
R21343 GND.n2436 GND.n2435 4.5
R21344 GND.n2430 GND.n2428 4.5
R21345 GND.n2476 GND.n2475 4.5
R21346 GND.n2999 GND.n2933 4.302
R21347 GND.n606 GND.n2 4.286
R21348 GND.n2673 GND.n2668 4.205
R21349 GND.n745 GND.n589 4.172
R21350 GND.n2882 GND.n2879 4.141
R21351 GND.n2740 GND.n2739 4.141
R21352 GND.n135 GND.n134 4.137
R21353 GND.n213 GND.n212 4.137
R21354 GND.n767 GND.n766 4.137
R21355 GND.n845 GND.n844 4.137
R21356 GND.n19 GND.n18 4.137
R21357 GND.n97 GND.n96 4.137
R21358 GND.n885 GND.n884 4.137
R21359 GND.n963 GND.n962 4.137
R21360 GND.n2171 GND.n2170 4.137
R21361 GND.n2249 GND.n2248 4.137
R21362 GND.n2054 GND.n2053 4.137
R21363 GND.n2132 GND.n2131 4.137
R21364 GND.n1937 GND.n1936 4.137
R21365 GND.n2015 GND.n2014 4.137
R21366 GND.n1820 GND.n1819 4.137
R21367 GND.n1898 GND.n1897 4.137
R21368 GND.n1703 GND.n1702 4.137
R21369 GND.n1781 GND.n1780 4.137
R21370 GND.n1586 GND.n1585 4.137
R21371 GND.n1664 GND.n1663 4.137
R21372 GND.n1469 GND.n1468 4.137
R21373 GND.n1547 GND.n1546 4.137
R21374 GND.n1352 GND.n1351 4.137
R21375 GND.n1430 GND.n1429 4.137
R21376 GND.n1235 GND.n1234 4.137
R21377 GND.n1313 GND.n1312 4.137
R21378 GND.n1118 GND.n1117 4.137
R21379 GND.n1196 GND.n1195 4.137
R21380 GND.n1002 GND.n1001 4.137
R21381 GND.n1080 GND.n1079 4.137
R21382 GND.n2517 GND.n2497 4.123
R21383 GND.n2289 GND.n2287 4.071
R21384 GND.n2998 GND.n2997 4.041
R21385 GND.n2391 GND.n2280 3.956
R21386 GND.n3046 GND.n3043 3.836
R21387 GND.n3023 GND.n3022 3.836
R21388 GND.n666 GND.n665 3.792
R21389 GND.n676 GND.n675 3.792
R21390 GND.n3069 GND.n3068 3.792
R21391 GND.n3076 GND.n3075 3.792
R21392 GND.n3114 GND.n3113 3.792
R21393 GND.n3107 GND.n3106 3.792
R21394 GND.n3013 GND.n3010 3.77
R21395 GND.n3039 GND.n3036 3.77
R21396 GND.n161 GND.n159 3.764
R21397 GND.n216 GND.n209 3.764
R21398 GND.n793 GND.n791 3.764
R21399 GND.n848 GND.n841 3.764
R21400 GND.n45 GND.n43 3.764
R21401 GND.n100 GND.n93 3.764
R21402 GND.n911 GND.n909 3.764
R21403 GND.n966 GND.n959 3.764
R21404 GND.n2197 GND.n2195 3.764
R21405 GND.n2252 GND.n2245 3.764
R21406 GND.n2080 GND.n2078 3.764
R21407 GND.n2135 GND.n2128 3.764
R21408 GND.n1963 GND.n1961 3.764
R21409 GND.n2018 GND.n2011 3.764
R21410 GND.n1846 GND.n1844 3.764
R21411 GND.n1901 GND.n1894 3.764
R21412 GND.n1729 GND.n1727 3.764
R21413 GND.n1784 GND.n1777 3.764
R21414 GND.n1612 GND.n1610 3.764
R21415 GND.n1667 GND.n1660 3.764
R21416 GND.n1495 GND.n1493 3.764
R21417 GND.n1550 GND.n1543 3.764
R21418 GND.n1378 GND.n1376 3.764
R21419 GND.n1433 GND.n1426 3.764
R21420 GND.n1261 GND.n1259 3.764
R21421 GND.n1316 GND.n1309 3.764
R21422 GND.n1144 GND.n1142 3.764
R21423 GND.n1199 GND.n1192 3.764
R21424 GND.n1028 GND.n1026 3.764
R21425 GND.n1083 GND.n1076 3.764
R21426 GND.n2856 GND.n2853 3.764
R21427 GND.n2787 GND.n2785 3.764
R21428 GND.n2517 GND.n0 3.734
R21429 GND.n2559 GND.n2558 3.734
R21430 GND.n2673 GND.n2672 3.734
R21431 GND.n2695 GND.n2565 3.734
R21432 GND.n672 GND.n669 3.716
R21433 GND.n682 GND.n679 3.716
R21434 GND.n465 GND.n462 3.716
R21435 GND.n490 GND.n487 3.716
R21436 GND.n3082 GND.n3074 3.702
R21437 GND.n3120 GND.n3119 3.702
R21438 GND.n3035 GND.n3028 3.648
R21439 GND.n3042 GND.n3041 3.648
R21440 GND.n3009 GND.n3002 3.581
R21441 GND.n3021 GND.n3020 3.581
R21442 GND.n2523 GND.n2522 3.555
R21443 GND.n2537 GND.n2536 3.555
R21444 GND.n2679 GND.n2678 3.555
R21445 GND.n2687 GND.n2686 3.555
R21446 GND.n3082 GND.n3081 3.517
R21447 GND.n3120 GND.n3112 3.517
R21448 GND.n3080 GND.n3078 3.495
R21449 GND.n3073 GND.n3071 3.495
R21450 GND.n3111 GND.n3109 3.495
R21451 GND.n3118 GND.n3116 3.495
R21452 GND.n139 GND.n138 3.388
R21453 GND.n227 GND.n226 3.388
R21454 GND.n771 GND.n770 3.388
R21455 GND.n859 GND.n858 3.388
R21456 GND.n23 GND.n22 3.388
R21457 GND.n111 GND.n110 3.388
R21458 GND.n889 GND.n888 3.388
R21459 GND.n977 GND.n976 3.388
R21460 GND.n2175 GND.n2174 3.388
R21461 GND.n2263 GND.n2262 3.388
R21462 GND.n2058 GND.n2057 3.388
R21463 GND.n2146 GND.n2145 3.388
R21464 GND.n1941 GND.n1940 3.388
R21465 GND.n2029 GND.n2028 3.388
R21466 GND.n1824 GND.n1823 3.388
R21467 GND.n1912 GND.n1911 3.388
R21468 GND.n1707 GND.n1706 3.388
R21469 GND.n1795 GND.n1794 3.388
R21470 GND.n1590 GND.n1589 3.388
R21471 GND.n1678 GND.n1677 3.388
R21472 GND.n1473 GND.n1472 3.388
R21473 GND.n1561 GND.n1560 3.388
R21474 GND.n1356 GND.n1355 3.388
R21475 GND.n1444 GND.n1443 3.388
R21476 GND.n1239 GND.n1238 3.388
R21477 GND.n1327 GND.n1326 3.388
R21478 GND.n1122 GND.n1121 3.388
R21479 GND.n1210 GND.n1209 3.388
R21480 GND.n1006 GND.n1005 3.388
R21481 GND.n1094 GND.n1093 3.388
R21482 GND.n2906 GND.n2903 3.388
R21483 GND.n2842 GND.n2841 3.388
R21484 GND.n2769 GND.n2768 3.388
R21485 GND.n2720 GND.n2719 3.388
R21486 GND.n652 GND.n651 3.318
R21487 GND.n690 GND.n689 3.318
R21488 GND.n574 GND.n453 3.294
R21489 GND.n332 GND.n1 3.206
R21490 GND.n2551 GND.n2550 3.081
R21491 GND.n2670 GND.n2669 3.081
R21492 GND.n2562 GND.n2561 3.081
R21493 GND.n139 GND.n137 3.011
R21494 GND.n147 GND.n144 3.011
R21495 GND.n227 GND.n225 3.011
R21496 GND.n771 GND.n769 3.011
R21497 GND.n779 GND.n776 3.011
R21498 GND.n859 GND.n857 3.011
R21499 GND.n23 GND.n21 3.011
R21500 GND.n31 GND.n28 3.011
R21501 GND.n111 GND.n109 3.011
R21502 GND.n889 GND.n887 3.011
R21503 GND.n897 GND.n894 3.011
R21504 GND.n977 GND.n975 3.011
R21505 GND.n2175 GND.n2173 3.011
R21506 GND.n2183 GND.n2180 3.011
R21507 GND.n2263 GND.n2261 3.011
R21508 GND.n2058 GND.n2056 3.011
R21509 GND.n2066 GND.n2063 3.011
R21510 GND.n2146 GND.n2144 3.011
R21511 GND.n1941 GND.n1939 3.011
R21512 GND.n1949 GND.n1946 3.011
R21513 GND.n2029 GND.n2027 3.011
R21514 GND.n1824 GND.n1822 3.011
R21515 GND.n1832 GND.n1829 3.011
R21516 GND.n1912 GND.n1910 3.011
R21517 GND.n1707 GND.n1705 3.011
R21518 GND.n1715 GND.n1712 3.011
R21519 GND.n1795 GND.n1793 3.011
R21520 GND.n1590 GND.n1588 3.011
R21521 GND.n1598 GND.n1595 3.011
R21522 GND.n1678 GND.n1676 3.011
R21523 GND.n1473 GND.n1471 3.011
R21524 GND.n1481 GND.n1478 3.011
R21525 GND.n1561 GND.n1559 3.011
R21526 GND.n1356 GND.n1354 3.011
R21527 GND.n1364 GND.n1361 3.011
R21528 GND.n1444 GND.n1442 3.011
R21529 GND.n1239 GND.n1237 3.011
R21530 GND.n1247 GND.n1244 3.011
R21531 GND.n1327 GND.n1325 3.011
R21532 GND.n1122 GND.n1120 3.011
R21533 GND.n1130 GND.n1127 3.011
R21534 GND.n1210 GND.n1208 3.011
R21535 GND.n1006 GND.n1004 3.011
R21536 GND.n1014 GND.n1011 3.011
R21537 GND.n1094 GND.n1092 3.011
R21538 GND.n2986 GND.n2984 3.011
R21539 GND.n2906 GND.n2905 3.011
R21540 GND.n2842 GND.n2839 3.011
R21541 GND.n2810 GND.n2808 3.011
R21542 GND.n2758 GND.n2757 3.011
R21543 GND.n2769 GND.n2767 3.011
R21544 GND.n2720 GND.n2718 3.011
R21545 GND.n2330 GND.n2329 2.909
R21546 GND.n2342 GND.n2341 2.909
R21547 GND.n638 GND.n637 2.844
R21548 GND.n704 GND.n703 2.844
R21549 GND.n161 GND.n160 2.635
R21550 GND.n205 GND.n204 2.635
R21551 GND.n216 GND.n215 2.635
R21552 GND.n793 GND.n792 2.635
R21553 GND.n837 GND.n836 2.635
R21554 GND.n848 GND.n847 2.635
R21555 GND.n45 GND.n44 2.635
R21556 GND.n89 GND.n88 2.635
R21557 GND.n100 GND.n99 2.635
R21558 GND.n911 GND.n910 2.635
R21559 GND.n955 GND.n954 2.635
R21560 GND.n966 GND.n965 2.635
R21561 GND.n2197 GND.n2196 2.635
R21562 GND.n2241 GND.n2240 2.635
R21563 GND.n2252 GND.n2251 2.635
R21564 GND.n2080 GND.n2079 2.635
R21565 GND.n2124 GND.n2123 2.635
R21566 GND.n2135 GND.n2134 2.635
R21567 GND.n1963 GND.n1962 2.635
R21568 GND.n2007 GND.n2006 2.635
R21569 GND.n2018 GND.n2017 2.635
R21570 GND.n1846 GND.n1845 2.635
R21571 GND.n1890 GND.n1889 2.635
R21572 GND.n1901 GND.n1900 2.635
R21573 GND.n1729 GND.n1728 2.635
R21574 GND.n1773 GND.n1772 2.635
R21575 GND.n1784 GND.n1783 2.635
R21576 GND.n1612 GND.n1611 2.635
R21577 GND.n1656 GND.n1655 2.635
R21578 GND.n1667 GND.n1666 2.635
R21579 GND.n1495 GND.n1494 2.635
R21580 GND.n1539 GND.n1538 2.635
R21581 GND.n1550 GND.n1549 2.635
R21582 GND.n1378 GND.n1377 2.635
R21583 GND.n1422 GND.n1421 2.635
R21584 GND.n1433 GND.n1432 2.635
R21585 GND.n1261 GND.n1260 2.635
R21586 GND.n1305 GND.n1304 2.635
R21587 GND.n1316 GND.n1315 2.635
R21588 GND.n1144 GND.n1143 2.635
R21589 GND.n1188 GND.n1187 2.635
R21590 GND.n1199 GND.n1198 2.635
R21591 GND.n1028 GND.n1027 2.635
R21592 GND.n1072 GND.n1071 2.635
R21593 GND.n1083 GND.n1082 2.635
R21594 GND.n2963 GND.n2962 2.635
R21595 GND.n2856 GND.n2855 2.635
R21596 GND.n2860 GND.n2859 2.635
R21597 GND.n2799 GND.n2798 2.635
R21598 GND.n2787 GND.n2786 2.635
R21599 GND.n589 GND.n579 2.607
R21600 GND.n300 GND.n289 2.607
R21601 GND.n493 GND.n491 2.607
R21602 GND.n453 GND.n441 2.607
R21603 GND.n2318 GND.n2317 2.521
R21604 GND.n2355 GND.n2354 2.521
R21605 GND.n3000 GND.n2999 2.46
R21606 GND.n624 GND.n623 2.37
R21607 GND.n718 GND.n717 2.37
R21608 GND.n266 GND.n256 2.37
R21609 GND.n258 GND.n257 2.37
R21610 GND.n467 GND.n466 2.37
R21611 GND.n473 GND.n471 2.37
R21612 GND.n532 GND.n531 2.37
R21613 GND.n541 GND.n540 2.37
R21614 GND.n550 GND.n549 2.37
R21615 GND.n2646 GND.n2644 2.37
R21616 GND.n2475 GND.n2473 2.37
R21617 GND.n2882 GND.n2881 2.258
R21618 GND.n2740 GND.n2738 2.258
R21619 GND.n3049 GND.n3048 2.25
R21620 GND.n3016 GND.n3015 2.25
R21621 GND.n2668 GND.n2667 2.25
R21622 GND.n2497 GND.n2496 2.25
R21623 GND.n3047 GND.n3046 2.246
R21624 GND.n3024 GND.n3023 2.246
R21625 GND.n3050 GND.n3039 2.245
R21626 GND.n3014 GND.n3013 2.245
R21627 GND.n2999 GND.n2998 2.219
R21628 GND.n2560 GND.n2392 2.178
R21629 GND.n617 GND.n610 2.133
R21630 GND.n739 GND.n732 2.133
R21631 GND.n326 GND.n325 2.133
R21632 GND.n325 GND.n318 2.133
R21633 GND.n278 GND.n267 2.133
R21634 GND.n481 GND.n480 2.133
R21635 GND.n502 GND.n501 2.133
R21636 GND.n512 GND.n510 2.133
R21637 GND.n566 GND.n559 2.133
R21638 GND.n568 GND.n566 2.133
R21639 GND.n2305 GND.n2304 2.133
R21640 GND.n2367 GND.n2366 2.133
R21641 GND.n2602 GND.n2601 2.133
R21642 GND.n2428 GND.n2427 2.133
R21643 GND.n2347 GND.n2346 1.956
R21644 GND.n2372 GND.n2371 1.956
R21645 GND.n2310 GND.n2309 1.956
R21646 GND.n2335 GND.n2334 1.956
R21647 GND.n2287 GND.n2282 1.939
R21648 GND.n2280 GND.n2274 1.939
R21649 GND.n610 GND.n609 1.896
R21650 GND.n732 GND.n731 1.896
R21651 GND.n326 GND.n316 1.896
R21652 GND.n318 GND.n317 1.896
R21653 GND.n278 GND.n277 1.896
R21654 GND.n269 GND.n268 1.896
R21655 GND.n512 GND.n511 1.896
R21656 GND.n559 GND.n558 1.896
R21657 GND.n568 GND.n567 1.896
R21658 GND.n2602 GND.n2593 1.896
R21659 GND.n2608 GND.n2606 1.896
R21660 GND.n2654 GND.n2653 1.896
R21661 GND.n2428 GND.n2419 1.896
R21662 GND.n2435 GND.n2433 1.896
R21663 GND.n2483 GND.n2482 1.896
R21664 GND.n2293 GND.n2292 1.745
R21665 GND.n2380 GND.n2379 1.745
R21666 GND.n3060 GND.n3059 1.706
R21667 GND.n3096 GND.n3095 1.706
R21668 GND.n631 GND.n624 1.659
R21669 GND.n725 GND.n718 1.659
R21670 GND.n266 GND.n265 1.659
R21671 GND.n265 GND.n258 1.659
R21672 GND.n467 GND.n458 1.659
R21673 GND.n522 GND.n521 1.659
R21674 GND.n532 GND.n530 1.659
R21675 GND.n548 GND.n541 1.659
R21676 GND.n550 GND.n548 1.659
R21677 GND.n2572 GND.n2571 1.659
R21678 GND.n2631 GND.n2630 1.659
R21679 GND.n2646 GND.n2645 1.659
R21680 GND.n2401 GND.n2400 1.659
R21681 GND.n2460 GND.n2459 1.659
R21682 GND.n2475 GND.n2474 1.659
R21683 GND.n2298 GND.n2293 1.551
R21684 GND.n2385 GND.n2380 1.551
R21685 GND.n2963 GND.n2961 1.505
R21686 GND.n2799 GND.n2797 1.505
R21687 GND.n230 GND.n229 1.5
R21688 GND.n163 GND.n162 1.5
R21689 GND.n862 GND.n861 1.5
R21690 GND.n795 GND.n794 1.5
R21691 GND.n114 GND.n113 1.5
R21692 GND.n47 GND.n46 1.5
R21693 GND.n980 GND.n979 1.5
R21694 GND.n913 GND.n912 1.5
R21695 GND.n2266 GND.n2265 1.5
R21696 GND.n2199 GND.n2198 1.5
R21697 GND.n2149 GND.n2148 1.5
R21698 GND.n2082 GND.n2081 1.5
R21699 GND.n2032 GND.n2031 1.5
R21700 GND.n1965 GND.n1964 1.5
R21701 GND.n1915 GND.n1914 1.5
R21702 GND.n1848 GND.n1847 1.5
R21703 GND.n1798 GND.n1797 1.5
R21704 GND.n1731 GND.n1730 1.5
R21705 GND.n1681 GND.n1680 1.5
R21706 GND.n1614 GND.n1613 1.5
R21707 GND.n1564 GND.n1563 1.5
R21708 GND.n1497 GND.n1496 1.5
R21709 GND.n1447 GND.n1446 1.5
R21710 GND.n1380 GND.n1379 1.5
R21711 GND.n1330 GND.n1329 1.5
R21712 GND.n1263 GND.n1262 1.5
R21713 GND.n1213 GND.n1212 1.5
R21714 GND.n1146 GND.n1145 1.5
R21715 GND.n1097 GND.n1096 1.5
R21716 GND.n1030 GND.n1029 1.5
R21717 GND.n2706 GND.n2704 1.5
R21718 GND.n2726 GND.n2725 1.5
R21719 GND.n2889 GND.n2888 1.5
R21720 GND.n2925 GND.n2924 1.5
R21721 GND.n2865 GND.n2864 1.5
R21722 GND.n2844 GND.n2843 1.5
R21723 GND.n2814 GND.n2813 1.5
R21724 GND.n2829 GND.n2828 1.5
R21725 GND.n2803 GND.n2802 1.5
R21726 GND.n2819 GND.n2818 1.5
R21727 GND.n2793 GND.n2792 1.5
R21728 GND.n2771 GND.n2770 1.5
R21729 GND.n2745 GND.n2744 1.5
R21730 GND.n2908 GND.n2907 1.5
R21731 GND.n2615 GND.n2614 1.5
R21732 GND.n2633 GND.n2632 1.5
R21733 GND.n2622 GND.n2621 1.5
R21734 GND.n2648 GND.n2647 1.5
R21735 GND.n2610 GND.n2609 1.5
R21736 GND.n2604 GND.n2603 1.5
R21737 GND.n2666 GND.n2665 1.5
R21738 GND.n2586 GND.n2585 1.5
R21739 GND.n2495 GND.n2494 1.5
R21740 GND.n2451 GND.n2450 1.5
R21741 GND.n2444 GND.n2443 1.5
R21742 GND.n2462 GND.n2461 1.5
R21743 GND.n2437 GND.n2436 1.5
R21744 GND.n2431 GND.n2430 1.5
R21745 GND.n2477 GND.n2476 1.5
R21746 GND.n2413 GND.n2412 1.5
R21747 GND.n579 GND.n578 1.422
R21748 GND.n300 GND.n299 1.422
R21749 GND.n292 GND.n291 1.422
R21750 GND.n291 GND.n290 1.422
R21751 GND.n270 GND.n269 1.422
R21752 GND.n493 GND.n492 1.422
R21753 GND.n441 GND.n440 1.422
R21754 GND.n2573 GND.n2572 1.422
R21755 GND.n2402 GND.n2401 1.422
R21756 GND.n2971 GND.n2970 1.399
R21757 GND.n2996 GND.n2993 1.395
R21758 GND.n2282 GND.n2281 1.357
R21759 GND.n2274 GND.n2273 1.357
R21760 GND.n3083 GND.n3082 1.254
R21761 GND.n645 GND.n638 1.185
R21762 GND.n711 GND.n704 1.185
R21763 GND.n299 GND.n292 1.185
R21764 GND.n481 GND.n478 1.185
R21765 GND.n503 GND.n502 1.185
R21766 GND.n523 GND.n522 1.185
R21767 GND.n530 GND.n523 1.185
R21768 GND.n3045 GND.n3044 1.185
R21769 GND.n3018 GND.n3017 1.185
R21770 GND.n2655 GND.n2654 1.185
R21771 GND.n2484 GND.n2483 1.185
R21772 GND.n2311 GND.n2305 1.163
R21773 GND.n2373 GND.n2367 1.163
R21774 GND.n336 GND.n335 1.142
R21775 GND.n3088 GND.n3087 1.138
R21776 GND.n576 GND.n575 1.137
R21777 GND.n355 GND.n354 1.137
R21778 GND.n365 GND.n364 1.137
R21779 GND.n372 GND.n371 1.137
R21780 GND.n380 GND.n379 1.137
R21781 GND.n386 GND.n385 1.137
R21782 GND.n391 GND.n390 1.137
R21783 GND.n399 GND.n398 1.137
R21784 GND.n408 GND.n407 1.137
R21785 GND.n415 GND.n414 1.137
R21786 GND.n424 GND.n423 1.137
R21787 GND.n429 GND.n428 1.137
R21788 GND.n435 GND.n434 1.137
R21789 GND.n347 GND.n346 1.137
R21790 GND.n341 GND.n340 1.137
R21791 GND.n2997 GND.n2996 1.137
R21792 GND.n2980 GND.n2979 1.137
R21793 GND.n2708 GND.n2707 1.137
R21794 GND.n2728 GND.n2727 1.137
R21795 GND.n2747 GND.n2746 1.137
R21796 GND.n2755 GND.n2754 1.137
R21797 GND.n2773 GND.n2772 1.137
R21798 GND.n2780 GND.n2779 1.137
R21799 GND.n2873 GND.n2872 1.137
R21800 GND.n2931 GND.n2930 1.137
R21801 GND.n2894 GND.n2893 1.137
R21802 GND.n2848 GND.n2847 1.137
R21803 GND.n2869 GND.n2868 1.137
R21804 GND.n2831 GND.n2830 1.137
R21805 GND.n2807 GND.n2806 1.137
R21806 GND.n2915 GND.n2914 1.137
R21807 GND.n3085 GND.n3084 1.137
R21808 GND.n3066 GND.n3065 1.137
R21809 GND.n3104 GND.n3103 1.137
R21810 GND.n3123 GND.n3122 1.137
R21811 GND.n3125 GND.n3124 1.135
R21812 GND.n2986 GND.n2985 1.129
R21813 GND.n2810 GND.n2809 1.129
R21814 GND.n3058 GND.n3057 1.065
R21815 GND.n3094 GND.n3093 1.065
R21816 GND.n1218 GND.n1101 1.063
R21817 GND.n750 GND.n234 1.037
R21818 GND.n1335 GND.n1334 1.036
R21819 GND.n1569 GND.n1568 1.036
R21820 GND.n1803 GND.n1802 1.036
R21821 GND.n2037 GND.n2036 1.036
R21822 GND.n2271 GND.n2270 1.036
R21823 GND.n868 GND.n118 1.036
R21824 GND.n867 GND.n866 1.034
R21825 GND.n985 GND.n984 1.034
R21826 GND.n2154 GND.n2153 1.034
R21827 GND.n1920 GND.n1919 1.034
R21828 GND.n1686 GND.n1685 1.034
R21829 GND.n1452 GND.n1451 1.034
R21830 GND.n1218 GND.n1217 1.034
R21831 GND.n3121 GND.n3120 0.962
R21832 GND.n473 GND.n472 0.948
R21833 GND.n3038 GND.n3037 0.948
R21834 GND.n3012 GND.n3011 0.948
R21835 GND.n2558 GND.n2551 0.948
R21836 GND.n2672 GND.n2670 0.948
R21837 GND.n2565 GND.n2562 0.948
R21838 GND.n2581 GND.n2573 0.948
R21839 GND.n2631 GND.n2628 0.948
R21840 GND.n2630 GND.n2629 0.948
R21841 GND.n2663 GND.n2655 0.948
R21842 GND.n2410 GND.n2402 0.948
R21843 GND.n2460 GND.n2457 0.948
R21844 GND.n2459 GND.n2458 0.948
R21845 GND.n2492 GND.n2484 0.948
R21846 GND.n575 GND.n574 0.867
R21847 GND.n335 GND.n332 0.866
R21848 GND.n2972 GND.n2971 0.862
R21849 GND.n233 GND.n232 0.853
R21850 GND.n865 GND.n864 0.853
R21851 GND.n117 GND.n116 0.853
R21852 GND.n983 GND.n982 0.853
R21853 GND.n2269 GND.n2268 0.853
R21854 GND.n2152 GND.n2151 0.853
R21855 GND.n2035 GND.n2034 0.853
R21856 GND.n1918 GND.n1917 0.853
R21857 GND.n1801 GND.n1800 0.853
R21858 GND.n1684 GND.n1683 0.853
R21859 GND.n1567 GND.n1566 0.853
R21860 GND.n1450 GND.n1449 0.853
R21861 GND.n1333 GND.n1332 0.853
R21862 GND.n1216 GND.n1215 0.853
R21863 GND.n1100 GND.n1099 0.853
R21864 GND.n746 GND.n745 0.827
R21865 GND.n2323 GND.n2318 0.775
R21866 GND.n2360 GND.n2355 0.775
R21867 GND.n3061 GND.n3060 0.756
R21868 GND.n133 GND.n132 0.752
R21869 GND.n211 GND.n210 0.752
R21870 GND.n765 GND.n764 0.752
R21871 GND.n843 GND.n842 0.752
R21872 GND.n17 GND.n16 0.752
R21873 GND.n95 GND.n94 0.752
R21874 GND.n883 GND.n882 0.752
R21875 GND.n961 GND.n960 0.752
R21876 GND.n2169 GND.n2168 0.752
R21877 GND.n2247 GND.n2246 0.752
R21878 GND.n2052 GND.n2051 0.752
R21879 GND.n2130 GND.n2129 0.752
R21880 GND.n1935 GND.n1934 0.752
R21881 GND.n2013 GND.n2012 0.752
R21882 GND.n1818 GND.n1817 0.752
R21883 GND.n1896 GND.n1895 0.752
R21884 GND.n1701 GND.n1700 0.752
R21885 GND.n1779 GND.n1778 0.752
R21886 GND.n1584 GND.n1583 0.752
R21887 GND.n1662 GND.n1661 0.752
R21888 GND.n1467 GND.n1466 0.752
R21889 GND.n1545 GND.n1544 0.752
R21890 GND.n1350 GND.n1349 0.752
R21891 GND.n1428 GND.n1427 0.752
R21892 GND.n1233 GND.n1232 0.752
R21893 GND.n1311 GND.n1310 0.752
R21894 GND.n1116 GND.n1115 0.752
R21895 GND.n1194 GND.n1193 0.752
R21896 GND.n1000 GND.n999 0.752
R21897 GND.n1078 GND.n1077 0.752
R21898 GND.n659 GND.n652 0.711
R21899 GND.n697 GND.n690 0.711
R21900 GND.n277 GND.n270 0.711
R21901 GND.n510 GND.n503 0.711
R21902 GND.n2608 GND.n2607 0.711
R21903 GND.n2435 GND.n2434 0.711
R21904 GND.n165 GND.n164 0.702
R21905 GND.n797 GND.n796 0.702
R21906 GND.n49 GND.n48 0.702
R21907 GND.n915 GND.n914 0.702
R21908 GND.n2201 GND.n2200 0.702
R21909 GND.n2084 GND.n2083 0.702
R21910 GND.n1967 GND.n1966 0.702
R21911 GND.n1850 GND.n1849 0.702
R21912 GND.n1733 GND.n1732 0.702
R21913 GND.n1616 GND.n1615 0.702
R21914 GND.n1499 GND.n1498 0.702
R21915 GND.n1382 GND.n1381 0.702
R21916 GND.n1265 GND.n1264 0.702
R21917 GND.n1148 GND.n1147 0.702
R21918 GND.n1032 GND.n1031 0.702
R21919 GND.n3127 GND.n3126 0.654
R21920 GND.n3097 GND.n3096 0.654
R21921 GND.n748 GND.n747 0.563
R21922 GND.n748 GND.n244 0.482
R21923 GND.n480 GND.n479 0.474
R21924 GND.n2530 GND.n2523 0.474
R21925 GND.n2544 GND.n2537 0.474
R21926 GND.n2681 GND.n2679 0.474
R21927 GND.n2689 GND.n2687 0.474
R21928 GND.n2601 GND.n2594 0.474
R21929 GND.n2427 GND.n2420 0.474
R21930 GND.n2286 GND.n2285 0.445
R21931 GND.n2336 GND.n2330 0.387
R21932 GND.n2348 GND.n2342 0.387
R21933 GND.n2297 GND.n2296 0.36
R21934 GND.n2384 GND.n2383 0.36
R21935 GND.n673 GND.n666 0.237
R21936 GND.n683 GND.n676 0.237
R21937 GND.n466 GND.n459 0.237
R21938 GND.n3036 GND.n3027 0.237
R21939 GND.n3043 GND.n3040 0.237
R21940 GND.n3010 GND.n3001 0.237
R21941 GND.n3022 GND.n3019 0.237
R21942 GND.n3074 GND.n3069 0.237
R21943 GND.n3081 GND.n3076 0.237
R21944 GND.n3119 GND.n3114 0.237
R21945 GND.n3112 GND.n3107 0.237
R21946 GND.n3053 GND.n3052 0.215
R21947 GND GND.n3127 0.191
R21948 GND.n2322 GND.n2321 0.184
R21949 GND.n2359 GND.n2358 0.184
R21950 GND.n2685 GND.n2682 0.162
R21951 GND.n2690 GND.n2685 0.162
R21952 GND.n2535 GND.n2531 0.159
R21953 GND.n2545 GND.n2535 0.159
R21954 GND.n2918 GND.n2917 0.155
R21955 GND.n2702 GND.n2701 0.155
R21956 GND.n2567 GND.n2566 0.148
R21957 GND.n2568 GND.n2567 0.148
R21958 GND.n2569 GND.n2568 0.148
R21959 GND.n2668 GND.n2569 0.148
R21960 GND.n2394 GND.n2393 0.148
R21961 GND.n2395 GND.n2394 0.148
R21962 GND.n3054 GND.n2272 0.147
R21963 GND.n2396 GND.n2395 0.147
R21964 GND.n2497 GND.n2396 0.145
R21965 GND.n2905 GND.n2904 0.144
R21966 GND.n2718 GND.n2717 0.144
R21967 GND.n2675 GND.n2673 0.136
R21968 GND.n2695 GND.n2694 0.136
R21969 GND.n2519 GND.n2517 0.134
R21970 GND.n2559 GND.n2549 0.134
R21971 GND.n2881 GND.n2880 0.133
R21972 GND.n2738 GND.n2737 0.132
R21973 GND.n684 GND.n674 0.132
R21974 GND.n2340 GND.n2337 0.132
R21975 GND.n2349 GND.n2340 0.132
R21976 GND.n745 GND.n744 0.115
R21977 GND.n2391 GND.n2390 0.115
R21978 GND.n3054 GND.n3053 0.108
R21979 GND.n620 GND.n618 0.1
R21980 GND.n634 GND.n632 0.1
R21981 GND.n648 GND.n646 0.1
R21982 GND.n662 GND.n660 0.1
R21983 GND.n698 GND.n688 0.1
R21984 GND.n712 GND.n702 0.1
R21985 GND.n726 GND.n716 0.1
R21986 GND.n740 GND.n730 0.1
R21987 GND.n2301 GND.n2299 0.1
R21988 GND.n2314 GND.n2312 0.1
R21989 GND.n2326 GND.n2324 0.1
R21990 GND.n2361 GND.n2353 0.1
R21991 GND.n2374 GND.n2365 0.1
R21992 GND.n2386 GND.n2378 0.1
R21993 GND GND.n3054 0.098
R21994 GND.n3084 GND.n3083 0.056
R21995 GND.n2614 GND.n2612 0.053
R21996 GND.n3122 GND.n3121 0.052
R21997 GND.n2861 GND.n2858 0.051
R21998 GND.n2632 GND.n2626 0.048
R21999 GND.n2443 GND.n2441 0.048
R22000 GND.n2461 GND.n2455 0.048
R22001 GND.n331 GND.n330 0.047
R22002 GND.n312 GND.n311 0.047
R22003 GND.n305 GND.n304 0.047
R22004 GND.n537 GND.n536 0.047
R22005 GND.n555 GND.n554 0.047
R22006 GND.n573 GND.n572 0.047
R22007 GND.n2802 GND.n2796 0.046
R22008 GND.n2846 GND.n2845 0.045
R22009 GND.n2830 GND.n2829 0.045
R22010 GND.n2931 GND.n2915 0.045
R22011 GND.n2831 GND.n2807 0.045
R22012 GND.n2728 GND.n2708 0.045
R22013 GND.n2813 GND.n2812 0.044
R22014 GND.n2745 GND.n2733 0.043
R22015 GND.n2885 GND.n2884 0.042
R22016 GND.n2790 GND.n2789 0.042
R22017 GND.n2726 GND.n2713 0.041
R22018 GND.n2722 GND.n2721 0.04
R22019 GND.n2930 GND.n2929 0.039
R22020 GND.n2707 GND.n2697 0.037
R22021 GND.n2992 GND.n2991 0.036
R22022 GND.n2969 GND.n2968 0.036
R22023 GND.n332 GND.n331 0.035
R22024 GND.n141 GND.n140 0.035
R22025 GND.n201 GND.n200 0.035
R22026 GND.n120 GND.n119 0.035
R22027 GND.n182 GND.n181 0.035
R22028 GND.n773 GND.n772 0.035
R22029 GND.n833 GND.n832 0.035
R22030 GND.n752 GND.n751 0.035
R22031 GND.n814 GND.n813 0.035
R22032 GND.n25 GND.n24 0.035
R22033 GND.n85 GND.n84 0.035
R22034 GND.n4 GND.n3 0.035
R22035 GND.n66 GND.n65 0.035
R22036 GND.n891 GND.n890 0.035
R22037 GND.n951 GND.n950 0.035
R22038 GND.n870 GND.n869 0.035
R22039 GND.n932 GND.n931 0.035
R22040 GND.n2177 GND.n2176 0.035
R22041 GND.n2237 GND.n2236 0.035
R22042 GND.n2156 GND.n2155 0.035
R22043 GND.n2218 GND.n2217 0.035
R22044 GND.n2060 GND.n2059 0.035
R22045 GND.n2120 GND.n2119 0.035
R22046 GND.n2039 GND.n2038 0.035
R22047 GND.n2101 GND.n2100 0.035
R22048 GND.n1943 GND.n1942 0.035
R22049 GND.n2003 GND.n2002 0.035
R22050 GND.n1922 GND.n1921 0.035
R22051 GND.n1984 GND.n1983 0.035
R22052 GND.n1826 GND.n1825 0.035
R22053 GND.n1886 GND.n1885 0.035
R22054 GND.n1805 GND.n1804 0.035
R22055 GND.n1867 GND.n1866 0.035
R22056 GND.n1709 GND.n1708 0.035
R22057 GND.n1769 GND.n1768 0.035
R22058 GND.n1688 GND.n1687 0.035
R22059 GND.n1750 GND.n1749 0.035
R22060 GND.n1592 GND.n1591 0.035
R22061 GND.n1652 GND.n1651 0.035
R22062 GND.n1571 GND.n1570 0.035
R22063 GND.n1633 GND.n1632 0.035
R22064 GND.n1475 GND.n1474 0.035
R22065 GND.n1535 GND.n1534 0.035
R22066 GND.n1454 GND.n1453 0.035
R22067 GND.n1516 GND.n1515 0.035
R22068 GND.n1358 GND.n1357 0.035
R22069 GND.n1418 GND.n1417 0.035
R22070 GND.n1337 GND.n1336 0.035
R22071 GND.n1399 GND.n1398 0.035
R22072 GND.n1241 GND.n1240 0.035
R22073 GND.n1301 GND.n1300 0.035
R22074 GND.n1220 GND.n1219 0.035
R22075 GND.n1282 GND.n1281 0.035
R22076 GND.n1124 GND.n1123 0.035
R22077 GND.n1184 GND.n1183 0.035
R22078 GND.n1103 GND.n1102 0.035
R22079 GND.n1165 GND.n1164 0.035
R22080 GND.n1008 GND.n1007 0.035
R22081 GND.n1068 GND.n1067 0.035
R22082 GND.n987 GND.n986 0.035
R22083 GND.n1049 GND.n1048 0.035
R22084 GND.n476 GND.n475 0.035
R22085 GND.n477 GND.n476 0.035
R22086 GND.n497 GND.n496 0.035
R22087 GND.n346 GND.n343 0.035
R22088 GND.n390 GND.n387 0.035
R22089 GND.n398 GND.n397 0.035
R22090 GND.n2949 GND.n2948 0.035
R22091 GND.n2958 GND.n2957 0.035
R22092 GND.n2936 GND.n2935 0.035
R22093 GND.n2941 GND.n2940 0.035
R22094 GND.n2922 GND.n2921 0.035
R22095 GND.n130 GND.n129 0.034
R22096 GND.n191 GND.n190 0.034
R22097 GND.n762 GND.n761 0.034
R22098 GND.n823 GND.n822 0.034
R22099 GND.n14 GND.n13 0.034
R22100 GND.n75 GND.n74 0.034
R22101 GND.n880 GND.n879 0.034
R22102 GND.n941 GND.n940 0.034
R22103 GND.n2166 GND.n2165 0.034
R22104 GND.n2227 GND.n2226 0.034
R22105 GND.n2049 GND.n2048 0.034
R22106 GND.n2110 GND.n2109 0.034
R22107 GND.n1932 GND.n1931 0.034
R22108 GND.n1993 GND.n1992 0.034
R22109 GND.n1815 GND.n1814 0.034
R22110 GND.n1876 GND.n1875 0.034
R22111 GND.n1698 GND.n1697 0.034
R22112 GND.n1759 GND.n1758 0.034
R22113 GND.n1581 GND.n1580 0.034
R22114 GND.n1642 GND.n1641 0.034
R22115 GND.n1464 GND.n1463 0.034
R22116 GND.n1525 GND.n1524 0.034
R22117 GND.n1347 GND.n1346 0.034
R22118 GND.n1408 GND.n1407 0.034
R22119 GND.n1230 GND.n1229 0.034
R22120 GND.n1291 GND.n1290 0.034
R22121 GND.n1113 GND.n1112 0.034
R22122 GND.n1174 GND.n1173 0.034
R22123 GND.n997 GND.n996 0.034
R22124 GND.n1058 GND.n1057 0.034
R22125 GND.n456 GND.n455 0.034
R22126 GND.n499 GND.n498 0.034
R22127 GND.n379 GND.n376 0.034
R22128 GND.n2928 GND.n2927 0.034
R22129 GND.n2821 GND.n2820 0.034
R22130 GND.n2712 GND.n2711 0.034
R22131 GND.n2677 GND.n2675 0.034
R22132 GND.n2694 GND.n2692 0.034
R22133 GND.n2521 GND.n2519 0.034
R22134 GND.n2549 GND.n2547 0.034
R22135 GND.n574 GND.n573 0.034
R22136 GND.n2699 GND.n2698 0.033
R22137 GND.n220 GND.n219 0.032
R22138 GND.n189 GND.n188 0.032
R22139 GND.n852 GND.n851 0.032
R22140 GND.n821 GND.n820 0.032
R22141 GND.n104 GND.n103 0.032
R22142 GND.n73 GND.n72 0.032
R22143 GND.n970 GND.n969 0.032
R22144 GND.n939 GND.n938 0.032
R22145 GND.n2256 GND.n2255 0.032
R22146 GND.n2225 GND.n2224 0.032
R22147 GND.n2139 GND.n2138 0.032
R22148 GND.n2108 GND.n2107 0.032
R22149 GND.n2022 GND.n2021 0.032
R22150 GND.n1991 GND.n1990 0.032
R22151 GND.n1905 GND.n1904 0.032
R22152 GND.n1874 GND.n1873 0.032
R22153 GND.n1788 GND.n1787 0.032
R22154 GND.n1757 GND.n1756 0.032
R22155 GND.n1671 GND.n1670 0.032
R22156 GND.n1640 GND.n1639 0.032
R22157 GND.n1554 GND.n1553 0.032
R22158 GND.n1523 GND.n1522 0.032
R22159 GND.n1437 GND.n1436 0.032
R22160 GND.n1406 GND.n1405 0.032
R22161 GND.n1320 GND.n1319 0.032
R22162 GND.n1289 GND.n1288 0.032
R22163 GND.n1203 GND.n1202 0.032
R22164 GND.n1172 GND.n1171 0.032
R22165 GND.n1087 GND.n1086 0.032
R22166 GND.n1056 GND.n1055 0.032
R22167 GND.n403 GND.n402 0.032
R22168 GND.n2925 GND.n2916 0.032
R22169 GND.n2804 GND.n2803 0.032
R22170 GND.n2794 GND.n2793 0.032
R22171 GND.n166 GND.n165 0.031
R22172 GND.n177 GND.n176 0.031
R22173 GND.n798 GND.n797 0.031
R22174 GND.n809 GND.n808 0.031
R22175 GND.n50 GND.n49 0.031
R22176 GND.n61 GND.n60 0.031
R22177 GND.n916 GND.n915 0.031
R22178 GND.n927 GND.n926 0.031
R22179 GND.n2202 GND.n2201 0.031
R22180 GND.n2213 GND.n2212 0.031
R22181 GND.n2085 GND.n2084 0.031
R22182 GND.n2096 GND.n2095 0.031
R22183 GND.n1968 GND.n1967 0.031
R22184 GND.n1979 GND.n1978 0.031
R22185 GND.n1851 GND.n1850 0.031
R22186 GND.n1862 GND.n1861 0.031
R22187 GND.n1734 GND.n1733 0.031
R22188 GND.n1745 GND.n1744 0.031
R22189 GND.n1617 GND.n1616 0.031
R22190 GND.n1628 GND.n1627 0.031
R22191 GND.n1500 GND.n1499 0.031
R22192 GND.n1511 GND.n1510 0.031
R22193 GND.n1383 GND.n1382 0.031
R22194 GND.n1394 GND.n1393 0.031
R22195 GND.n1266 GND.n1265 0.031
R22196 GND.n1277 GND.n1276 0.031
R22197 GND.n1149 GND.n1148 0.031
R22198 GND.n1160 GND.n1159 0.031
R22199 GND.n1033 GND.n1032 0.031
R22200 GND.n1044 GND.n1043 0.031
R22201 GND.n2901 GND.n2900 0.031
R22202 GND.n2764 GND.n2763 0.031
R22203 GND.n154 GND.n153 0.03
R22204 GND.n223 GND.n221 0.03
R22205 GND.n128 GND.n127 0.03
R22206 GND.n187 GND.n186 0.03
R22207 GND.n786 GND.n785 0.03
R22208 GND.n855 GND.n853 0.03
R22209 GND.n760 GND.n759 0.03
R22210 GND.n819 GND.n818 0.03
R22211 GND.n38 GND.n37 0.03
R22212 GND.n107 GND.n105 0.03
R22213 GND.n12 GND.n11 0.03
R22214 GND.n71 GND.n70 0.03
R22215 GND.n904 GND.n903 0.03
R22216 GND.n973 GND.n971 0.03
R22217 GND.n878 GND.n877 0.03
R22218 GND.n937 GND.n936 0.03
R22219 GND.n2190 GND.n2189 0.03
R22220 GND.n2259 GND.n2257 0.03
R22221 GND.n2164 GND.n2163 0.03
R22222 GND.n2223 GND.n2222 0.03
R22223 GND.n2073 GND.n2072 0.03
R22224 GND.n2142 GND.n2140 0.03
R22225 GND.n2047 GND.n2046 0.03
R22226 GND.n2106 GND.n2105 0.03
R22227 GND.n1956 GND.n1955 0.03
R22228 GND.n2025 GND.n2023 0.03
R22229 GND.n1930 GND.n1929 0.03
R22230 GND.n1989 GND.n1988 0.03
R22231 GND.n1839 GND.n1838 0.03
R22232 GND.n1908 GND.n1906 0.03
R22233 GND.n1813 GND.n1812 0.03
R22234 GND.n1872 GND.n1871 0.03
R22235 GND.n1722 GND.n1721 0.03
R22236 GND.n1791 GND.n1789 0.03
R22237 GND.n1696 GND.n1695 0.03
R22238 GND.n1755 GND.n1754 0.03
R22239 GND.n1605 GND.n1604 0.03
R22240 GND.n1674 GND.n1672 0.03
R22241 GND.n1579 GND.n1578 0.03
R22242 GND.n1638 GND.n1637 0.03
R22243 GND.n1488 GND.n1487 0.03
R22244 GND.n1557 GND.n1555 0.03
R22245 GND.n1462 GND.n1461 0.03
R22246 GND.n1521 GND.n1520 0.03
R22247 GND.n1371 GND.n1370 0.03
R22248 GND.n1440 GND.n1438 0.03
R22249 GND.n1345 GND.n1344 0.03
R22250 GND.n1404 GND.n1403 0.03
R22251 GND.n1254 GND.n1253 0.03
R22252 GND.n1323 GND.n1321 0.03
R22253 GND.n1228 GND.n1227 0.03
R22254 GND.n1287 GND.n1286 0.03
R22255 GND.n1137 GND.n1136 0.03
R22256 GND.n1206 GND.n1204 0.03
R22257 GND.n1111 GND.n1110 0.03
R22258 GND.n1170 GND.n1169 0.03
R22259 GND.n1021 GND.n1020 0.03
R22260 GND.n1090 GND.n1088 0.03
R22261 GND.n995 GND.n994 0.03
R22262 GND.n1054 GND.n1053 0.03
R22263 GND.n664 GND.n662 0.03
R22264 GND.n688 GND.n686 0.03
R22265 GND.n360 GND.n359 0.03
R22266 GND.n369 GND.n368 0.03
R22267 GND.n750 GND.n749 0.03
R22268 GND.n2946 GND.n2945 0.03
R22269 GND.n2911 GND.n2910 0.03
R22270 GND.n2844 GND.n2834 0.03
R22271 GND.n2815 GND.n2814 0.03
R22272 GND.n372 GND.n365 0.029
R22273 GND.n415 GND.n408 0.029
R22274 GND.n2715 GND.n2714 0.029
R22275 GND.n2724 GND.n2723 0.029
R22276 GND.n157 GND.n155 0.028
R22277 GND.n143 GND.n142 0.028
R22278 GND.n203 GND.n202 0.028
R22279 GND.n125 GND.n124 0.028
R22280 GND.n122 GND.n121 0.028
R22281 GND.n184 GND.n183 0.028
R22282 GND.n230 GND.n191 0.028
R22283 GND.n789 GND.n787 0.028
R22284 GND.n775 GND.n774 0.028
R22285 GND.n835 GND.n834 0.028
R22286 GND.n757 GND.n756 0.028
R22287 GND.n754 GND.n753 0.028
R22288 GND.n816 GND.n815 0.028
R22289 GND.n862 GND.n823 0.028
R22290 GND.n41 GND.n39 0.028
R22291 GND.n27 GND.n26 0.028
R22292 GND.n87 GND.n86 0.028
R22293 GND.n9 GND.n8 0.028
R22294 GND.n6 GND.n5 0.028
R22295 GND.n68 GND.n67 0.028
R22296 GND.n114 GND.n75 0.028
R22297 GND.n907 GND.n905 0.028
R22298 GND.n893 GND.n892 0.028
R22299 GND.n953 GND.n952 0.028
R22300 GND.n875 GND.n874 0.028
R22301 GND.n872 GND.n871 0.028
R22302 GND.n934 GND.n933 0.028
R22303 GND.n980 GND.n941 0.028
R22304 GND.n2193 GND.n2191 0.028
R22305 GND.n2179 GND.n2178 0.028
R22306 GND.n2239 GND.n2238 0.028
R22307 GND.n2161 GND.n2160 0.028
R22308 GND.n2158 GND.n2157 0.028
R22309 GND.n2220 GND.n2219 0.028
R22310 GND.n2266 GND.n2227 0.028
R22311 GND.n2076 GND.n2074 0.028
R22312 GND.n2062 GND.n2061 0.028
R22313 GND.n2122 GND.n2121 0.028
R22314 GND.n2044 GND.n2043 0.028
R22315 GND.n2041 GND.n2040 0.028
R22316 GND.n2103 GND.n2102 0.028
R22317 GND.n2149 GND.n2110 0.028
R22318 GND.n1959 GND.n1957 0.028
R22319 GND.n1945 GND.n1944 0.028
R22320 GND.n2005 GND.n2004 0.028
R22321 GND.n1927 GND.n1926 0.028
R22322 GND.n1924 GND.n1923 0.028
R22323 GND.n1986 GND.n1985 0.028
R22324 GND.n2032 GND.n1993 0.028
R22325 GND.n1842 GND.n1840 0.028
R22326 GND.n1828 GND.n1827 0.028
R22327 GND.n1888 GND.n1887 0.028
R22328 GND.n1810 GND.n1809 0.028
R22329 GND.n1807 GND.n1806 0.028
R22330 GND.n1869 GND.n1868 0.028
R22331 GND.n1915 GND.n1876 0.028
R22332 GND.n1725 GND.n1723 0.028
R22333 GND.n1711 GND.n1710 0.028
R22334 GND.n1771 GND.n1770 0.028
R22335 GND.n1693 GND.n1692 0.028
R22336 GND.n1690 GND.n1689 0.028
R22337 GND.n1752 GND.n1751 0.028
R22338 GND.n1798 GND.n1759 0.028
R22339 GND.n1608 GND.n1606 0.028
R22340 GND.n1594 GND.n1593 0.028
R22341 GND.n1654 GND.n1653 0.028
R22342 GND.n1576 GND.n1575 0.028
R22343 GND.n1573 GND.n1572 0.028
R22344 GND.n1635 GND.n1634 0.028
R22345 GND.n1681 GND.n1642 0.028
R22346 GND.n1491 GND.n1489 0.028
R22347 GND.n1477 GND.n1476 0.028
R22348 GND.n1537 GND.n1536 0.028
R22349 GND.n1459 GND.n1458 0.028
R22350 GND.n1456 GND.n1455 0.028
R22351 GND.n1518 GND.n1517 0.028
R22352 GND.n1564 GND.n1525 0.028
R22353 GND.n1374 GND.n1372 0.028
R22354 GND.n1360 GND.n1359 0.028
R22355 GND.n1420 GND.n1419 0.028
R22356 GND.n1342 GND.n1341 0.028
R22357 GND.n1339 GND.n1338 0.028
R22358 GND.n1401 GND.n1400 0.028
R22359 GND.n1447 GND.n1408 0.028
R22360 GND.n1257 GND.n1255 0.028
R22361 GND.n1243 GND.n1242 0.028
R22362 GND.n1303 GND.n1302 0.028
R22363 GND.n1225 GND.n1224 0.028
R22364 GND.n1222 GND.n1221 0.028
R22365 GND.n1284 GND.n1283 0.028
R22366 GND.n1330 GND.n1291 0.028
R22367 GND.n1140 GND.n1138 0.028
R22368 GND.n1126 GND.n1125 0.028
R22369 GND.n1186 GND.n1185 0.028
R22370 GND.n1108 GND.n1107 0.028
R22371 GND.n1105 GND.n1104 0.028
R22372 GND.n1167 GND.n1166 0.028
R22373 GND.n1213 GND.n1174 0.028
R22374 GND.n1024 GND.n1022 0.028
R22375 GND.n1010 GND.n1009 0.028
R22376 GND.n1070 GND.n1069 0.028
R22377 GND.n992 GND.n991 0.028
R22378 GND.n989 GND.n988 0.028
R22379 GND.n1051 GND.n1050 0.028
R22380 GND.n1097 GND.n1058 0.028
R22381 GND.n516 GND.n515 0.028
R22382 GND.n354 GND.n353 0.028
R22383 GND.n407 GND.n406 0.028
R22384 GND.n412 GND.n411 0.028
R22385 GND.n423 GND.n420 0.028
R22386 GND.n434 GND.n431 0.028
R22387 GND.n2960 GND.n2959 0.028
R22388 GND.n2943 GND.n2942 0.028
R22389 GND.n2732 GND.n2731 0.028
R22390 GND.n2895 GND.n2894 0.028
R22391 GND.n2848 GND.n2833 0.028
R22392 GND.n2781 GND.n2780 0.028
R22393 GND.n2747 GND.n2730 0.028
R22394 GND.n2328 GND.n2326 0.028
R22395 GND.n2353 GND.n2351 0.028
R22396 GND.n164 GND.n163 0.028
R22397 GND.n796 GND.n795 0.028
R22398 GND.n48 GND.n47 0.028
R22399 GND.n914 GND.n913 0.028
R22400 GND.n2200 GND.n2199 0.028
R22401 GND.n2083 GND.n2082 0.028
R22402 GND.n1966 GND.n1965 0.028
R22403 GND.n1849 GND.n1848 0.028
R22404 GND.n1732 GND.n1731 0.028
R22405 GND.n1615 GND.n1614 0.028
R22406 GND.n1498 GND.n1497 0.028
R22407 GND.n1381 GND.n1380 0.028
R22408 GND.n1264 GND.n1263 0.028
R22409 GND.n1147 GND.n1146 0.028
R22410 GND.n1031 GND.n1030 0.028
R22411 GND.n170 GND.n169 0.027
R22412 GND.n173 GND.n172 0.027
R22413 GND.n802 GND.n801 0.027
R22414 GND.n805 GND.n804 0.027
R22415 GND.n54 GND.n53 0.027
R22416 GND.n57 GND.n56 0.027
R22417 GND.n920 GND.n919 0.027
R22418 GND.n923 GND.n922 0.027
R22419 GND.n2206 GND.n2205 0.027
R22420 GND.n2209 GND.n2208 0.027
R22421 GND.n2089 GND.n2088 0.027
R22422 GND.n2092 GND.n2091 0.027
R22423 GND.n1972 GND.n1971 0.027
R22424 GND.n1975 GND.n1974 0.027
R22425 GND.n1855 GND.n1854 0.027
R22426 GND.n1858 GND.n1857 0.027
R22427 GND.n1738 GND.n1737 0.027
R22428 GND.n1741 GND.n1740 0.027
R22429 GND.n1621 GND.n1620 0.027
R22430 GND.n1624 GND.n1623 0.027
R22431 GND.n1504 GND.n1503 0.027
R22432 GND.n1507 GND.n1506 0.027
R22433 GND.n1387 GND.n1386 0.027
R22434 GND.n1390 GND.n1389 0.027
R22435 GND.n1270 GND.n1269 0.027
R22436 GND.n1273 GND.n1272 0.027
R22437 GND.n1153 GND.n1152 0.027
R22438 GND.n1156 GND.n1155 0.027
R22439 GND.n1037 GND.n1036 0.027
R22440 GND.n1040 GND.n1039 0.027
R22441 GND.n1335 GND.n1218 0.027
R22442 GND.n1452 GND.n1335 0.027
R22443 GND.n1569 GND.n1452 0.027
R22444 GND.n1686 GND.n1569 0.027
R22445 GND.n1803 GND.n1686 0.027
R22446 GND.n1920 GND.n1803 0.027
R22447 GND.n2037 GND.n1920 0.027
R22448 GND.n2154 GND.n2037 0.027
R22449 GND.n2271 GND.n2154 0.027
R22450 GND.n985 GND.n868 0.027
R22451 GND.n868 GND.n867 0.027
R22452 GND.n867 GND.n750 0.027
R22453 GND.n2621 GND.n2619 0.027
R22454 GND.n2450 GND.n2448 0.027
R22455 GND.n163 GND.n130 0.026
R22456 GND.n795 GND.n762 0.026
R22457 GND.n47 GND.n14 0.026
R22458 GND.n913 GND.n880 0.026
R22459 GND.n2199 GND.n2166 0.026
R22460 GND.n2082 GND.n2049 0.026
R22461 GND.n1965 GND.n1932 0.026
R22462 GND.n1848 GND.n1815 0.026
R22463 GND.n1731 GND.n1698 0.026
R22464 GND.n1614 GND.n1581 0.026
R22465 GND.n1497 GND.n1464 0.026
R22466 GND.n1380 GND.n1347 0.026
R22467 GND.n1263 GND.n1230 0.026
R22468 GND.n1146 GND.n1113 0.026
R22469 GND.n1030 GND.n997 0.026
R22470 GND.n650 GND.n648 0.026
R22471 GND.n702 GND.n700 0.026
R22472 GND.n314 GND.n313 0.026
R22473 GND.n284 GND.n283 0.026
R22474 GND.n518 GND.n517 0.026
R22475 GND.n556 GND.n555 0.026
R22476 GND.n364 GND.n363 0.026
R22477 GND.n371 GND.n367 0.026
R22478 GND.n2899 GND.n2898 0.026
R22479 GND.n2878 GND.n2877 0.026
R22480 GND.n2886 GND.n2885 0.026
R22481 GND.n2743 GND.n2742 0.026
R22482 GND.n2913 GND.n2912 0.026
R22483 GND.n286 GND.n285 0.024
R22484 GND.n536 GND.n535 0.024
R22485 GND.n410 GND.n409 0.024
R22486 GND.n414 GND.n410 0.024
R22487 GND.n428 GND.n427 0.024
R22488 GND.n2888 GND.n2878 0.024
R22489 GND.n2735 GND.n2734 0.024
R22490 GND.n2744 GND.n2743 0.024
R22491 GND.n2893 GND.n2892 0.024
R22492 GND.n2871 GND.n2870 0.024
R22493 GND.n2868 GND.n2867 0.024
R22494 GND.n2779 GND.n2778 0.024
R22495 GND.n2754 GND.n2753 0.024
R22496 GND.n2710 GND.n2709 0.024
R22497 GND.n2873 GND.n2869 0.024
R22498 GND.n2773 GND.n2755 0.024
R22499 GND.n2316 GND.n2314 0.024
R22500 GND.n2365 GND.n2363 0.024
R22501 GND.n3052 GND.n3026 0.024
R22502 GND.n2855 GND.n2854 0.024
R22503 GND.n2767 GND.n2766 0.024
R22504 GND.n2584 GND.n2583 0.023
R22505 GND.n2647 GND.n2634 0.023
R22506 GND.n2636 GND.n2635 0.023
R22507 GND.n2399 GND.n2398 0.023
R22508 GND.n2476 GND.n2463 0.023
R22509 GND.n2465 GND.n2464 0.023
R22510 GND.n199 GND.n195 0.022
R22511 GND.n180 GND.n179 0.022
R22512 GND.n232 GND.n230 0.022
R22513 GND.n831 GND.n827 0.022
R22514 GND.n812 GND.n811 0.022
R22515 GND.n864 GND.n862 0.022
R22516 GND.n83 GND.n79 0.022
R22517 GND.n64 GND.n63 0.022
R22518 GND.n116 GND.n114 0.022
R22519 GND.n949 GND.n945 0.022
R22520 GND.n930 GND.n929 0.022
R22521 GND.n982 GND.n980 0.022
R22522 GND.n2235 GND.n2231 0.022
R22523 GND.n2216 GND.n2215 0.022
R22524 GND.n2268 GND.n2266 0.022
R22525 GND.n2118 GND.n2114 0.022
R22526 GND.n2099 GND.n2098 0.022
R22527 GND.n2151 GND.n2149 0.022
R22528 GND.n2001 GND.n1997 0.022
R22529 GND.n1982 GND.n1981 0.022
R22530 GND.n2034 GND.n2032 0.022
R22531 GND.n1884 GND.n1880 0.022
R22532 GND.n1865 GND.n1864 0.022
R22533 GND.n1917 GND.n1915 0.022
R22534 GND.n1767 GND.n1763 0.022
R22535 GND.n1748 GND.n1747 0.022
R22536 GND.n1800 GND.n1798 0.022
R22537 GND.n1650 GND.n1646 0.022
R22538 GND.n1631 GND.n1630 0.022
R22539 GND.n1683 GND.n1681 0.022
R22540 GND.n1533 GND.n1529 0.022
R22541 GND.n1514 GND.n1513 0.022
R22542 GND.n1566 GND.n1564 0.022
R22543 GND.n1416 GND.n1412 0.022
R22544 GND.n1397 GND.n1396 0.022
R22545 GND.n1449 GND.n1447 0.022
R22546 GND.n1299 GND.n1295 0.022
R22547 GND.n1280 GND.n1279 0.022
R22548 GND.n1332 GND.n1330 0.022
R22549 GND.n1182 GND.n1178 0.022
R22550 GND.n1163 GND.n1162 0.022
R22551 GND.n1215 GND.n1213 0.022
R22552 GND.n1066 GND.n1062 0.022
R22553 GND.n1047 GND.n1046 0.022
R22554 GND.n1099 GND.n1097 0.022
R22555 GND.n636 GND.n634 0.022
R22556 GND.n716 GND.n714 0.022
R22557 GND.n304 GND.n303 0.022
R22558 GND.n285 GND.n284 0.022
R22559 GND.n345 GND.n344 0.022
R22560 GND.n363 GND.n362 0.022
R22561 GND.n367 GND.n366 0.022
R22562 GND.n2956 GND.n2954 0.022
R22563 GND.n2939 GND.n2938 0.022
R22564 GND.n2980 GND.n2976 0.022
R22565 GND.n2974 GND.n2973 0.022
R22566 GND.n2864 GND.n2852 0.022
R22567 GND.n2862 GND.n2861 0.022
R22568 GND.n2771 GND.n2756 0.022
R22569 GND.n239 GND.n238 0.021
R22570 GND.n236 GND.n235 0.021
R22571 GND.n243 GND.n242 0.021
R22572 GND.n244 GND.n241 0.02
R22573 GND.n195 GND.n193 0.02
R22574 GND.n179 GND.n178 0.02
R22575 GND.n827 GND.n825 0.02
R22576 GND.n811 GND.n810 0.02
R22577 GND.n79 GND.n77 0.02
R22578 GND.n63 GND.n62 0.02
R22579 GND.n945 GND.n943 0.02
R22580 GND.n929 GND.n928 0.02
R22581 GND.n2231 GND.n2229 0.02
R22582 GND.n2215 GND.n2214 0.02
R22583 GND.n2114 GND.n2112 0.02
R22584 GND.n2098 GND.n2097 0.02
R22585 GND.n1997 GND.n1995 0.02
R22586 GND.n1981 GND.n1980 0.02
R22587 GND.n1880 GND.n1878 0.02
R22588 GND.n1864 GND.n1863 0.02
R22589 GND.n1763 GND.n1761 0.02
R22590 GND.n1747 GND.n1746 0.02
R22591 GND.n1646 GND.n1644 0.02
R22592 GND.n1630 GND.n1629 0.02
R22593 GND.n1529 GND.n1527 0.02
R22594 GND.n1513 GND.n1512 0.02
R22595 GND.n1412 GND.n1410 0.02
R22596 GND.n1396 GND.n1395 0.02
R22597 GND.n1295 GND.n1293 0.02
R22598 GND.n1279 GND.n1278 0.02
R22599 GND.n1178 GND.n1176 0.02
R22600 GND.n1162 GND.n1161 0.02
R22601 GND.n1062 GND.n1060 0.02
R22602 GND.n1046 GND.n1045 0.02
R22603 GND.n302 GND.n301 0.02
R22604 GND.n494 GND.n484 0.02
R22605 GND.n517 GND.n516 0.02
R22606 GND.n353 GND.n352 0.02
R22607 GND.n406 GND.n405 0.02
R22608 GND.n420 GND.n419 0.02
R22609 GND.n2954 GND.n2951 0.02
R22610 GND.n2938 GND.n2937 0.02
R22611 GND.n2907 GND.n2899 0.02
R22612 GND.n2843 GND.n2838 0.02
R22613 GND.n2827 GND.n2826 0.02
R22614 GND.n2826 GND.n2823 0.02
R22615 GND.n2760 GND.n2759 0.02
R22616 GND.n2770 GND.n2765 0.02
R22617 GND.n2725 GND.n2724 0.02
R22618 GND.n2303 GND.n2301 0.02
R22619 GND.n2378 GND.n2376 0.02
R22620 GND.n2590 GND.n2589 0.02
R22621 GND.n2591 GND.n2590 0.02
R22622 GND.n2603 GND.n2592 0.02
R22623 GND.n2637 GND.n2636 0.02
R22624 GND.n2652 GND.n2651 0.02
R22625 GND.n2417 GND.n2416 0.02
R22626 GND.n2418 GND.n2417 0.02
R22627 GND.n2430 GND.n2429 0.02
R22628 GND.n2466 GND.n2465 0.02
R22629 GND.n2481 GND.n2480 0.02
R22630 GND.n3067 GND.n3066 0.02
R22631 GND.n3085 GND.n3067 0.02
R22632 GND.n3123 GND.n3105 0.02
R22633 GND.n3105 GND.n3104 0.02
R22634 GND.n237 GND.n236 0.02
R22635 GND.n233 GND.n177 0.019
R22636 GND.n234 GND.n233 0.019
R22637 GND.n865 GND.n809 0.019
R22638 GND.n866 GND.n865 0.019
R22639 GND.n117 GND.n61 0.019
R22640 GND.n118 GND.n117 0.019
R22641 GND.n983 GND.n927 0.019
R22642 GND.n984 GND.n983 0.019
R22643 GND.n2269 GND.n2213 0.019
R22644 GND.n2270 GND.n2269 0.019
R22645 GND.n2152 GND.n2096 0.019
R22646 GND.n2153 GND.n2152 0.019
R22647 GND.n2035 GND.n1979 0.019
R22648 GND.n2036 GND.n2035 0.019
R22649 GND.n1918 GND.n1862 0.019
R22650 GND.n1919 GND.n1918 0.019
R22651 GND.n1801 GND.n1745 0.019
R22652 GND.n1802 GND.n1801 0.019
R22653 GND.n1684 GND.n1628 0.019
R22654 GND.n1685 GND.n1684 0.019
R22655 GND.n1567 GND.n1511 0.019
R22656 GND.n1568 GND.n1567 0.019
R22657 GND.n1450 GND.n1394 0.019
R22658 GND.n1451 GND.n1450 0.019
R22659 GND.n1333 GND.n1277 0.019
R22660 GND.n1334 GND.n1333 0.019
R22661 GND.n1216 GND.n1160 0.019
R22662 GND.n1217 GND.n1216 0.019
R22663 GND.n1100 GND.n1044 0.019
R22664 GND.n1101 GND.n1100 0.019
R22665 GND.n162 GND.n131 0.018
R22666 GND.n158 GND.n157 0.018
R22667 GND.n155 GND.n154 0.018
R22668 GND.n217 GND.n208 0.018
R22669 GND.n129 GND.n128 0.018
R22670 GND.n794 GND.n763 0.018
R22671 GND.n790 GND.n789 0.018
R22672 GND.n787 GND.n786 0.018
R22673 GND.n849 GND.n840 0.018
R22674 GND.n761 GND.n760 0.018
R22675 GND.n46 GND.n15 0.018
R22676 GND.n42 GND.n41 0.018
R22677 GND.n39 GND.n38 0.018
R22678 GND.n101 GND.n92 0.018
R22679 GND.n13 GND.n12 0.018
R22680 GND.n912 GND.n881 0.018
R22681 GND.n908 GND.n907 0.018
R22682 GND.n905 GND.n904 0.018
R22683 GND.n967 GND.n958 0.018
R22684 GND.n879 GND.n878 0.018
R22685 GND.n2198 GND.n2167 0.018
R22686 GND.n2194 GND.n2193 0.018
R22687 GND.n2191 GND.n2190 0.018
R22688 GND.n2253 GND.n2244 0.018
R22689 GND.n2165 GND.n2164 0.018
R22690 GND.n2081 GND.n2050 0.018
R22691 GND.n2077 GND.n2076 0.018
R22692 GND.n2074 GND.n2073 0.018
R22693 GND.n2136 GND.n2127 0.018
R22694 GND.n2048 GND.n2047 0.018
R22695 GND.n1964 GND.n1933 0.018
R22696 GND.n1960 GND.n1959 0.018
R22697 GND.n1957 GND.n1956 0.018
R22698 GND.n2019 GND.n2010 0.018
R22699 GND.n1931 GND.n1930 0.018
R22700 GND.n1847 GND.n1816 0.018
R22701 GND.n1843 GND.n1842 0.018
R22702 GND.n1840 GND.n1839 0.018
R22703 GND.n1902 GND.n1893 0.018
R22704 GND.n1814 GND.n1813 0.018
R22705 GND.n1730 GND.n1699 0.018
R22706 GND.n1726 GND.n1725 0.018
R22707 GND.n1723 GND.n1722 0.018
R22708 GND.n1785 GND.n1776 0.018
R22709 GND.n1697 GND.n1696 0.018
R22710 GND.n1613 GND.n1582 0.018
R22711 GND.n1609 GND.n1608 0.018
R22712 GND.n1606 GND.n1605 0.018
R22713 GND.n1668 GND.n1659 0.018
R22714 GND.n1580 GND.n1579 0.018
R22715 GND.n1496 GND.n1465 0.018
R22716 GND.n1492 GND.n1491 0.018
R22717 GND.n1489 GND.n1488 0.018
R22718 GND.n1551 GND.n1542 0.018
R22719 GND.n1463 GND.n1462 0.018
R22720 GND.n1379 GND.n1348 0.018
R22721 GND.n1375 GND.n1374 0.018
R22722 GND.n1372 GND.n1371 0.018
R22723 GND.n1434 GND.n1425 0.018
R22724 GND.n1346 GND.n1345 0.018
R22725 GND.n1262 GND.n1231 0.018
R22726 GND.n1258 GND.n1257 0.018
R22727 GND.n1255 GND.n1254 0.018
R22728 GND.n1317 GND.n1308 0.018
R22729 GND.n1229 GND.n1228 0.018
R22730 GND.n1145 GND.n1114 0.018
R22731 GND.n1141 GND.n1140 0.018
R22732 GND.n1138 GND.n1137 0.018
R22733 GND.n1200 GND.n1191 0.018
R22734 GND.n1112 GND.n1111 0.018
R22735 GND.n1029 GND.n998 0.018
R22736 GND.n1025 GND.n1024 0.018
R22737 GND.n1022 GND.n1021 0.018
R22738 GND.n1084 GND.n1075 0.018
R22739 GND.n996 GND.n995 0.018
R22740 GND.n622 GND.n620 0.018
R22741 GND.n730 GND.n728 0.018
R22742 GND.n309 GND.n308 0.018
R22743 GND.n469 GND.n468 0.018
R22744 GND.n474 GND.n470 0.018
R22745 GND.n534 GND.n533 0.018
R22746 GND.n552 GND.n551 0.018
R22747 GND.n384 GND.n383 0.018
R22748 GND.n356 GND.n355 0.018
R22749 GND.n380 GND.n374 0.018
R22750 GND.n400 GND.n399 0.018
R22751 GND.n424 GND.n417 0.018
R22752 GND.n2967 GND.n2966 0.018
R22753 GND.n2603 GND.n2591 0.018
R22754 GND.n2609 GND.n2605 0.018
R22755 GND.n2665 GND.n2652 0.018
R22756 GND.n2430 GND.n2418 0.018
R22757 GND.n2436 GND.n2432 0.018
R22758 GND.n2494 GND.n2481 0.018
R22759 GND.n2706 GND.n2705 0.017
R22760 GND.n151 GND.n150 0.017
R22761 GND.n221 GND.n220 0.017
R22762 GND.n224 GND.n223 0.017
R22763 GND.n229 GND.n228 0.017
R22764 GND.n127 GND.n126 0.017
R22765 GND.n188 GND.n187 0.017
R22766 GND.n190 GND.n189 0.017
R22767 GND.n783 GND.n782 0.017
R22768 GND.n853 GND.n852 0.017
R22769 GND.n856 GND.n855 0.017
R22770 GND.n861 GND.n860 0.017
R22771 GND.n759 GND.n758 0.017
R22772 GND.n820 GND.n819 0.017
R22773 GND.n822 GND.n821 0.017
R22774 GND.n35 GND.n34 0.017
R22775 GND.n105 GND.n104 0.017
R22776 GND.n108 GND.n107 0.017
R22777 GND.n113 GND.n112 0.017
R22778 GND.n11 GND.n10 0.017
R22779 GND.n72 GND.n71 0.017
R22780 GND.n74 GND.n73 0.017
R22781 GND.n901 GND.n900 0.017
R22782 GND.n971 GND.n970 0.017
R22783 GND.n974 GND.n973 0.017
R22784 GND.n979 GND.n978 0.017
R22785 GND.n877 GND.n876 0.017
R22786 GND.n938 GND.n937 0.017
R22787 GND.n940 GND.n939 0.017
R22788 GND.n2187 GND.n2186 0.017
R22789 GND.n2257 GND.n2256 0.017
R22790 GND.n2260 GND.n2259 0.017
R22791 GND.n2265 GND.n2264 0.017
R22792 GND.n2163 GND.n2162 0.017
R22793 GND.n2224 GND.n2223 0.017
R22794 GND.n2226 GND.n2225 0.017
R22795 GND.n2070 GND.n2069 0.017
R22796 GND.n2140 GND.n2139 0.017
R22797 GND.n2143 GND.n2142 0.017
R22798 GND.n2148 GND.n2147 0.017
R22799 GND.n2046 GND.n2045 0.017
R22800 GND.n2107 GND.n2106 0.017
R22801 GND.n2109 GND.n2108 0.017
R22802 GND.n1953 GND.n1952 0.017
R22803 GND.n2023 GND.n2022 0.017
R22804 GND.n2026 GND.n2025 0.017
R22805 GND.n2031 GND.n2030 0.017
R22806 GND.n1929 GND.n1928 0.017
R22807 GND.n1990 GND.n1989 0.017
R22808 GND.n1992 GND.n1991 0.017
R22809 GND.n1836 GND.n1835 0.017
R22810 GND.n1906 GND.n1905 0.017
R22811 GND.n1909 GND.n1908 0.017
R22812 GND.n1914 GND.n1913 0.017
R22813 GND.n1812 GND.n1811 0.017
R22814 GND.n1873 GND.n1872 0.017
R22815 GND.n1875 GND.n1874 0.017
R22816 GND.n1719 GND.n1718 0.017
R22817 GND.n1789 GND.n1788 0.017
R22818 GND.n1792 GND.n1791 0.017
R22819 GND.n1797 GND.n1796 0.017
R22820 GND.n1695 GND.n1694 0.017
R22821 GND.n1756 GND.n1755 0.017
R22822 GND.n1758 GND.n1757 0.017
R22823 GND.n1602 GND.n1601 0.017
R22824 GND.n1672 GND.n1671 0.017
R22825 GND.n1675 GND.n1674 0.017
R22826 GND.n1680 GND.n1679 0.017
R22827 GND.n1578 GND.n1577 0.017
R22828 GND.n1639 GND.n1638 0.017
R22829 GND.n1641 GND.n1640 0.017
R22830 GND.n1485 GND.n1484 0.017
R22831 GND.n1555 GND.n1554 0.017
R22832 GND.n1558 GND.n1557 0.017
R22833 GND.n1563 GND.n1562 0.017
R22834 GND.n1461 GND.n1460 0.017
R22835 GND.n1522 GND.n1521 0.017
R22836 GND.n1524 GND.n1523 0.017
R22837 GND.n1368 GND.n1367 0.017
R22838 GND.n1438 GND.n1437 0.017
R22839 GND.n1441 GND.n1440 0.017
R22840 GND.n1446 GND.n1445 0.017
R22841 GND.n1344 GND.n1343 0.017
R22842 GND.n1405 GND.n1404 0.017
R22843 GND.n1407 GND.n1406 0.017
R22844 GND.n1251 GND.n1250 0.017
R22845 GND.n1321 GND.n1320 0.017
R22846 GND.n1324 GND.n1323 0.017
R22847 GND.n1329 GND.n1328 0.017
R22848 GND.n1227 GND.n1226 0.017
R22849 GND.n1288 GND.n1287 0.017
R22850 GND.n1290 GND.n1289 0.017
R22851 GND.n1134 GND.n1133 0.017
R22852 GND.n1204 GND.n1203 0.017
R22853 GND.n1207 GND.n1206 0.017
R22854 GND.n1212 GND.n1211 0.017
R22855 GND.n1110 GND.n1109 0.017
R22856 GND.n1171 GND.n1170 0.017
R22857 GND.n1173 GND.n1172 0.017
R22858 GND.n1018 GND.n1017 0.017
R22859 GND.n1088 GND.n1087 0.017
R22860 GND.n1091 GND.n1090 0.017
R22861 GND.n1096 GND.n1095 0.017
R22862 GND.n994 GND.n993 0.017
R22863 GND.n1055 GND.n1054 0.017
R22864 GND.n1057 GND.n1056 0.017
R22865 GND.n618 GND.n608 0.017
R22866 GND.n742 GND.n740 0.017
R22867 GND.n306 GND.n305 0.017
R22868 GND.n282 GND.n281 0.017
R22869 GND.n280 GND.n279 0.017
R22870 GND.n483 GND.n482 0.017
R22871 GND.n513 GND.n500 0.017
R22872 GND.n554 GND.n553 0.017
R22873 GND.n339 GND.n338 0.017
R22874 GND.n359 GND.n358 0.017
R22875 GND.n389 GND.n388 0.017
R22876 GND.n423 GND.n422 0.017
R22877 GND.n439 GND.n438 0.017
R22878 GND.n2272 GND.n2271 0.017
R22879 GND.n2990 GND.n2989 0.017
R22880 GND.n2996 GND.n2995 0.017
R22881 GND.n2912 GND.n2911 0.017
R22882 GND.n2291 GND.n2289 0.017
R22883 GND.n2390 GND.n2388 0.017
R22884 GND.n347 GND.n341 0.016
R22885 GND.n391 GND.n386 0.016
R22886 GND.n435 GND.n429 0.016
R22887 GND.n2585 GND.n2584 0.016
R22888 GND.n2632 GND.n2627 0.016
R22889 GND.n2647 GND.n2637 0.016
R22890 GND.n2412 GND.n2399 0.016
R22891 GND.n2461 GND.n2456 0.016
R22892 GND.n2476 GND.n2466 0.016
R22893 GND.n152 GND.n151 0.015
R22894 GND.n149 GND.n148 0.015
R22895 GND.n229 GND.n224 0.015
R22896 GND.n124 GND.n123 0.015
R22897 GND.n784 GND.n783 0.015
R22898 GND.n781 GND.n780 0.015
R22899 GND.n861 GND.n856 0.015
R22900 GND.n756 GND.n755 0.015
R22901 GND.n36 GND.n35 0.015
R22902 GND.n33 GND.n32 0.015
R22903 GND.n113 GND.n108 0.015
R22904 GND.n8 GND.n7 0.015
R22905 GND.n902 GND.n901 0.015
R22906 GND.n899 GND.n898 0.015
R22907 GND.n979 GND.n974 0.015
R22908 GND.n874 GND.n873 0.015
R22909 GND.n2188 GND.n2187 0.015
R22910 GND.n2185 GND.n2184 0.015
R22911 GND.n2265 GND.n2260 0.015
R22912 GND.n2160 GND.n2159 0.015
R22913 GND.n2071 GND.n2070 0.015
R22914 GND.n2068 GND.n2067 0.015
R22915 GND.n2148 GND.n2143 0.015
R22916 GND.n2043 GND.n2042 0.015
R22917 GND.n1954 GND.n1953 0.015
R22918 GND.n1951 GND.n1950 0.015
R22919 GND.n2031 GND.n2026 0.015
R22920 GND.n1926 GND.n1925 0.015
R22921 GND.n1837 GND.n1836 0.015
R22922 GND.n1834 GND.n1833 0.015
R22923 GND.n1914 GND.n1909 0.015
R22924 GND.n1809 GND.n1808 0.015
R22925 GND.n1720 GND.n1719 0.015
R22926 GND.n1717 GND.n1716 0.015
R22927 GND.n1797 GND.n1792 0.015
R22928 GND.n1692 GND.n1691 0.015
R22929 GND.n1603 GND.n1602 0.015
R22930 GND.n1600 GND.n1599 0.015
R22931 GND.n1680 GND.n1675 0.015
R22932 GND.n1575 GND.n1574 0.015
R22933 GND.n1486 GND.n1485 0.015
R22934 GND.n1483 GND.n1482 0.015
R22935 GND.n1563 GND.n1558 0.015
R22936 GND.n1458 GND.n1457 0.015
R22937 GND.n1369 GND.n1368 0.015
R22938 GND.n1366 GND.n1365 0.015
R22939 GND.n1446 GND.n1441 0.015
R22940 GND.n1341 GND.n1340 0.015
R22941 GND.n1252 GND.n1251 0.015
R22942 GND.n1249 GND.n1248 0.015
R22943 GND.n1329 GND.n1324 0.015
R22944 GND.n1224 GND.n1223 0.015
R22945 GND.n1135 GND.n1134 0.015
R22946 GND.n1132 GND.n1131 0.015
R22947 GND.n1212 GND.n1207 0.015
R22948 GND.n1107 GND.n1106 0.015
R22949 GND.n1019 GND.n1018 0.015
R22950 GND.n1016 GND.n1015 0.015
R22951 GND.n1096 GND.n1091 0.015
R22952 GND.n991 GND.n990 0.015
R22953 GND.n608 GND.n606 0.015
R22954 GND.n744 GND.n742 0.015
R22955 GND.n328 GND.n327 0.015
R22956 GND.n311 GND.n310 0.015
R22957 GND.n281 GND.n280 0.015
R22958 GND.n455 GND.n454 0.015
R22959 GND.n500 GND.n499 0.015
R22960 GND.n514 GND.n513 0.015
R22961 GND.n538 GND.n537 0.015
R22962 GND.n570 GND.n569 0.015
R22963 GND.n334 GND.n333 0.015
R22964 GND.n354 GND.n351 0.015
R22965 GND.n376 GND.n375 0.015
R22966 GND.n379 GND.n378 0.015
R22967 GND.n413 GND.n412 0.015
R22968 GND.n419 GND.n418 0.015
R22969 GND.n433 GND.n432 0.015
R22970 GND.n2988 GND.n2987 0.015
R22971 GND.n2978 GND.n2977 0.015
R22972 GND.n2802 GND.n2801 0.015
R22973 GND.n2770 GND.n2761 0.015
R22974 GND.n2867 GND.n2866 0.015
R22975 GND.n2778 GND.n2777 0.015
R22976 GND.n2299 GND.n2291 0.015
R22977 GND.n2388 GND.n2386 0.015
R22978 GND.n244 GND.n243 0.014
R22979 GND.n2933 GND.n2932 0.014
R22980 GND.n2896 GND.n2895 0.014
R22981 GND.n2833 GND.n2832 0.014
R22982 GND.n2782 GND.n2781 0.014
R22983 GND.n2730 GND.n2729 0.014
R22984 GND.n2971 GND.n2946 0.013
R22985 GND.n162 GND.n158 0.013
R22986 GND.n207 GND.n206 0.013
R22987 GND.n218 GND.n217 0.013
R22988 GND.n186 GND.n185 0.013
R22989 GND.n794 GND.n790 0.013
R22990 GND.n839 GND.n838 0.013
R22991 GND.n850 GND.n849 0.013
R22992 GND.n818 GND.n817 0.013
R22993 GND.n46 GND.n42 0.013
R22994 GND.n91 GND.n90 0.013
R22995 GND.n102 GND.n101 0.013
R22996 GND.n70 GND.n69 0.013
R22997 GND.n912 GND.n908 0.013
R22998 GND.n957 GND.n956 0.013
R22999 GND.n968 GND.n967 0.013
R23000 GND.n936 GND.n935 0.013
R23001 GND.n2198 GND.n2194 0.013
R23002 GND.n2243 GND.n2242 0.013
R23003 GND.n2254 GND.n2253 0.013
R23004 GND.n2222 GND.n2221 0.013
R23005 GND.n2081 GND.n2077 0.013
R23006 GND.n2126 GND.n2125 0.013
R23007 GND.n2137 GND.n2136 0.013
R23008 GND.n2105 GND.n2104 0.013
R23009 GND.n1964 GND.n1960 0.013
R23010 GND.n2009 GND.n2008 0.013
R23011 GND.n2020 GND.n2019 0.013
R23012 GND.n1988 GND.n1987 0.013
R23013 GND.n1847 GND.n1843 0.013
R23014 GND.n1892 GND.n1891 0.013
R23015 GND.n1903 GND.n1902 0.013
R23016 GND.n1871 GND.n1870 0.013
R23017 GND.n1730 GND.n1726 0.013
R23018 GND.n1775 GND.n1774 0.013
R23019 GND.n1786 GND.n1785 0.013
R23020 GND.n1754 GND.n1753 0.013
R23021 GND.n1613 GND.n1609 0.013
R23022 GND.n1658 GND.n1657 0.013
R23023 GND.n1669 GND.n1668 0.013
R23024 GND.n1637 GND.n1636 0.013
R23025 GND.n1496 GND.n1492 0.013
R23026 GND.n1541 GND.n1540 0.013
R23027 GND.n1552 GND.n1551 0.013
R23028 GND.n1520 GND.n1519 0.013
R23029 GND.n1379 GND.n1375 0.013
R23030 GND.n1424 GND.n1423 0.013
R23031 GND.n1435 GND.n1434 0.013
R23032 GND.n1403 GND.n1402 0.013
R23033 GND.n1262 GND.n1258 0.013
R23034 GND.n1307 GND.n1306 0.013
R23035 GND.n1318 GND.n1317 0.013
R23036 GND.n1286 GND.n1285 0.013
R23037 GND.n1145 GND.n1141 0.013
R23038 GND.n1190 GND.n1189 0.013
R23039 GND.n1201 GND.n1200 0.013
R23040 GND.n1169 GND.n1168 0.013
R23041 GND.n1029 GND.n1025 0.013
R23042 GND.n1074 GND.n1073 0.013
R23043 GND.n1085 GND.n1084 0.013
R23044 GND.n1053 GND.n1052 0.013
R23045 GND.n632 GND.n622 0.013
R23046 GND.n728 GND.n726 0.013
R23047 GND.n329 GND.n328 0.013
R23048 GND.n308 GND.n307 0.013
R23049 GND.n468 GND.n457 0.013
R23050 GND.n498 GND.n497 0.013
R23051 GND.n533 GND.n520 0.013
R23052 GND.n551 GND.n539 0.013
R23053 GND.n571 GND.n570 0.013
R23054 GND.n361 GND.n360 0.013
R23055 GND.n370 GND.n369 0.013
R23056 GND.n398 GND.n395 0.013
R23057 GND.n397 GND.n396 0.013
R23058 GND.n2965 GND.n2964 0.013
R23059 GND.n2945 GND.n2944 0.013
R23060 GND.n2884 GND.n2883 0.013
R23061 GND.n2864 GND.n2863 0.013
R23062 GND.n2836 GND.n2835 0.013
R23063 GND.n2838 GND.n2837 0.013
R23064 GND.n2801 GND.n2800 0.013
R23065 GND.n2791 GND.n2790 0.013
R23066 GND.n2772 GND.n2771 0.013
R23067 GND.n2753 GND.n2752 0.013
R23068 GND.n2587 GND.n2586 0.013
R23069 GND.n2666 GND.n2650 0.013
R23070 GND.n2414 GND.n2413 0.013
R23071 GND.n2495 GND.n2479 0.013
R23072 GND.n239 GND.n237 0.013
R23073 GND.n2841 GND.n2840 0.012
R23074 GND.n2785 GND.n2784 0.012
R23075 GND.n171 GND.n170 0.012
R23076 GND.n172 GND.n171 0.012
R23077 GND.n803 GND.n802 0.012
R23078 GND.n804 GND.n803 0.012
R23079 GND.n55 GND.n54 0.012
R23080 GND.n56 GND.n55 0.012
R23081 GND.n921 GND.n920 0.012
R23082 GND.n922 GND.n921 0.012
R23083 GND.n2207 GND.n2206 0.012
R23084 GND.n2208 GND.n2207 0.012
R23085 GND.n2090 GND.n2089 0.012
R23086 GND.n2091 GND.n2090 0.012
R23087 GND.n1973 GND.n1972 0.012
R23088 GND.n1974 GND.n1973 0.012
R23089 GND.n1856 GND.n1855 0.012
R23090 GND.n1857 GND.n1856 0.012
R23091 GND.n1739 GND.n1738 0.012
R23092 GND.n1740 GND.n1739 0.012
R23093 GND.n1622 GND.n1621 0.012
R23094 GND.n1623 GND.n1622 0.012
R23095 GND.n1505 GND.n1504 0.012
R23096 GND.n1506 GND.n1505 0.012
R23097 GND.n1388 GND.n1387 0.012
R23098 GND.n1389 GND.n1388 0.012
R23099 GND.n1271 GND.n1270 0.012
R23100 GND.n1272 GND.n1271 0.012
R23101 GND.n1154 GND.n1153 0.012
R23102 GND.n1155 GND.n1154 0.012
R23103 GND.n1038 GND.n1037 0.012
R23104 GND.n1039 GND.n1038 0.012
R23105 GND.n2696 GND.n2560 0.012
R23106 GND.n232 GND.n231 0.012
R23107 GND.n864 GND.n863 0.012
R23108 GND.n116 GND.n115 0.012
R23109 GND.n982 GND.n981 0.012
R23110 GND.n2268 GND.n2267 0.012
R23111 GND.n2151 GND.n2150 0.012
R23112 GND.n2034 GND.n2033 0.012
R23113 GND.n1917 GND.n1916 0.012
R23114 GND.n1800 GND.n1799 0.012
R23115 GND.n1683 GND.n1682 0.012
R23116 GND.n1566 GND.n1565 0.012
R23117 GND.n1449 GND.n1448 0.012
R23118 GND.n1332 GND.n1331 0.012
R23119 GND.n1215 GND.n1214 0.012
R23120 GND.n1099 GND.n1098 0.012
R23121 GND.n747 GND.n746 0.012
R23122 GND.n150 GND.n149 0.011
R23123 GND.n208 GND.n207 0.011
R23124 GND.n168 GND.n167 0.011
R23125 GND.n175 GND.n174 0.011
R23126 GND.n782 GND.n781 0.011
R23127 GND.n840 GND.n839 0.011
R23128 GND.n800 GND.n799 0.011
R23129 GND.n807 GND.n806 0.011
R23130 GND.n34 GND.n33 0.011
R23131 GND.n92 GND.n91 0.011
R23132 GND.n52 GND.n51 0.011
R23133 GND.n59 GND.n58 0.011
R23134 GND.n900 GND.n899 0.011
R23135 GND.n958 GND.n957 0.011
R23136 GND.n918 GND.n917 0.011
R23137 GND.n925 GND.n924 0.011
R23138 GND.n2186 GND.n2185 0.011
R23139 GND.n2244 GND.n2243 0.011
R23140 GND.n2204 GND.n2203 0.011
R23141 GND.n2211 GND.n2210 0.011
R23142 GND.n2069 GND.n2068 0.011
R23143 GND.n2127 GND.n2126 0.011
R23144 GND.n2087 GND.n2086 0.011
R23145 GND.n2094 GND.n2093 0.011
R23146 GND.n1952 GND.n1951 0.011
R23147 GND.n2010 GND.n2009 0.011
R23148 GND.n1970 GND.n1969 0.011
R23149 GND.n1977 GND.n1976 0.011
R23150 GND.n1835 GND.n1834 0.011
R23151 GND.n1893 GND.n1892 0.011
R23152 GND.n1853 GND.n1852 0.011
R23153 GND.n1860 GND.n1859 0.011
R23154 GND.n1718 GND.n1717 0.011
R23155 GND.n1776 GND.n1775 0.011
R23156 GND.n1736 GND.n1735 0.011
R23157 GND.n1743 GND.n1742 0.011
R23158 GND.n1601 GND.n1600 0.011
R23159 GND.n1659 GND.n1658 0.011
R23160 GND.n1619 GND.n1618 0.011
R23161 GND.n1626 GND.n1625 0.011
R23162 GND.n1484 GND.n1483 0.011
R23163 GND.n1542 GND.n1541 0.011
R23164 GND.n1502 GND.n1501 0.011
R23165 GND.n1509 GND.n1508 0.011
R23166 GND.n1367 GND.n1366 0.011
R23167 GND.n1425 GND.n1424 0.011
R23168 GND.n1385 GND.n1384 0.011
R23169 GND.n1392 GND.n1391 0.011
R23170 GND.n1250 GND.n1249 0.011
R23171 GND.n1308 GND.n1307 0.011
R23172 GND.n1268 GND.n1267 0.011
R23173 GND.n1275 GND.n1274 0.011
R23174 GND.n1133 GND.n1132 0.011
R23175 GND.n1191 GND.n1190 0.011
R23176 GND.n1151 GND.n1150 0.011
R23177 GND.n1158 GND.n1157 0.011
R23178 GND.n1017 GND.n1016 0.011
R23179 GND.n1075 GND.n1074 0.011
R23180 GND.n1035 GND.n1034 0.011
R23181 GND.n1042 GND.n1041 0.011
R23182 GND.n301 GND.n288 0.011
R23183 GND.n288 GND.n287 0.011
R23184 GND.n495 GND.n494 0.011
R23185 GND.n520 GND.n519 0.011
R23186 GND.n395 GND.n394 0.011
R23187 GND.n404 GND.n403 0.011
R23188 GND.n2989 GND.n2988 0.011
R23189 GND.n2951 GND.n2949 0.011
R23190 GND.n2966 GND.n2965 0.011
R23191 GND.n2937 GND.n2936 0.011
R23192 GND.n2924 GND.n2923 0.011
R23193 GND.n2923 GND.n2922 0.011
R23194 GND.n2921 GND.n2920 0.011
R23195 GND.n2902 GND.n2901 0.011
R23196 GND.n2763 GND.n2762 0.011
R23197 GND.n2716 GND.n2715 0.011
R23198 GND.n2700 GND.n2699 0.011
R23199 GND.n2704 GND.n2700 0.011
R23200 GND.n2891 GND.n2890 0.011
R23201 GND.n2872 GND.n2871 0.011
R23202 GND.n2868 GND.n2865 0.011
R23203 GND.n2803 GND.n2794 0.011
R23204 GND.n2312 GND.n2303 0.011
R23205 GND.n2376 GND.n2374 0.011
R23206 GND.n3051 GND.n3050 0.011
R23207 GND.n3050 GND.n3049 0.011
R23208 GND.n3016 GND.n3014 0.011
R23209 GND.n3049 GND.n3047 0.01
R23210 GND.n3025 GND.n3024 0.01
R23211 GND.n3024 GND.n3016 0.01
R23212 GND.n3059 GND.n3056 0.009
R23213 GND.n3095 GND.n3092 0.009
R23214 GND.n240 GND.n239 0.009
R23215 GND.n241 GND.n240 0.009
R23216 GND.n200 GND.n199 0.009
R23217 GND.n181 GND.n180 0.009
R23218 GND.n832 GND.n831 0.009
R23219 GND.n813 GND.n812 0.009
R23220 GND.n84 GND.n83 0.009
R23221 GND.n65 GND.n64 0.009
R23222 GND.n950 GND.n949 0.009
R23223 GND.n931 GND.n930 0.009
R23224 GND.n2236 GND.n2235 0.009
R23225 GND.n2217 GND.n2216 0.009
R23226 GND.n2119 GND.n2118 0.009
R23227 GND.n2100 GND.n2099 0.009
R23228 GND.n2002 GND.n2001 0.009
R23229 GND.n1983 GND.n1982 0.009
R23230 GND.n1885 GND.n1884 0.009
R23231 GND.n1866 GND.n1865 0.009
R23232 GND.n1768 GND.n1767 0.009
R23233 GND.n1749 GND.n1748 0.009
R23234 GND.n1651 GND.n1650 0.009
R23235 GND.n1632 GND.n1631 0.009
R23236 GND.n1534 GND.n1533 0.009
R23237 GND.n1515 GND.n1514 0.009
R23238 GND.n1417 GND.n1416 0.009
R23239 GND.n1398 GND.n1397 0.009
R23240 GND.n1300 GND.n1299 0.009
R23241 GND.n1281 GND.n1280 0.009
R23242 GND.n1183 GND.n1182 0.009
R23243 GND.n1164 GND.n1163 0.009
R23244 GND.n1067 GND.n1066 0.009
R23245 GND.n1048 GND.n1047 0.009
R23246 GND.n646 GND.n636 0.009
R23247 GND.n714 GND.n712 0.009
R23248 GND.n315 GND.n314 0.009
R23249 GND.n310 GND.n309 0.009
R23250 GND.n287 GND.n286 0.009
R23251 GND.n553 GND.n552 0.009
R23252 GND.n557 GND.n556 0.009
R23253 GND.n572 GND.n571 0.009
R23254 GND.n335 GND.n334 0.009
R23255 GND.n351 GND.n350 0.009
R23256 GND.n364 GND.n361 0.009
R23257 GND.n371 GND.n370 0.009
R23258 GND.n378 GND.n377 0.009
R23259 GND.n407 GND.n404 0.009
R23260 GND.n414 GND.n413 0.009
R23261 GND.n434 GND.n433 0.009
R23262 GND.n357 GND.n356 0.009
R23263 GND.n374 GND.n373 0.009
R23264 GND.n401 GND.n400 0.009
R23265 GND.n417 GND.n416 0.009
R23266 GND.n2272 GND.n985 0.009
R23267 GND.n2957 GND.n2956 0.009
R23268 GND.n2940 GND.n2939 0.009
R23269 GND.n2982 GND.n2981 0.009
R23270 GND.n2976 GND.n2975 0.009
R23271 GND.n2975 GND.n2974 0.009
R23272 GND.n2930 GND.n2925 0.009
R23273 GND.n2929 GND.n2928 0.009
R23274 GND.n2914 GND.n2913 0.009
R23275 GND.n2754 GND.n2750 0.009
R23276 GND.n2727 GND.n2710 0.009
R23277 GND.n2707 GND.n2706 0.009
R23278 GND.n2626 GND.n2625 0.009
R23279 GND.n2441 GND.n2440 0.009
R23280 GND.n2455 GND.n2454 0.009
R23281 GND.n2894 GND.n2875 0.008
R23282 GND.n2874 GND.n2873 0.008
R23283 GND.n2869 GND.n2850 0.008
R23284 GND.n2849 GND.n2848 0.008
R23285 GND.n2780 GND.n2775 0.008
R23286 GND.n2774 GND.n2773 0.008
R23287 GND.n2755 GND.n2749 0.008
R23288 GND.n2748 GND.n2747 0.008
R23289 GND.n3060 GND.n3055 0.008
R23290 GND.n3096 GND.n3091 0.008
R23291 GND.n142 GND.n141 0.007
R23292 GND.n202 GND.n201 0.007
R23293 GND.n121 GND.n120 0.007
R23294 GND.n183 GND.n182 0.007
R23295 GND.n774 GND.n773 0.007
R23296 GND.n834 GND.n833 0.007
R23297 GND.n753 GND.n752 0.007
R23298 GND.n815 GND.n814 0.007
R23299 GND.n26 GND.n25 0.007
R23300 GND.n86 GND.n85 0.007
R23301 GND.n5 GND.n4 0.007
R23302 GND.n67 GND.n66 0.007
R23303 GND.n892 GND.n891 0.007
R23304 GND.n952 GND.n951 0.007
R23305 GND.n871 GND.n870 0.007
R23306 GND.n933 GND.n932 0.007
R23307 GND.n2178 GND.n2177 0.007
R23308 GND.n2238 GND.n2237 0.007
R23309 GND.n2157 GND.n2156 0.007
R23310 GND.n2219 GND.n2218 0.007
R23311 GND.n2061 GND.n2060 0.007
R23312 GND.n2121 GND.n2120 0.007
R23313 GND.n2040 GND.n2039 0.007
R23314 GND.n2102 GND.n2101 0.007
R23315 GND.n1944 GND.n1943 0.007
R23316 GND.n2004 GND.n2003 0.007
R23317 GND.n1923 GND.n1922 0.007
R23318 GND.n1985 GND.n1984 0.007
R23319 GND.n1827 GND.n1826 0.007
R23320 GND.n1887 GND.n1886 0.007
R23321 GND.n1806 GND.n1805 0.007
R23322 GND.n1868 GND.n1867 0.007
R23323 GND.n1710 GND.n1709 0.007
R23324 GND.n1770 GND.n1769 0.007
R23325 GND.n1689 GND.n1688 0.007
R23326 GND.n1751 GND.n1750 0.007
R23327 GND.n1593 GND.n1592 0.007
R23328 GND.n1653 GND.n1652 0.007
R23329 GND.n1572 GND.n1571 0.007
R23330 GND.n1634 GND.n1633 0.007
R23331 GND.n1476 GND.n1475 0.007
R23332 GND.n1536 GND.n1535 0.007
R23333 GND.n1455 GND.n1454 0.007
R23334 GND.n1517 GND.n1516 0.007
R23335 GND.n1359 GND.n1358 0.007
R23336 GND.n1419 GND.n1418 0.007
R23337 GND.n1338 GND.n1337 0.007
R23338 GND.n1400 GND.n1399 0.007
R23339 GND.n1242 GND.n1241 0.007
R23340 GND.n1302 GND.n1301 0.007
R23341 GND.n1221 GND.n1220 0.007
R23342 GND.n1283 GND.n1282 0.007
R23343 GND.n1125 GND.n1124 0.007
R23344 GND.n1185 GND.n1184 0.007
R23345 GND.n1104 GND.n1103 0.007
R23346 GND.n1166 GND.n1165 0.007
R23347 GND.n1009 GND.n1008 0.007
R23348 GND.n1069 GND.n1068 0.007
R23349 GND.n988 GND.n987 0.007
R23350 GND.n1050 GND.n1049 0.007
R23351 GND.n330 GND.n329 0.007
R23352 GND.n327 GND.n315 0.007
R23353 GND.n307 GND.n306 0.007
R23354 GND.n482 GND.n477 0.007
R23355 GND.n519 GND.n518 0.007
R23356 GND.n539 GND.n538 0.007
R23357 GND.n569 GND.n557 0.007
R23358 GND.n340 GND.n339 0.007
R23359 GND.n343 GND.n342 0.007
R23360 GND.n390 GND.n389 0.007
R23361 GND.n422 GND.n421 0.007
R23362 GND.n431 GND.n430 0.007
R23363 GND.n575 GND.n439 0.007
R23364 GND.n2948 GND.n2947 0.007
R23365 GND.n2959 GND.n2958 0.007
R23366 GND.n2935 GND.n2934 0.007
R23367 GND.n2942 GND.n2941 0.007
R23368 GND.n2816 GND.n2815 0.007
R23369 GND.n2805 GND.n2804 0.007
R23370 GND.n2324 GND.n2316 0.007
R23371 GND.n2363 GND.n2361 0.007
R23372 GND.n2610 GND.n2604 0.007
R23373 GND.n2622 GND.n2615 0.007
R23374 GND.n2648 GND.n2633 0.007
R23375 GND.n2437 GND.n2431 0.007
R23376 GND.n2451 GND.n2444 0.007
R23377 GND.n2477 GND.n2462 0.007
R23378 GND.n3064 GND.n3063 0.007
R23379 GND.n3124 GND.n3100 0.007
R23380 GND.n2585 GND.n2582 0.007
R23381 GND.n2412 GND.n2411 0.007
R23382 GND.n2665 GND.n2664 0.006
R23383 GND.n2494 GND.n2493 0.006
R23384 GND.n167 GND.n166 0.006
R23385 GND.n169 GND.n168 0.006
R23386 GND.n174 GND.n173 0.006
R23387 GND.n176 GND.n175 0.006
R23388 GND.n799 GND.n798 0.006
R23389 GND.n801 GND.n800 0.006
R23390 GND.n806 GND.n805 0.006
R23391 GND.n808 GND.n807 0.006
R23392 GND.n51 GND.n50 0.006
R23393 GND.n53 GND.n52 0.006
R23394 GND.n58 GND.n57 0.006
R23395 GND.n60 GND.n59 0.006
R23396 GND.n917 GND.n916 0.006
R23397 GND.n919 GND.n918 0.006
R23398 GND.n924 GND.n923 0.006
R23399 GND.n926 GND.n925 0.006
R23400 GND.n2203 GND.n2202 0.006
R23401 GND.n2205 GND.n2204 0.006
R23402 GND.n2210 GND.n2209 0.006
R23403 GND.n2212 GND.n2211 0.006
R23404 GND.n2086 GND.n2085 0.006
R23405 GND.n2088 GND.n2087 0.006
R23406 GND.n2093 GND.n2092 0.006
R23407 GND.n2095 GND.n2094 0.006
R23408 GND.n1969 GND.n1968 0.006
R23409 GND.n1971 GND.n1970 0.006
R23410 GND.n1976 GND.n1975 0.006
R23411 GND.n1978 GND.n1977 0.006
R23412 GND.n1852 GND.n1851 0.006
R23413 GND.n1854 GND.n1853 0.006
R23414 GND.n1859 GND.n1858 0.006
R23415 GND.n1861 GND.n1860 0.006
R23416 GND.n1735 GND.n1734 0.006
R23417 GND.n1737 GND.n1736 0.006
R23418 GND.n1742 GND.n1741 0.006
R23419 GND.n1744 GND.n1743 0.006
R23420 GND.n1618 GND.n1617 0.006
R23421 GND.n1620 GND.n1619 0.006
R23422 GND.n1625 GND.n1624 0.006
R23423 GND.n1627 GND.n1626 0.006
R23424 GND.n1501 GND.n1500 0.006
R23425 GND.n1503 GND.n1502 0.006
R23426 GND.n1508 GND.n1507 0.006
R23427 GND.n1510 GND.n1509 0.006
R23428 GND.n1384 GND.n1383 0.006
R23429 GND.n1386 GND.n1385 0.006
R23430 GND.n1391 GND.n1390 0.006
R23431 GND.n1393 GND.n1392 0.006
R23432 GND.n1267 GND.n1266 0.006
R23433 GND.n1269 GND.n1268 0.006
R23434 GND.n1274 GND.n1273 0.006
R23435 GND.n1276 GND.n1275 0.006
R23436 GND.n1150 GND.n1149 0.006
R23437 GND.n1152 GND.n1151 0.006
R23438 GND.n1157 GND.n1156 0.006
R23439 GND.n1159 GND.n1158 0.006
R23440 GND.n1034 GND.n1033 0.006
R23441 GND.n1036 GND.n1035 0.006
R23442 GND.n1041 GND.n1040 0.006
R23443 GND.n1043 GND.n1042 0.006
R23444 GND.n2907 GND.n2902 0.006
R23445 GND.n2888 GND.n2887 0.006
R23446 GND.n2887 GND.n2886 0.006
R23447 GND.n2852 GND.n2851 0.006
R23448 GND.n2765 GND.n2764 0.006
R23449 GND.n2736 GND.n2735 0.006
R23450 GND.n2744 GND.n2736 0.006
R23451 GND.n2742 GND.n2741 0.006
R23452 GND.n2725 GND.n2716 0.006
R23453 GND.n2611 GND.n2610 0.006
R23454 GND.n2615 GND.n2611 0.006
R23455 GND.n2633 GND.n2624 0.006
R23456 GND.n2438 GND.n2437 0.006
R23457 GND.n2444 GND.n2439 0.006
R23458 GND.n2452 GND.n2451 0.006
R23459 GND.n2462 GND.n2453 0.006
R23460 GND.n3000 GND.n2696 0.006
R23461 GND.n3026 GND.n3000 0.006
R23462 GND.n3126 GND.n3125 0.006
R23463 GND.n660 GND.n650 0.005
R23464 GND.n700 GND.n698 0.005
R23465 GND.n303 GND.n302 0.005
R23466 GND.n283 GND.n282 0.005
R23467 GND.n470 GND.n469 0.005
R23468 GND.n475 GND.n474 0.005
R23469 GND.n484 GND.n483 0.005
R23470 GND.n515 GND.n514 0.005
R23471 GND.n535 GND.n534 0.005
R23472 GND.n385 GND.n384 0.005
R23473 GND.n341 GND.n337 0.005
R23474 GND.n348 GND.n347 0.005
R23475 GND.n355 GND.n349 0.005
R23476 GND.n381 GND.n380 0.005
R23477 GND.n386 GND.n382 0.005
R23478 GND.n392 GND.n391 0.005
R23479 GND.n399 GND.n393 0.005
R23480 GND.n425 GND.n424 0.005
R23481 GND.n429 GND.n426 0.005
R23482 GND.n436 GND.n435 0.005
R23483 GND.n576 GND.n437 0.005
R23484 GND.n2997 GND.n2982 0.005
R23485 GND.n2981 GND.n2980 0.005
R23486 GND.n2973 GND.n2972 0.005
R23487 GND.n2914 GND.n2908 0.005
R23488 GND.n2893 GND.n2889 0.005
R23489 GND.n2820 GND.n2819 0.005
R23490 GND.n2746 GND.n2745 0.005
R23491 GND.n2733 GND.n2732 0.005
R23492 GND.n2727 GND.n2726 0.005
R23493 GND.n2875 GND.n2874 0.005
R23494 GND.n2850 GND.n2849 0.005
R23495 GND.n2775 GND.n2774 0.005
R23496 GND.n2749 GND.n2748 0.005
R23497 GND.n2604 GND.n2588 0.005
R23498 GND.n2623 GND.n2622 0.005
R23499 GND.n2431 GND.n2415 0.005
R23500 GND.n2478 GND.n2477 0.005
R23501 GND.n3059 GND.n3058 0.005
R23502 GND.n3095 GND.n3094 0.005
R23503 GND.n2924 GND.n2919 0.005
R23504 GND.n2704 GND.n2703 0.005
R23505 GND.n2993 GND.n2990 0.005
R23506 GND.n3062 GND.n3061 0.004
R23507 GND.n3090 GND.n3089 0.004
R23508 GND.n3088 GND.n3062 0.004
R23509 GND.n3089 GND.n3088 0.004
R23510 GND.n3099 GND.n3098 0.004
R23511 GND.n3098 GND.n3097 0.004
R23512 GND.n2970 GND.n2967 0.004
R23513 GND.n2898 GND.n2897 0.004
R23514 GND.n2877 GND.n2876 0.004
R23515 GND.n2858 GND.n2857 0.004
R23516 GND.n2843 GND.n2836 0.004
R23517 GND.n2828 GND.n2827 0.004
R23518 GND.n2682 GND.n2677 0.004
R23519 GND.n2692 GND.n2690 0.004
R23520 GND.n2586 GND.n2570 0.004
R23521 GND.n2649 GND.n2648 0.004
R23522 GND.n2413 GND.n2397 0.004
R23523 GND.n2531 GND.n2521 0.004
R23524 GND.n2547 GND.n2545 0.004
R23525 GND.n3102 GND.n3101 0.004
R23526 GND.n3125 GND.n3099 0.003
R23527 GND.n3087 GND.n3086 0.003
R23528 GND.n153 GND.n152 0.003
R23529 GND.n206 GND.n203 0.003
R23530 GND.n219 GND.n218 0.003
R23531 GND.n185 GND.n184 0.003
R23532 GND.n785 GND.n784 0.003
R23533 GND.n838 GND.n835 0.003
R23534 GND.n851 GND.n850 0.003
R23535 GND.n817 GND.n816 0.003
R23536 GND.n37 GND.n36 0.003
R23537 GND.n90 GND.n87 0.003
R23538 GND.n103 GND.n102 0.003
R23539 GND.n69 GND.n68 0.003
R23540 GND.n903 GND.n902 0.003
R23541 GND.n956 GND.n953 0.003
R23542 GND.n969 GND.n968 0.003
R23543 GND.n935 GND.n934 0.003
R23544 GND.n2189 GND.n2188 0.003
R23545 GND.n2242 GND.n2239 0.003
R23546 GND.n2255 GND.n2254 0.003
R23547 GND.n2221 GND.n2220 0.003
R23548 GND.n2072 GND.n2071 0.003
R23549 GND.n2125 GND.n2122 0.003
R23550 GND.n2138 GND.n2137 0.003
R23551 GND.n2104 GND.n2103 0.003
R23552 GND.n1955 GND.n1954 0.003
R23553 GND.n2008 GND.n2005 0.003
R23554 GND.n2021 GND.n2020 0.003
R23555 GND.n1987 GND.n1986 0.003
R23556 GND.n1838 GND.n1837 0.003
R23557 GND.n1891 GND.n1888 0.003
R23558 GND.n1904 GND.n1903 0.003
R23559 GND.n1870 GND.n1869 0.003
R23560 GND.n1721 GND.n1720 0.003
R23561 GND.n1774 GND.n1771 0.003
R23562 GND.n1787 GND.n1786 0.003
R23563 GND.n1753 GND.n1752 0.003
R23564 GND.n1604 GND.n1603 0.003
R23565 GND.n1657 GND.n1654 0.003
R23566 GND.n1670 GND.n1669 0.003
R23567 GND.n1636 GND.n1635 0.003
R23568 GND.n1487 GND.n1486 0.003
R23569 GND.n1540 GND.n1537 0.003
R23570 GND.n1553 GND.n1552 0.003
R23571 GND.n1519 GND.n1518 0.003
R23572 GND.n1370 GND.n1369 0.003
R23573 GND.n1423 GND.n1420 0.003
R23574 GND.n1436 GND.n1435 0.003
R23575 GND.n1402 GND.n1401 0.003
R23576 GND.n1253 GND.n1252 0.003
R23577 GND.n1306 GND.n1303 0.003
R23578 GND.n1319 GND.n1318 0.003
R23579 GND.n1285 GND.n1284 0.003
R23580 GND.n1136 GND.n1135 0.003
R23581 GND.n1189 GND.n1186 0.003
R23582 GND.n1202 GND.n1201 0.003
R23583 GND.n1168 GND.n1167 0.003
R23584 GND.n1020 GND.n1019 0.003
R23585 GND.n1073 GND.n1070 0.003
R23586 GND.n1086 GND.n1085 0.003
R23587 GND.n1052 GND.n1051 0.003
R23588 GND.n337 GND.n336 0.003
R23589 GND.n349 GND.n348 0.003
R23590 GND.n382 GND.n381 0.003
R23591 GND.n393 GND.n392 0.003
R23592 GND.n426 GND.n425 0.003
R23593 GND.n437 GND.n436 0.003
R23594 GND.n2964 GND.n2960 0.003
R23595 GND.n2944 GND.n2943 0.003
R23596 GND.n2927 GND.n2926 0.003
R23597 GND.n2910 GND.n2909 0.003
R23598 GND.n2892 GND.n2891 0.003
R23599 GND.n2847 GND.n2846 0.003
R23600 GND.n2845 GND.n2844 0.003
R23601 GND.n2829 GND.n2821 0.003
R23602 GND.n2932 GND.n2931 0.003
R23603 GND.n2915 GND.n2896 0.003
R23604 GND.n2832 GND.n2831 0.003
R23605 GND.n2807 GND.n2782 0.003
R23606 GND.n2729 GND.n2728 0.003
R23607 GND.n2337 GND.n2328 0.003
R23608 GND.n2351 GND.n2349 0.003
R23609 GND.n2650 GND.n2649 0.003
R23610 GND.n2667 GND.n2666 0.003
R23611 GND.n2479 GND.n2478 0.003
R23612 GND.n2496 GND.n2495 0.003
R23613 GND.n365 GND.n357 0.002
R23614 GND.n373 GND.n372 0.002
R23615 GND.n408 GND.n401 0.002
R23616 GND.n416 GND.n415 0.002
R23617 GND.n2863 GND.n2862 0.002
R23618 GND.n2812 GND.n2811 0.002
R23619 GND.n2796 GND.n2795 0.002
R23620 GND.n2792 GND.n2791 0.002
R23621 GND.n2789 GND.n2788 0.002
R23622 GND.n2761 GND.n2760 0.002
R23623 GND.n2723 GND.n2722 0.002
R23624 GND.n2588 GND.n2587 0.002
R23625 GND.n2415 GND.n2414 0.002
R23626 GND.n3066 GND.n3064 0.002
R23627 GND.n3086 GND.n3085 0.002
R23628 GND.n3124 GND.n3123 0.002
R23629 GND.n3104 GND.n3102 0.002
R23630 GND.n148 GND.n143 0.001
R23631 GND.n126 GND.n125 0.001
R23632 GND.n123 GND.n122 0.001
R23633 GND.n780 GND.n775 0.001
R23634 GND.n758 GND.n757 0.001
R23635 GND.n755 GND.n754 0.001
R23636 GND.n32 GND.n27 0.001
R23637 GND.n10 GND.n9 0.001
R23638 GND.n7 GND.n6 0.001
R23639 GND.n898 GND.n893 0.001
R23640 GND.n876 GND.n875 0.001
R23641 GND.n873 GND.n872 0.001
R23642 GND.n2184 GND.n2179 0.001
R23643 GND.n2162 GND.n2161 0.001
R23644 GND.n2159 GND.n2158 0.001
R23645 GND.n2067 GND.n2062 0.001
R23646 GND.n2045 GND.n2044 0.001
R23647 GND.n2042 GND.n2041 0.001
R23648 GND.n1950 GND.n1945 0.001
R23649 GND.n1928 GND.n1927 0.001
R23650 GND.n1925 GND.n1924 0.001
R23651 GND.n1833 GND.n1828 0.001
R23652 GND.n1811 GND.n1810 0.001
R23653 GND.n1808 GND.n1807 0.001
R23654 GND.n1716 GND.n1711 0.001
R23655 GND.n1694 GND.n1693 0.001
R23656 GND.n1691 GND.n1690 0.001
R23657 GND.n1599 GND.n1594 0.001
R23658 GND.n1577 GND.n1576 0.001
R23659 GND.n1574 GND.n1573 0.001
R23660 GND.n1482 GND.n1477 0.001
R23661 GND.n1460 GND.n1459 0.001
R23662 GND.n1457 GND.n1456 0.001
R23663 GND.n1365 GND.n1360 0.001
R23664 GND.n1343 GND.n1342 0.001
R23665 GND.n1340 GND.n1339 0.001
R23666 GND.n1248 GND.n1243 0.001
R23667 GND.n1226 GND.n1225 0.001
R23668 GND.n1223 GND.n1222 0.001
R23669 GND.n1131 GND.n1126 0.001
R23670 GND.n1109 GND.n1108 0.001
R23671 GND.n1106 GND.n1105 0.001
R23672 GND.n1015 GND.n1010 0.001
R23673 GND.n993 GND.n992 0.001
R23674 GND.n990 GND.n989 0.001
R23675 GND.n674 GND.n664 0.001
R23676 GND.n686 GND.n684 0.001
R23677 GND.n313 GND.n312 0.001
R23678 GND.n457 GND.n456 0.001
R23679 GND.n496 GND.n495 0.001
R23680 GND.n346 GND.n345 0.001
R23681 GND.n749 GND.n748 0.001
R23682 GND.n748 GND.n577 0.001
R23683 GND.n2987 GND.n2983 0.001
R23684 GND.n2995 GND.n2994 0.001
R23685 GND.n2979 GND.n2978 0.001
R23686 GND.n2830 GND.n2816 0.001
R23687 GND.n2806 GND.n2805 0.001
R23688 GND.n2793 GND.n2783 0.001
R23689 GND.n2779 GND.n2776 0.001
R23690 GND.n2752 GND.n2751 0.001
R23691 GND.n2713 GND.n2712 0.001
R23692 GND.n2624 GND.n2623 0.001
R23693 GND.n2439 GND.n2438 0.001
R23694 GND.n2453 GND.n2452 0.001
R23695 VBP.n3 VBP.t13 308.184
R23696 VBP.n13 VBP.t18 308.184
R23697 VBP.n16 VBP.t16 307.987
R23698 VBP.n15 VBP.t11 307.987
R23699 VBP.n14 VBP.t17 307.987
R23700 VBP.n13 VBP.t10 307.987
R23701 VBP.n4 VBP.t14 307.987
R23702 VBP.n6 VBP.t15 307.987
R23703 VBP.n17 VBP.t9 307.986
R23704 VBP.n3 VBP.t6 307.986
R23705 VBP.n5 VBP.t8 307.986
R23706 VBP.n7 VBP.t7 307.986
R23707 VBP.n24 VBP.t5 248.432
R23708 VBP.n24 VBP.t12 248.427
R23709 VBP.n94 VBP.n93 175.251
R23710 VBP.n295 VBP.n294 175.251
R23711 VBP.n156 VBP.n155 175.251
R23712 VBP.n93 VBP.t0 131.474
R23713 VBP.n294 VBP.t4 131.474
R23714 VBP.n155 VBP.t3 131.474
R23715 VBP.n54 VBP.t2 124.695
R23716 VBP.n34 VBP.t1 124.695
R23717 VBP.n53 VBP.n52 92.5
R23718 VBP.n33 VBP.n32 92.5
R23719 VBP.n63 VBP.n62 31.034
R23720 VBP.n43 VBP.n42 31.034
R23721 VBP.n54 VBP.n53 15.431
R23722 VBP.n34 VBP.n33 15.431
R23723 VBP.n192 VBP.n191 9.3
R23724 VBP.n69 VBP.n68 9.3
R23725 VBP.n58 VBP.n57 9.3
R23726 VBP.n56 VBP.n55 9.3
R23727 VBP.n65 VBP.n64 9.3
R23728 VBP.n64 VBP.n63 9.3
R23729 VBP.n67 VBP.n66 9.3
R23730 VBP.n71 VBP.n70 9.3
R23731 VBP.n47 VBP.n46 9.3
R23732 VBP.n38 VBP.n37 9.3
R23733 VBP.n36 VBP.n35 9.3
R23734 VBP.n45 VBP.n44 9.3
R23735 VBP.n44 VBP.n43 9.3
R23736 VBP.n49 VBP.n48 9.3
R23737 VBP.n51 VBP.n50 9.3
R23738 VBP.n77 VBP.n76 9.013
R23739 VBP.n256 VBP.n255 9.013
R23740 VBP.n344 VBP.n343 9.013
R23741 VBP.n329 VBP.n328 9.013
R23742 VBP.n151 VBP.n150 9.013
R23743 VBP.n223 VBP.n222 9.013
R23744 VBP.n95 VBP.n94 6.413
R23745 VBP.n296 VBP.n295 6.413
R23746 VBP.n157 VBP.n156 6.413
R23747 VBP.n64 VBP.n60 5.647
R23748 VBP.n44 VBP.n40 5.647
R23749 VBP.n383 VBP.n31 4.699
R23750 VBP.n72 VBP.n51 4.659
R23751 VBP.n72 VBP.n71 4.647
R23752 VBP.n160 VBP.n159 4.5
R23753 VBP.n177 VBP.n176 4.5
R23754 VBP.n168 VBP.n167 4.5
R23755 VBP.n173 VBP.n172 4.5
R23756 VBP.n184 VBP.n183 4.5
R23757 VBP.n98 VBP.n97 4.5
R23758 VBP.n376 VBP.n373 4.5
R23759 VBP.n108 VBP.n107 4.5
R23760 VBP.n126 VBP.n124 4.5
R23761 VBP.n369 VBP.n366 4.5
R23762 VBP.n359 VBP.n356 4.5
R23763 VBP.n299 VBP.n298 4.5
R23764 VBP.n281 VBP.n263 4.5
R23765 VBP.n286 VBP.n259 4.5
R23766 VBP.n283 VBP.n261 4.5
R23767 VBP.n278 VBP.n266 4.5
R23768 VBP.n273 VBP.n270 4.5
R23769 VBP.n195 VBP.n194 4.5
R23770 VBP.n62 VBP.n61 4.137
R23771 VBP.n42 VBP.n41 4.137
R23772 VBP.n345 VBP.n344 3.992
R23773 VBP.n330 VBP.n329 3.992
R23774 VBP.n78 VBP.n77 3.882
R23775 VBP.n224 VBP.n223 3.882
R23776 VBP.n95 VBP.n91 3
R23777 VBP.n296 VBP.n292 3
R23778 VBP.n192 VBP.n190 3
R23779 VBP.n382 VBP.n381 2.844
R23780 VBP.n199 VBP.n151 2.797
R23781 VBP.n94 VBP.n92 2.787
R23782 VBP.n295 VBP.n293 2.787
R23783 VBP.n303 VBP.n256 2.742
R23784 VBP.n124 VBP.n123 2.656
R23785 VBP.n149 VBP.n148 2.535
R23786 VBP.n254 VBP.n253 2.415
R23787 VBP.n106 VBP.n105 2.26
R23788 VBP.n365 VBP.n364 2.26
R23789 VBP.n96 VBP.n95 2.26
R23790 VBP.n355 VBP.n354 2.26
R23791 VBP.n258 VBP.n257 2.26
R23792 VBP.n265 VBP.n264 2.26
R23793 VBP.n297 VBP.n296 2.26
R23794 VBP.n269 VBP.n268 2.26
R23795 VBP.n158 VBP.n157 2.26
R23796 VBP.n166 VBP.n165 2.26
R23797 VBP.n182 VBP.n181 2.26
R23798 VBP.n193 VBP.n192 2.26
R23799 VBP.n12 VBP.n10 2.25
R23800 VBP.n12 VBP.n11 2.25
R23801 VBP.n383 VBP.n382 1.851
R23802 VBP.n26 VBP.n25 1.705
R23803 VBP.n56 VBP.n54 1.57
R23804 VBP.n36 VBP.n34 1.57
R23805 VBP.n127 VBP.n126 1.501
R23806 VBP.n228 VBP.n227 1.5
R23807 VBP.n377 VBP.n376 1.5
R23808 VBP.n109 VBP.n108 1.5
R23809 VBP.n370 VBP.n369 1.5
R23810 VBP.n99 VBP.n98 1.5
R23811 VBP.n360 VBP.n359 1.5
R23812 VBP.n347 VBP.n346 1.5
R23813 VBP.n82 VBP.n81 1.5
R23814 VBP.n332 VBP.n331 1.5
R23815 VBP.n96 VBP.n90 1.449
R23816 VBP.n297 VBP.n291 1.449
R23817 VBP.n158 VBP.n154 1.449
R23818 VBP VBP.n23 1.378
R23819 VBP.n77 VBP.n75 1.328
R23820 VBP.n355 VBP.n353 1.328
R23821 VBP.n256 VBP.n254 1.328
R23822 VBP.n269 VBP.n267 1.328
R23823 VBP.n223 VBP.n221 1.328
R23824 VBP.n193 VBP.n189 1.328
R23825 VBP.n25 VBP.n24 1.208
R23826 VBP.n124 VBP.n112 1.207
R23827 VBP.n366 VBP.n365 1.207
R23828 VBP.n344 VBP.n342 1.207
R23829 VBP.n261 VBP.n260 1.207
R23830 VBP.n266 VBP.n265 1.207
R23831 VBP.n329 VBP.n327 1.207
R23832 VBP.n172 VBP.n171 1.207
R23833 VBP.n183 VBP.n182 1.207
R23834 VBP.n151 VBP.n149 1.207
R23835 VBP.n382 VBP.n72 1.163
R23836 VBP.n22 VBP.n21 1.135
R23837 VBP.n107 VBP.n106 1.086
R23838 VBP.n373 VBP.n372 1.086
R23839 VBP.n259 VBP.n258 1.086
R23840 VBP.n263 VBP.n262 1.086
R23841 VBP.n167 VBP.n166 1.086
R23842 VBP.n176 VBP.n175 1.086
R23843 VBP VBP.n383 1.086
R23844 VBP.n60 VBP.n59 0.752
R23845 VBP.n40 VBP.n39 0.752
R23846 VBP.n356 VBP.n355 0.724
R23847 VBP.n270 VBP.n269 0.724
R23848 VBP.n194 VBP.n193 0.724
R23849 VBP.n304 VBP.n303 0.722
R23850 VBP.n200 VBP.n199 0.722
R23851 VBP.n181 VBP.n180 0.604
R23852 VBP.n97 VBP.n96 0.603
R23853 VBP.n298 VBP.n297 0.603
R23854 VBP.n159 VBP.n158 0.603
R23855 VBP.n30 VBP.n28 0.476
R23856 VBP.n4 VBP.n3 0.197
R23857 VBP.n5 VBP.n4 0.197
R23858 VBP.n6 VBP.n5 0.197
R23859 VBP.n17 VBP.n16 0.197
R23860 VBP.n16 VBP.n15 0.197
R23861 VBP.n15 VBP.n14 0.197
R23862 VBP.n14 VBP.n13 0.197
R23863 VBP.n7 VBP.n6 0.196
R23864 VBP.n18 VBP.n17 0.188
R23865 VBP.n8 VBP.n7 0.184
R23866 VBP.n67 VBP.n65 0.144
R23867 VBP.n47 VBP.n45 0.144
R23868 VBP.n231 VBP.n230 0.129
R23869 VBP.n335 VBP.n334 0.128
R23870 VBP.n335 VBP.n242 0.05
R23871 VBP.n231 VBP.n138 0.05
R23872 VBP.n302 VBP.n301 0.048
R23873 VBP.n289 VBP.n288 0.048
R23874 VBP.n276 VBP.n275 0.048
R23875 VBP.n163 VBP.n162 0.048
R23876 VBP.n187 VBP.n186 0.048
R23877 VBP.n198 VBP.n197 0.048
R23878 VBP.n282 VBP.n281 0.044
R23879 VBP.n177 VBP.n174 0.044
R23880 VBP.n126 VBP.n125 0.042
R23881 VBP.n283 VBP.n282 0.042
R23882 VBP.n174 VBP.n173 0.042
R23883 VBP.n65 VBP.n58 0.04
R23884 VBP.n45 VBP.n38 0.04
R23885 VBP.n108 VBP.n104 0.036
R23886 VBP.n287 VBP.n286 0.036
R23887 VBP.n168 VBP.n164 0.036
R23888 VBP.n71 VBP.n69 0.035
R23889 VBP.n51 VBP.n49 0.035
R23890 VBP.n28 VBP.n26 0.034
R23891 VBP.n369 VBP.n368 0.034
R23892 VBP.n278 VBP.n277 0.034
R23893 VBP.n185 VBP.n184 0.034
R23894 VBP.n379 VBP.n335 0.033
R23895 VBP.n379 VBP.n231 0.032
R23896 VBP.n303 VBP.n302 0.028
R23897 VBP.n98 VBP.n87 0.028
R23898 VBP.n300 VBP.n299 0.028
R23899 VBP.n160 VBP.n153 0.028
R23900 VBP.n199 VBP.n198 0.027
R23901 VBP.n359 VBP.n358 0.026
R23902 VBP.n273 VBP.n272 0.026
R23903 VBP.n196 VBP.n195 0.026
R23904 VBP.n28 VBP.n27 0.026
R23905 VBP.n89 VBP.n88 0.023
R23906 VBP.n358 VBP.n357 0.023
R23907 VBP.n290 VBP.n289 0.023
R23908 VBP.n272 VBP.n271 0.023
R23909 VBP.n162 VBP.n161 0.023
R23910 VBP.n197 VBP.n196 0.023
R23911 VBP.n80 VBP.n79 0.021
R23912 VBP.n87 VBP.n86 0.021
R23913 VBP.n352 VBP.n351 0.021
R23914 VBP.n301 VBP.n300 0.021
R23915 VBP.n275 VBP.n274 0.021
R23916 VBP.n226 VBP.n225 0.021
R23917 VBP.n153 VBP.n152 0.021
R23918 VBP.n188 VBP.n187 0.021
R23919 VBP.n305 VBP.n304 0.019
R23920 VBP.n126 VBP.n111 0.019
R23921 VBP.n341 VBP.n340 0.019
R23922 VBP.n284 VBP.n283 0.019
R23923 VBP.n279 VBP.n278 0.019
R23924 VBP.n326 VBP.n325 0.019
R23925 VBP.n173 VBP.n170 0.019
R23926 VBP.n184 VBP.n179 0.019
R23927 VBP.n2 VBP.n1 0.018
R23928 VBP.n376 VBP.n375 0.017
R23929 VBP.n286 VBP.n285 0.017
R23930 VBP.n281 VBP.n280 0.017
R23931 VBP.n169 VBP.n168 0.017
R23932 VBP.n178 VBP.n177 0.017
R23933 VBP.n201 VBP.n200 0.017
R23934 VBP.n368 VBP.n367 0.015
R23935 VBP.n277 VBP.n276 0.015
R23936 VBP.n186 VBP.n185 0.015
R23937 VBP.n309 VBP.n308 0.015
R23938 VBP.n101 VBP.n100 0.015
R23939 VBP.n216 VBP.n215 0.015
R23940 VBP.n22 VBP.n2 0.015
R23941 VBP.n127 VBP.n109 0.014
R23942 VBP.n315 VBP.n314 0.014
R23943 VBP.n320 VBP.n319 0.014
R23944 VBP.n378 VBP.n377 0.014
R23945 VBP.n362 VBP.n361 0.014
R23946 VBP.n210 VBP.n209 0.014
R23947 VBP.n205 VBP.n204 0.014
R23948 VBP.n104 VBP.n103 0.013
R23949 VBP.n346 VBP.n341 0.013
R23950 VBP.n288 VBP.n287 0.013
R23951 VBP.n331 VBP.n326 0.013
R23952 VBP.n164 VBP.n163 0.013
R23953 VBP.n314 VBP.n313 0.013
R23954 VBP.n332 VBP.n324 0.013
R23955 VBP.n83 VBP.n82 0.013
R23956 VBP.n84 VBP.n83 0.013
R23957 VBP.n348 VBP.n347 0.013
R23958 VBP.n228 VBP.n220 0.013
R23959 VBP.n220 VBP.n219 0.013
R23960 VBP.n211 VBP.n210 0.013
R23961 VBP.n379 VBP.n127 0.012
R23962 VBP.n324 VBP.n323 0.012
R23963 VBP.n349 VBP.n348 0.012
R23964 VBP.n81 VBP.n80 0.011
R23965 VBP.n359 VBP.n352 0.011
R23966 VBP.n274 VBP.n273 0.011
R23967 VBP.n227 VBP.n226 0.011
R23968 VBP.n195 VBP.n188 0.011
R23969 VBP.n311 VBP.n310 0.011
R23970 VBP.n318 VBP.n317 0.011
R23971 VBP.n321 VBP.n320 0.011
R23972 VBP.n109 VBP.n102 0.011
R23973 VBP.n370 VBP.n363 0.011
R23974 VBP.n361 VBP.n360 0.011
R23975 VBP.n214 VBP.n213 0.011
R23976 VBP.n207 VBP.n206 0.011
R23977 VBP.n204 VBP.n203 0.011
R23978 VBP.n19 VBP.n18 0.01
R23979 VBP.n308 VBP.n307 0.01
R23980 VBP.n100 VBP.n99 0.01
R23981 VBP.n217 VBP.n216 0.01
R23982 VBP.n69 VBP.n67 0.01
R23983 VBP.n49 VBP.n47 0.01
R23984 VBP.n23 VBP.n22 0.009
R23985 VBP.n98 VBP.n89 0.009
R23986 VBP.n299 VBP.n290 0.009
R23987 VBP.n161 VBP.n160 0.009
R23988 VBP.n307 VBP.n306 0.009
R23989 VBP.n99 VBP.n85 0.009
R23990 VBP.n218 VBP.n217 0.009
R23991 VBP.n312 VBP.n311 0.008
R23992 VBP.n317 VBP.n316 0.008
R23993 VBP.n322 VBP.n321 0.008
R23994 VBP.n371 VBP.n370 0.008
R23995 VBP.n360 VBP.n350 0.008
R23996 VBP.n213 VBP.n212 0.008
R23997 VBP.n208 VBP.n207 0.008
R23998 VBP.n203 VBP.n202 0.008
R23999 VBP.n233 VBP.n232 0.007
R24000 VBP.n234 VBP.n233 0.007
R24001 VBP.n235 VBP.n234 0.007
R24002 VBP.n236 VBP.n235 0.007
R24003 VBP.n237 VBP.n236 0.007
R24004 VBP.n238 VBP.n237 0.007
R24005 VBP.n239 VBP.n238 0.007
R24006 VBP.n240 VBP.n239 0.007
R24007 VBP.n241 VBP.n240 0.007
R24008 VBP.n242 VBP.n241 0.007
R24009 VBP.n111 VBP.n110 0.007
R24010 VBP.n375 VBP.n374 0.007
R24011 VBP.n138 VBP.n137 0.007
R24012 VBP.n137 VBP.n136 0.007
R24013 VBP.n136 VBP.n135 0.007
R24014 VBP.n135 VBP.n134 0.007
R24015 VBP.n134 VBP.n133 0.007
R24016 VBP.n133 VBP.n132 0.007
R24017 VBP.n132 VBP.n131 0.007
R24018 VBP.n131 VBP.n130 0.007
R24019 VBP.n130 VBP.n129 0.007
R24020 VBP.n129 VBP.n128 0.007
R24021 VBP.n285 VBP.n284 0.007
R24022 VBP.n280 VBP.n279 0.007
R24023 VBP.n170 VBP.n169 0.007
R24024 VBP.n179 VBP.n178 0.007
R24025 VBP.n323 VBP.n322 0.007
R24026 VBP.n350 VBP.n349 0.007
R24027 VBP.n202 VBP.n201 0.007
R24028 VBP.n227 VBP.n224 0.007
R24029 VBP.n81 VBP.n78 0.007
R24030 VBP.n346 VBP.n345 0.006
R24031 VBP.n331 VBP.n330 0.006
R24032 VBP.n31 VBP.n30 0.006
R24033 VBP.n306 VBP.n305 0.006
R24034 VBP.n313 VBP.n312 0.006
R24035 VBP.n333 VBP.n332 0.006
R24036 VBP.n82 VBP.n74 0.006
R24037 VBP.n85 VBP.n84 0.006
R24038 VBP.n347 VBP.n339 0.006
R24039 VBP.n229 VBP.n228 0.006
R24040 VBP.n219 VBP.n218 0.006
R24041 VBP.n212 VBP.n211 0.006
R24042 VBP.n1 VBP.n0 0.006
R24043 VBP.n316 VBP.n315 0.005
R24044 VBP.n377 VBP.n371 0.005
R24045 VBP.n209 VBP.n208 0.005
R24046 VBP.n58 VBP.n56 0.005
R24047 VBP.n38 VBP.n36 0.005
R24048 VBP.n21 VBP.n9 0.005
R24049 VBP.n9 VBP.n8 0.005
R24050 VBP.n74 VBP.n73 0.004
R24051 VBP.n230 VBP.n229 0.004
R24052 VBP.n334 VBP.n333 0.004
R24053 VBP.n339 VBP.n338 0.004
R24054 VBP.n114 VBP.n113 0.004
R24055 VBP.n123 VBP.n114 0.004
R24056 VBP.n119 VBP.n118 0.004
R24057 VBP.n123 VBP.n119 0.004
R24058 VBP.n116 VBP.n115 0.004
R24059 VBP.n121 VBP.n120 0.004
R24060 VBP.n253 VBP.n252 0.004
R24061 VBP.n252 VBP.n251 0.004
R24062 VBP.n247 VBP.n246 0.004
R24063 VBP.n251 VBP.n247 0.004
R24064 VBP.n244 VBP.n243 0.004
R24065 VBP.n249 VBP.n248 0.004
R24066 VBP.n148 VBP.n147 0.004
R24067 VBP.n147 VBP.n146 0.004
R24068 VBP.n145 VBP.n144 0.004
R24069 VBP.n146 VBP.n145 0.004
R24070 VBP.n142 VBP.n141 0.004
R24071 VBP.n140 VBP.n139 0.004
R24072 VBP.n146 VBP.n140 0.004
R24073 VBP.n310 VBP.n309 0.004
R24074 VBP.n319 VBP.n318 0.004
R24075 VBP.n102 VBP.n101 0.004
R24076 VBP.n363 VBP.n362 0.004
R24077 VBP.n215 VBP.n214 0.004
R24078 VBP.n206 VBP.n205 0.004
R24079 VBP.n30 VBP.n29 0.004
R24080 VBP.n122 VBP.n121 0.002
R24081 VBP.n117 VBP.n116 0.002
R24082 VBP.n123 VBP.n117 0.002
R24083 VBP.n123 VBP.n122 0.002
R24084 VBP.n250 VBP.n249 0.002
R24085 VBP.n245 VBP.n244 0.002
R24086 VBP.n251 VBP.n245 0.002
R24087 VBP.n251 VBP.n250 0.002
R24088 VBP.n143 VBP.n142 0.002
R24089 VBP.n146 VBP.n143 0.002
R24090 VBP.n379 VBP.n337 0.002
R24091 VBP.n381 VBP.n380 0.002
R24092 VBP.n337 VBP.n336 0.002
R24093 VBP.n380 VBP.n379 0.002
R24094 VBP.n20 VBP.n19 0.001
R24095 VBP.n21 VBP.n20 0.001
R24096 VBP.n379 VBP.n378 0.001
R24097 VBP.n19 VBP.n12 0.001
R24098 VON.n61 VON.t4 734.909
R24099 VON.n61 VON.t5 238
R24100 VON.n48 VON.t2 28.565
R24101 VON.n7 VON.t3 17.4
R24102 VON.n170 VON.n169 13.176
R24103 VON.n583 VON.n582 13.176
R24104 VON.n152 VON.n151 9.3
R24105 VON.n296 VON.n295 9.3
R24106 VON.n374 VON.n373 9.3
R24107 VON.n520 VON.n519 9.3
R24108 VON.n522 VON.n521 9.3
R24109 VON.n270 VON.n269 9.3
R24110 VON.n163 VON.n162 9.3
R24111 VON.n150 VON.n149 9.3
R24112 VON.n282 VON.n281 9.3
R24113 VON.n293 VON.n292 9.3
R24114 VON.n388 VON.n387 9.3
R24115 VON.n351 VON.n350 9.3
R24116 VON.n376 VON.n375 9.3
R24117 VON.n534 VON.n533 9.3
R24118 VON.n546 VON.n545 9.3
R24119 VON.n581 VON.n580 9.3
R24120 VON.n731 VON.n730 9.3
R24121 VON.n772 VON.n771 9.3
R24122 VON.n49 VON.n48 9.02
R24123 VON.n8 VON.n7 8.5
R24124 VON.n31 VON.n30 8.282
R24125 VON.n669 VON.n668 8.043
R24126 VON.n796 VON.n795 7.029
R24127 VON.n362 VON.n361 5.417
R24128 VON.n519 VON.n518 5.081
R24129 VON.n814 VON.n813 4.767
R24130 VON.n295 VON.n294 4.704
R24131 VON.n92 VON.n89 4.703
R24132 VON.n341 VON.n340 4.65
R24133 VON.n573 VON.n572 4.65
R24134 VON.n751 VON.n750 4.65
R24135 VON.n656 VON.n655 4.5
R24136 VON.n93 VON.n92 4.5
R24137 VON.n84 VON.n83 4.5
R24138 VON.n454 VON.n453 4.5
R24139 VON.n446 VON.n445 4.5
R24140 VON.n97 VON.n78 4.5
R24141 VON.n182 VON.n181 4.5
R24142 VON.n172 VON.n171 4.5
R24143 VON.n156 VON.n155 4.5
R24144 VON.n143 VON.n142 4.5
R24145 VON.n137 VON.n136 4.5
R24146 VON.n278 VON.n277 4.5
R24147 VON.n290 VON.n289 4.5
R24148 VON.n308 VON.n307 4.5
R24149 VON.n328 VON.n327 4.5
R24150 VON.n321 VON.n320 4.5
R24151 VON.n314 VON.n313 4.5
R24152 VON.n336 VON.n335 4.5
R24153 VON.n392 VON.n391 4.5
R24154 VON.n354 VON.n353 4.5
R24155 VON.n381 VON.n380 4.5
R24156 VON.n369 VON.n365 4.5
R24157 VON.n484 VON.n474 4.5
R24158 VON.n462 VON.n461 4.5
R24159 VON.n479 VON.n476 4.5
R24160 VON.n526 VON.n525 4.5
R24161 VON.n551 VON.n550 4.5
R24162 VON.n538 VON.n537 4.5
R24163 VON.n621 VON.n620 4.5
R24164 VON.n585 VON.n584 4.5
R24165 VON.n629 VON.n628 4.5
R24166 VON.n644 VON.n643 4.5
R24167 VON.n636 VON.n635 4.5
R24168 VON.n102 VON.n101 4.5
R24169 VON.n10 VON.n9 4.5
R24170 VON.n3 VON.n2 4.5
R24171 VON.n35 VON.n31 4.5
R24172 VON.n41 VON.n40 4.5
R24173 VON.n55 VON.n46 4.5
R24174 VON.n52 VON.n50 4.5
R24175 VON.n807 VON.n806 4.5
R24176 VON.n788 VON.n787 4.5
R24177 VON.n778 VON.n777 4.5
R24178 VON.n766 VON.n765 4.5
R24179 VON.n717 VON.n716 4.5
R24180 VON.n727 VON.n726 4.5
R24181 VON.n759 VON.n758 4.5
R24182 VON.n753 VON.n752 4.5
R24183 VON.n749 VON.n748 4.5
R24184 VON.n745 VON.n744 4.5
R24185 VON.n739 VON.n738 4.5
R24186 VON.n677 VON.n676 4.5
R24187 VON.n679 VON.n669 4.473
R24188 VON.n668 VON.t1 4.35
R24189 VON.n136 VON.n133 4.328
R24190 VON.n643 VON.n642 4.326
R24191 VON.n9 VON.n6 4.141
R24192 VON.n50 VON.n47 4.141
R24193 VON.n716 VON.n713 4.141
R24194 VON.n787 VON.n786 4.141
R24195 VON.n628 VON.n627 3.951
R24196 VON.n365 VON.n363 3.946
R24197 VON.n91 VON.n90 3.764
R24198 VON.n40 VON.n39 3.764
R24199 VON.n31 VON.n29 3.764
R24200 VON.n726 VON.n723 3.764
R24201 VON.n765 VON.n763 3.764
R24202 VON.n453 VON.n450 3.572
R24203 VON.n335 VON.n334 3.569
R24204 VON.n312 VON.n311 3.388
R24205 VON.n2 VON.n1 3.388
R24206 VON.n46 VON.n45 3.388
R24207 VON.n676 VON.n673 3.388
R24208 VON.n738 VON.n737 3.388
R24209 VON.n777 VON.n776 3.388
R24210 VON.n806 VON.n805 3.388
R24211 VON.n474 VON.n471 3.197
R24212 VON.n320 VON.n319 3.195
R24213 VON.n300 VON.n299 3.033
R24214 VON.n398 VON.n362 3.033
R24215 VON.n345 VON.n344 3.033
R24216 VON.n574 VON.n570 3.033
R24217 VON.n662 VON.n661 3.033
R24218 VON.n452 VON.n451 3.011
R24219 VON.n676 VON.n675 3.011
R24220 VON.n738 VON.n735 3.011
R24221 VON.n744 VON.n742 3.011
R24222 VON.n771 VON.n770 3.011
R24223 VON.n777 VON.n775 3.011
R24224 VON.n806 VON.n804 3.011
R24225 VON.n360 VON.t0 2.856
R24226 VON.n307 VON.n306 2.82
R24227 VON.n814 VON.n667 2.722
R24228 VON.n78 VON.n77 2.635
R24229 VON.n634 VON.n633 2.635
R24230 VON.n40 VON.n38 2.635
R24231 VON.n726 VON.n725 2.635
R24232 VON.n730 VON.n729 2.635
R24233 VON.n758 VON.n757 2.635
R24234 VON.n765 VON.n764 2.635
R24235 VON.n815 VON.n814 2.448
R24236 VON.n307 VON.n305 2.258
R24237 VON.n655 VON.n654 2.258
R24238 VON.n9 VON.n8 2.258
R24239 VON.n50 VON.n49 2.258
R24240 VON.n716 VON.n715 2.258
R24241 VON.n787 VON.n785 2.258
R24242 VON.n83 VON.n82 1.882
R24243 VON.n445 VON.n444 1.882
R24244 VON.n474 VON.n473 1.882
R24245 VON.n361 VON.n360 1.844
R24246 VON.n135 VON.n134 1.505
R24247 VON.n320 VON.n318 1.505
R24248 VON.n327 VON.n326 1.505
R24249 VON.n626 VON.n625 1.505
R24250 VON.n628 VON.n626 1.505
R24251 VON.n635 VON.n634 1.505
R24252 VON.n758 VON.n756 1.505
R24253 VON.n657 VON.n656 1.5
R24254 VON.n183 VON.n182 1.5
R24255 VON.n173 VON.n172 1.5
R24256 VON.n485 VON.n484 1.5
R24257 VON.n463 VON.n462 1.5
R24258 VON.n552 VON.n551 1.5
R24259 VON.n586 VON.n585 1.5
R24260 VON.n663 VON.n662 1.5
R24261 VON.n645 VON.n644 1.5
R24262 VON.n103 VON.n102 1.5
R24263 VON.n12 VON.n11 1.384
R24264 VON.n43 VON.n42 1.384
R24265 VON.n60 VON.n59 1.148
R24266 VON.n13 VON.n12 1.146
R24267 VON.n23 VON.n22 1.137
R24268 VON.n19 VON.n18 1.137
R24269 VON.n44 VON.n43 1.137
R24270 VON.n136 VON.n135 1.129
R24271 VON.n142 VON.n141 1.129
R24272 VON.n277 VON.n276 1.129
R24273 VON.n326 VON.n325 1.129
R24274 VON.n444 VON.n443 1.129
R24275 VON.n453 VON.n452 1.129
R24276 VON.n461 VON.n460 1.129
R24277 VON.n537 VON.n536 1.129
R24278 VON.n744 VON.n743 1.129
R24279 VON.n808 VON.n807 1.125
R24280 VON.n408 VON.n398 1.042
R24281 VON.n60 VON.n44 1.019
R24282 VON VON.n60 0.876
R24283 VON.n189 VON.n188 0.853
R24284 VON.n234 VON.n233 0.853
R24285 VON.n409 VON.n408 0.853
R24286 VON.n488 VON.n487 0.853
R24287 VON.n588 VON.n587 0.853
R24288 VON.n666 VON.n665 0.853
R24289 VON.n289 VON.n288 0.752
R24290 VON.n305 VON.n304 0.752
R24291 VON.n313 VON.n312 0.752
R24292 VON.n335 VON.n333 0.752
R24293 VON.n353 VON.n352 0.752
R24294 VON.n391 VON.n390 0.752
R24295 VON.n473 VON.n472 0.752
R24296 VON.n620 VON.n619 0.752
R24297 VON.n643 VON.n641 0.752
R24298 VON.n680 VON.n679 0.75
R24299 VON.n105 VON.n104 0.704
R24300 VON.n795 VON.n794 0.445
R24301 VON.n58 VON.n55 0.443
R24302 VON.n675 VON.n674 0.414
R24303 VON.n804 VON.n803 0.414
R24304 VON.n715 VON.n714 0.382
R24305 VON.n785 VON.n784 0.382
R24306 VON.n101 VON.n100 0.376
R24307 VON.n77 VON.n76 0.376
R24308 VON.n92 VON.n91 0.376
R24309 VON.n155 VON.n154 0.376
R24310 VON.n171 VON.n170 0.376
R24311 VON.n181 VON.n180 0.376
R24312 VON.n380 VON.n379 0.376
R24313 VON.n365 VON.n364 0.376
R24314 VON.n476 VON.n475 0.376
R24315 VON.n525 VON.n524 0.376
R24316 VON.n550 VON.n549 0.376
R24317 VON.n584 VON.n583 0.376
R24318 VON.n654 VON.n653 0.376
R24319 VON.n59 VON.n58 0.288
R24320 VON VON.n815 0.251
R24321 VON.n162 VON.n161 0.189
R24322 VON.n269 VON.n268 0.189
R24323 VON.n545 VON.n544 0.189
R24324 VON.n580 VON.n579 0.189
R24325 VON.n149 VON.n148 0.177
R24326 VON.n281 VON.n280 0.177
R24327 VON.n533 VON.n532 0.177
R24328 VON.n572 VON.n571 0.177
R24329 VON.n379 VON.n378 0.121
R24330 VON.n344 VON.n343 0.121
R24331 VON.n679 VON.n678 0.113
R24332 VON.n390 VON.n389 0.109
R24333 VON.n689 VON.n688 0.1
R24334 VON.n703 VON.n702 0.1
R24335 VON.n725 VON.n724 0.072
R24336 VON.n775 VON.n774 0.072
R24337 VON.n58 VON.n57 0.067
R24338 VON.n671 VON.n670 0.06
R24339 VON.n720 VON.n719 0.06
R24340 VON.n732 VON.n731 0.06
R24341 VON.n772 VON.n769 0.06
R24342 VON.n782 VON.n781 0.06
R24343 VON.n792 VON.n791 0.06
R24344 VON.n801 VON.n800 0.06
R24345 VON.n682 VON.n681 0.06
R24346 VON.n686 VON.n685 0.06
R24347 VON.n706 VON.n705 0.06
R24348 VON.n710 VON.n709 0.06
R24349 VON.n810 VON.n809 0.06
R24350 VON.n692 VON.n691 0.055
R24351 VON.n696 VON.n695 0.055
R24352 VON.n700 VON.n699 0.055
R24353 VON.n681 VON.n680 0.052
R24354 VON.n809 VON.n808 0.052
R24355 VON.n749 VON.n747 0.05
R24356 VON.n759 VON.n755 0.05
R24357 VON.n695 VON.n694 0.05
R24358 VON.n699 VON.n698 0.05
R24359 VON.n808 VON.n710 0.05
R24360 VON.n746 VON.n745 0.048
R24361 VON.n754 VON.n753 0.048
R24362 VON.n693 VON.n692 0.048
R24363 VON.n697 VON.n696 0.048
R24364 VON.n166 VON.n165 0.047
R24365 VON.n297 VON.n296 0.047
R24366 VON.n567 VON.n566 0.047
R24367 VON.n264 VON.n263 0.047
R24368 VON.n300 VON.n298 0.045
R24369 VON.n357 VON.n356 0.045
R24370 VON.n359 VON.n358 0.045
R24371 VON.n531 VON.n530 0.045
R24372 VON.n219 VON.n218 0.045
R24373 VON.n404 VON.n403 0.045
R24374 VON.n145 VON.n144 0.043
R24375 VON.n284 VON.n283 0.043
R24376 VON.n323 VON.n322 0.043
R24377 VON.n397 VON.n396 0.043
R24378 VON.n395 VON.n394 0.043
R24379 VON.n449 VON.n448 0.043
R24380 VON.n479 VON.n478 0.043
R24381 VON.n618 VON.n617 0.043
R24382 VON.n122 VON.n121 0.043
R24383 VON.n229 VON.n228 0.043
R24384 VON.n439 VON.n438 0.043
R24385 VON.n468 VON.n467 0.043
R24386 VON.n605 VON.n604 0.043
R24387 VON.n685 VON.n684 0.043
R24388 VON.n709 VON.n708 0.043
R24389 VON.n813 VON.n812 0.043
R24390 VON.n398 VON.n397 0.041
R24391 VON.n529 VON.n528 0.041
R24392 VON.n408 VON.n407 0.041
R24393 VON.n505 VON.n504 0.041
R24394 VON.n683 VON.n682 0.04
R24395 VON.n691 VON.n690 0.04
R24396 VON.n707 VON.n706 0.04
R24397 VON.n811 VON.n810 0.04
R24398 VON.n158 VON.n157 0.039
R24399 VON.n286 VON.n285 0.039
R24400 VON.n314 VON.n310 0.039
R24401 VON.n398 VON.n359 0.039
R24402 VON.n129 VON.n128 0.039
R24403 VON.n212 VON.n211 0.039
R24404 VON.n233 VON.n232 0.039
R24405 VON.n408 VON.n267 0.039
R24406 VON.n426 VON.n425 0.039
R24407 VON.n486 VON.n485 0.039
R24408 VON.n701 VON.n700 0.038
R24409 VON.n160 VON.n159 0.037
R24410 VON.n309 VON.n308 0.037
R24411 VON.n341 VON.n339 0.037
R24412 VON.n346 VON.n345 0.037
R24413 VON.n383 VON.n382 0.037
R24414 VON.n462 VON.n459 0.037
R24415 VON.n543 VON.n542 0.037
R24416 VON.n576 VON.n575 0.037
R24417 VON.n223 VON.n222 0.037
R24418 VON.n256 VON.n255 0.037
R24419 VON.n487 VON.n463 0.037
R24420 VON.n561 VON.n560 0.037
R24421 VON.n737 VON.n736 0.036
R24422 VON.n763 VON.n762 0.036
R24423 VON.n791 VON.n790 0.036
R24424 VON.n800 VON.n799 0.036
R24425 VON.n272 VON.n271 0.035
R24426 VON.n374 VON.n372 0.035
R24427 VON.n578 VON.n577 0.035
R24428 VON.n184 VON.n183 0.035
R24429 VON.n553 VON.n552 0.035
R24430 VON.n34 VON.n33 0.035
R24431 VON.n33 VON.n32 0.035
R24432 VON.n22 VON.n21 0.035
R24433 VON.n104 VON.n103 0.035
R24434 VON.n167 VON.n166 0.034
R24435 VON.n328 VON.n324 0.034
R24436 VON.n338 VON.n337 0.034
R24437 VON.n131 VON.n130 0.034
R24438 VON.n188 VON.n187 0.034
R24439 VON.n221 VON.n220 0.034
R24440 VON.n251 VON.n250 0.034
R24441 VON.n266 VON.n265 0.034
R24442 VON.n406 VON.n405 0.034
R24443 VON.n470 VON.n469 0.034
R24444 VON.n586 VON.n564 0.034
R24445 VON.n563 VON.n562 0.034
R24446 VON.n672 VON.n671 0.033
R24447 VON.n781 VON.n780 0.033
R24448 VON.n705 VON.n704 0.033
R24449 VON.n371 VON.n370 0.032
R24450 VON.n447 VON.n446 0.032
R24451 VON.n568 VON.n567 0.032
R24452 VON.n574 VON.n573 0.032
R24453 VON.n173 VON.n132 0.032
R24454 VON.n210 VON.n209 0.032
R24455 VON.n231 VON.n230 0.032
R24456 VON.n253 VON.n252 0.032
R24457 VON.n254 VON.n253 0.032
R24458 VON.n428 VON.n427 0.032
R24459 VON.n429 VON.n428 0.032
R24460 VON.n431 VON.n430 0.032
R24461 VON.n507 VON.n506 0.032
R24462 VON.n587 VON.n556 0.032
R24463 VON.n106 VON.n105 0.031
R24464 VON.n117 VON.n116 0.031
R24465 VON.n191 VON.n190 0.031
R24466 VON.n202 VON.n201 0.031
R24467 VON.n236 VON.n235 0.031
R24468 VON.n247 VON.n246 0.031
R24469 VON.n411 VON.n410 0.031
R24470 VON.n422 VON.n421 0.031
R24471 VON.n490 VON.n489 0.031
R24472 VON.n501 VON.n500 0.031
R24473 VON.n590 VON.n589 0.031
R24474 VON.n601 VON.n600 0.031
R24475 VON.n721 VON.n720 0.031
R24476 VON.n793 VON.n792 0.031
R24477 VON.n802 VON.n801 0.031
R24478 VON.n687 VON.n686 0.031
R24479 VON.n688 VON.n687 0.031
R24480 VON.n153 VON.n152 0.03
R24481 VON.n172 VON.n163 0.03
R24482 VON.n349 VON.n348 0.03
R24483 VON.n585 VON.n581 0.03
R24484 VON.n662 VON.n660 0.03
R24485 VON.n120 VON.n119 0.03
R24486 VON.n126 VON.n125 0.03
R24487 VON.n186 VON.n185 0.03
R24488 VON.n206 VON.n205 0.03
R24489 VON.n216 VON.n215 0.03
R24490 VON.n441 VON.n440 0.03
R24491 VON.n465 VON.n464 0.03
R24492 VON.n511 VON.n510 0.03
R24493 VON.n558 VON.n557 0.03
R24494 VON.n665 VON.n663 0.03
R24495 VON.n102 VON.n99 0.028
R24496 VON.n96 VON.n95 0.028
R24497 VON.n354 VON.n351 0.028
R24498 VON.n392 VON.n388 0.028
R24499 VON.n386 VON.n385 0.028
R24500 VON.n652 VON.n651 0.028
R24501 VON.n72 VON.n71 0.028
R24502 VON.n555 VON.n554 0.028
R24503 VON.n607 VON.n606 0.028
R24504 VON.n649 VON.n648 0.028
R24505 VON.n719 VON.n718 0.028
R24506 VON.n753 VON.n751 0.028
R24507 VON.n704 VON.n703 0.028
R24508 VON.n110 VON.n109 0.027
R24509 VON.n113 VON.n112 0.027
R24510 VON.n195 VON.n194 0.027
R24511 VON.n198 VON.n197 0.027
R24512 VON.n240 VON.n239 0.027
R24513 VON.n243 VON.n242 0.027
R24514 VON.n415 VON.n414 0.027
R24515 VON.n418 VON.n417 0.027
R24516 VON.n494 VON.n493 0.027
R24517 VON.n497 VON.n496 0.027
R24518 VON.n594 VON.n593 0.027
R24519 VON.n597 VON.n596 0.027
R24520 VON.n23 VON.n19 0.027
R24521 VON.n94 VON.n93 0.026
R24522 VON.n342 VON.n341 0.026
R24523 VON.n377 VON.n376 0.026
R24524 VON.n616 VON.n615 0.026
R24525 VON.n603 VON.n602 0.026
R24526 VON.n751 VON.n749 0.026
R24527 VON.n783 VON.n782 0.026
R24528 VON.n140 VON.n139 0.024
R24529 VON.n147 VON.n146 0.024
R24530 VON.n275 VON.n274 0.024
R24531 VON.n302 VON.n301 0.024
R24532 VON.n482 VON.n481 0.024
R24533 VON.n540 VON.n539 0.024
R24534 VON.n623 VON.n622 0.024
R24535 VON.n636 VON.n632 0.024
R24536 VON.n74 VON.n73 0.024
R24537 VON.n124 VON.n123 0.024
R24538 VON.n612 VON.n611 0.024
R24539 VON.n727 VON.n722 0.024
R24540 VON.n731 VON.n728 0.024
R24541 VON.n766 VON.n761 0.024
R24542 VON.n769 VON.n768 0.024
R24543 VON.n702 VON.n701 0.024
R24544 VON.n84 VON.n81 0.022
R24545 VON.n81 VON.n80 0.022
R24546 VON.n632 VON.n631 0.022
R24547 VON.n65 VON.n64 0.022
R24548 VON.n64 VON.n63 0.022
R24549 VON.n611 VON.n610 0.022
R24550 VON.n645 VON.n614 0.022
R24551 VON.n658 VON.n657 0.022
R24552 VON.n678 VON.n677 0.021
R24553 VON.n733 VON.n732 0.021
R24554 VON.n734 VON.n733 0.021
R24555 VON.n740 VON.n739 0.021
R24556 VON.n768 VON.n767 0.021
R24557 VON.n773 VON.n772 0.021
R24558 VON.n779 VON.n778 0.021
R24559 VON.n807 VON.n802 0.021
R24560 VON.n690 VON.n689 0.021
R24561 VON.n95 VON.n94 0.02
R24562 VON.n80 VON.n79 0.02
R24563 VON.n150 VON.n147 0.02
R24564 VON.n526 VON.n523 0.02
R24565 VON.n631 VON.n630 0.02
R24566 VON.n651 VON.n650 0.02
R24567 VON.n71 VON.n70 0.02
R24568 VON.n68 VON.n67 0.02
R24569 VON.n63 VON.n62 0.02
R24570 VON.n208 VON.n207 0.02
R24571 VON.n503 VON.n502 0.02
R24572 VON.n515 VON.n514 0.02
R24573 VON.n610 VON.n609 0.02
R24574 VON.n648 VON.n647 0.02
R24575 VON.n663 VON.n658 0.02
R24576 VON.n10 VON.n5 0.02
R24577 VON.n53 VON.n52 0.02
R24578 VON.n189 VON.n117 0.019
R24579 VON.n190 VON.n189 0.019
R24580 VON.n234 VON.n202 0.019
R24581 VON.n235 VON.n234 0.019
R24582 VON.n409 VON.n247 0.019
R24583 VON.n410 VON.n409 0.019
R24584 VON.n488 VON.n422 0.019
R24585 VON.n489 VON.n488 0.019
R24586 VON.n588 VON.n501 0.019
R24587 VON.n589 VON.n588 0.019
R24588 VON.n677 VON.n672 0.019
R24589 VON.n717 VON.n712 0.019
R24590 VON.n739 VON.n734 0.019
R24591 VON.n745 VON.n741 0.019
R24592 VON.n778 VON.n773 0.019
R24593 VON.n789 VON.n788 0.019
R24594 VON.n807 VON.n793 0.019
R24595 VON.n798 VON.n797 0.019
R24596 VON.n684 VON.n683 0.019
R24597 VON.n708 VON.n707 0.019
R24598 VON.n812 VON.n811 0.019
R24599 VON.n88 VON.n87 0.018
R24600 VON.n291 VON.n290 0.018
R24601 VON.n385 VON.n384 0.018
R24602 VON.n541 VON.n540 0.018
R24603 VON.n640 VON.n639 0.018
R24604 VON.n103 VON.n74 0.018
R24605 VON.n175 VON.n174 0.018
R24606 VON.n214 VON.n213 0.018
R24607 VON.n401 VON.n400 0.018
R24608 VON.n424 VON.n423 0.018
R24609 VON.n509 VON.n508 0.018
R24610 VON.n512 VON.n511 0.018
R24611 VON.n556 VON.n555 0.018
R24612 VON.n41 VON.n37 0.018
R24613 VON.n36 VON.n35 0.018
R24614 VON.n274 VON.n273 0.017
R24615 VON.n316 VON.n315 0.017
R24616 VON.n331 VON.n330 0.017
R24617 VON.n348 VON.n347 0.017
R24618 VON.n370 VON.n369 0.017
R24619 VON.n367 VON.n366 0.017
R24620 VON.n457 VON.n456 0.017
R24621 VON.n547 VON.n546 0.017
R24622 VON.n630 VON.n629 0.017
R24623 VON.n70 VON.n69 0.017
R24624 VON.n67 VON.n66 0.017
R24625 VON.n125 VON.n124 0.017
R24626 VON.n187 VON.n186 0.017
R24627 VON.n177 VON.n176 0.017
R24628 VON.n205 VON.n204 0.017
R24629 VON.n215 VON.n214 0.017
R24630 VON.n227 VON.n226 0.017
R24631 VON.n226 VON.n225 0.017
R24632 VON.n258 VON.n257 0.017
R24633 VON.n259 VON.n258 0.017
R24634 VON.n261 VON.n260 0.017
R24635 VON.n432 VON.n431 0.017
R24636 VON.n434 VON.n433 0.017
R24637 VON.n437 VON.n436 0.017
R24638 VON.n514 VON.n513 0.017
R24639 VON.n517 VON.n516 0.017
R24640 VON.n609 VON.n608 0.017
R24641 VON.n614 VON.n613 0.017
R24642 VON.n647 VON.n646 0.017
R24643 VON.n4 VON.n3 0.017
R24644 VON.n17 VON.n16 0.017
R24645 VON.n55 VON.n54 0.017
R24646 VON.n666 VON.n601 0.016
R24647 VON.n728 VON.n727 0.016
R24648 VON.n760 VON.n759 0.016
R24649 VON.n767 VON.n766 0.016
R24650 VON.n317 VON.n316 0.015
R24651 VON.n337 VON.n336 0.015
R24652 VON.n456 VON.n455 0.015
R24653 VON.n188 VON.n173 0.015
R24654 VON.n250 VON.n249 0.015
R24655 VON.n262 VON.n261 0.015
R24656 VON.n402 VON.n401 0.015
R24657 VON.n435 VON.n434 0.015
R24658 VON.n436 VON.n435 0.015
R24659 VON.n587 VON.n586 0.015
R24660 VON.n608 VON.n607 0.015
R24661 VON.n43 VON.n28 0.015
R24662 VON.n27 VON.n26 0.015
R24663 VON.n16 VON.n15 0.015
R24664 VON.n667 VON.n666 0.014
R24665 VON.n718 VON.n717 0.014
R24666 VON.n741 VON.n740 0.014
R24667 VON.n761 VON.n760 0.014
R24668 VON.n788 VON.n783 0.014
R24669 VON.n98 VON.n97 0.013
R24670 VON.n87 VON.n86 0.013
R24671 VON.n168 VON.n167 0.013
R24672 VON.n182 VON.n179 0.013
R24673 VON.n279 VON.n278 0.013
R24674 VON.n282 VON.n279 0.013
R24675 VON.n535 VON.n534 0.013
R24676 VON.n538 VON.n535 0.013
R24677 VON.n551 VON.n547 0.013
R24678 VON.n569 VON.n568 0.013
R24679 VON.n639 VON.n638 0.013
R24680 VON.n119 VON.n118 0.013
R24681 VON.n183 VON.n177 0.013
R24682 VON.n207 VON.n206 0.013
R24683 VON.n217 VON.n216 0.013
R24684 VON.n225 VON.n224 0.013
R24685 VON.n249 VON.n248 0.013
R24686 VON.n260 VON.n259 0.013
R24687 VON.n463 VON.n441 0.013
R24688 VON.n508 VON.n507 0.013
R24689 VON.n510 VON.n509 0.013
R24690 VON.n552 VON.n517 0.013
R24691 VON.n42 VON.n41 0.013
R24692 VON.n12 VON.n0 0.013
R24693 VON.n57 VON.n56 0.013
R24694 VON.n111 VON.n110 0.012
R24695 VON.n112 VON.n111 0.012
R24696 VON.n196 VON.n195 0.012
R24697 VON.n197 VON.n196 0.012
R24698 VON.n241 VON.n240 0.012
R24699 VON.n242 VON.n241 0.012
R24700 VON.n416 VON.n415 0.012
R24701 VON.n417 VON.n416 0.012
R24702 VON.n495 VON.n494 0.012
R24703 VON.n496 VON.n495 0.012
R24704 VON.n595 VON.n594 0.012
R24705 VON.n596 VON.n595 0.012
R24706 VON.n271 VON.n270 0.011
R24707 VON.n273 VON.n272 0.011
R24708 VON.n308 VON.n303 0.011
R24709 VON.n347 VON.n346 0.011
R24710 VON.n372 VON.n371 0.011
R24711 VON.n577 VON.n576 0.011
R24712 VON.n575 VON.n574 0.011
R24713 VON.n656 VON.n652 0.011
R24714 VON.n176 VON.n175 0.011
R24715 VON.n204 VON.n203 0.011
R24716 VON.n209 VON.n208 0.011
R24717 VON.n232 VON.n231 0.011
R24718 VON.n257 VON.n256 0.011
R24719 VON.n267 VON.n266 0.011
R24720 VON.n400 VON.n399 0.011
R24721 VON.n430 VON.n429 0.011
R24722 VON.n433 VON.n432 0.011
R24723 VON.n466 VON.n465 0.011
R24724 VON.n562 VON.n561 0.011
R24725 VON.n560 VON.n559 0.011
R24726 VON.n657 VON.n649 0.011
R24727 VON.n108 VON.n107 0.011
R24728 VON.n115 VON.n114 0.011
R24729 VON.n193 VON.n192 0.011
R24730 VON.n200 VON.n199 0.011
R24731 VON.n238 VON.n237 0.011
R24732 VON.n245 VON.n244 0.011
R24733 VON.n413 VON.n412 0.011
R24734 VON.n420 VON.n419 0.011
R24735 VON.n492 VON.n491 0.011
R24736 VON.n499 VON.n498 0.011
R24737 VON.n592 VON.n591 0.011
R24738 VON.n599 VON.n598 0.011
R24739 VON.n11 VON.n10 0.011
R24740 VON.n52 VON.n51 0.011
R24741 VON.n97 VON.n96 0.009
R24742 VON.n157 VON.n156 0.009
R24743 VON.n159 VON.n158 0.009
R24744 VON.n293 VON.n291 0.009
R24745 VON.n332 VON.n331 0.009
R24746 VON.n339 VON.n338 0.009
R24747 VON.n384 VON.n383 0.009
R24748 VON.n368 VON.n367 0.009
R24749 VON.n446 VON.n442 0.009
R24750 VON.n484 VON.n483 0.009
R24751 VON.n523 VON.n522 0.009
R24752 VON.n542 VON.n541 0.009
R24753 VON.n546 VON.n543 0.009
R24754 VON.n73 VON.n72 0.009
R24755 VON.n69 VON.n68 0.009
R24756 VON.n128 VON.n127 0.009
R24757 VON.n130 VON.n129 0.009
R24758 VON.n213 VON.n212 0.009
R24759 VON.n252 VON.n251 0.009
R24760 VON.n407 VON.n406 0.009
R24761 VON.n425 VON.n424 0.009
R24762 VON.n513 VON.n512 0.009
R24763 VON.n516 VON.n515 0.009
R24764 VON.n28 VON.n27 0.009
R24765 VON.n44 VON.n25 0.009
R24766 VON.n24 VON.n23 0.009
R24767 VON.n19 VON.n14 0.009
R24768 VON.n747 VON.n746 0.009
R24769 VON.n755 VON.n754 0.009
R24770 VON.n694 VON.n693 0.009
R24771 VON.n698 VON.n697 0.009
R24772 VON.n665 VON.n664 0.008
R24773 VON.n139 VON.n138 0.007
R24774 VON.n283 VON.n282 0.007
R24775 VON.n310 VON.n309 0.007
R24776 VON.n321 VON.n317 0.007
R24777 VON.n329 VON.n328 0.007
R24778 VON.n459 VON.n458 0.007
R24779 VON.n624 VON.n623 0.007
R24780 VON.n629 VON.n624 0.007
R24781 VON.n127 VON.n126 0.007
R24782 VON.n233 VON.n223 0.007
R24783 VON.n487 VON.n486 0.007
R24784 VON.n504 VON.n503 0.007
R24785 VON.n646 VON.n645 0.007
R24786 VON.n18 VON.n17 0.007
R24787 VON.n712 VON.n711 0.007
R24788 VON.n722 VON.n721 0.007
R24789 VON.n780 VON.n779 0.007
R24790 VON.n790 VON.n789 0.007
R24791 VON.n107 VON.n106 0.006
R24792 VON.n109 VON.n108 0.006
R24793 VON.n114 VON.n113 0.006
R24794 VON.n116 VON.n115 0.006
R24795 VON.n192 VON.n191 0.006
R24796 VON.n194 VON.n193 0.006
R24797 VON.n199 VON.n198 0.006
R24798 VON.n201 VON.n200 0.006
R24799 VON.n237 VON.n236 0.006
R24800 VON.n239 VON.n238 0.006
R24801 VON.n244 VON.n243 0.006
R24802 VON.n246 VON.n245 0.006
R24803 VON.n412 VON.n411 0.006
R24804 VON.n414 VON.n413 0.006
R24805 VON.n419 VON.n418 0.006
R24806 VON.n421 VON.n420 0.006
R24807 VON.n491 VON.n490 0.006
R24808 VON.n493 VON.n492 0.006
R24809 VON.n498 VON.n497 0.006
R24810 VON.n500 VON.n499 0.006
R24811 VON.n591 VON.n590 0.006
R24812 VON.n593 VON.n592 0.006
R24813 VON.n598 VON.n597 0.006
R24814 VON.n600 VON.n599 0.006
R24815 VON.n85 VON.n84 0.005
R24816 VON.n138 VON.n137 0.005
R24817 VON.n143 VON.n140 0.005
R24818 VON.n278 VON.n275 0.005
R24819 VON.n287 VON.n286 0.005
R24820 VON.n324 VON.n323 0.005
R24821 VON.n330 VON.n329 0.005
R24822 VON.n345 VON.n342 0.005
R24823 VON.n388 VON.n386 0.005
R24824 VON.n448 VON.n447 0.005
R24825 VON.n455 VON.n454 0.005
R24826 VON.n462 VON.n457 0.005
R24827 VON.n478 VON.n477 0.005
R24828 VON.n528 VON.n527 0.005
R24829 VON.n534 VON.n531 0.005
R24830 VON.n539 VON.n538 0.005
R24831 VON.n566 VON.n565 0.005
R24832 VON.n66 VON.n65 0.005
R24833 VON.n222 VON.n221 0.005
R24834 VON.n228 VON.n227 0.005
R24835 VON.n255 VON.n254 0.005
R24836 VON.n438 VON.n437 0.005
R24837 VON.n469 VON.n468 0.005
R24838 VON.n467 VON.n466 0.005
R24839 VON.n554 VON.n553 0.005
R24840 VON.n559 VON.n558 0.005
R24841 VON.n37 VON.n36 0.005
R24842 VON.n35 VON.n34 0.005
R24843 VON.n5 VON.n4 0.005
R24844 VON.n22 VON.n20 0.005
R24845 VON.n25 VON.n24 0.005
R24846 VON.n14 VON.n13 0.005
R24847 VON.n54 VON.n53 0.005
R24848 VON.n797 VON.n796 0.005
R24849 VON.n799 VON.n798 0.004
R24850 VON.n86 VON.n85 0.003
R24851 VON.n146 VON.n145 0.003
R24852 VON.n165 VON.n164 0.003
R24853 VON.n285 VON.n284 0.003
R24854 VON.n290 VON.n287 0.003
R24855 VON.n296 VON.n293 0.003
R24856 VON.n298 VON.n297 0.003
R24857 VON.n301 VON.n300 0.003
R24858 VON.n303 VON.n302 0.003
R24859 VON.n315 VON.n314 0.003
R24860 VON.n336 VON.n332 0.003
R24861 VON.n351 VON.n349 0.003
R24862 VON.n396 VON.n395 0.003
R24863 VON.n381 VON.n377 0.003
R24864 VON.n454 VON.n449 0.003
R24865 VON.n483 VON.n482 0.003
R24866 VON.n481 VON.n480 0.003
R24867 VON.n581 VON.n578 0.003
R24868 VON.n621 VON.n618 0.003
R24869 VON.n622 VON.n621 0.003
R24870 VON.n637 VON.n636 0.003
R24871 VON.n638 VON.n637 0.003
R24872 VON.n644 VON.n640 0.003
R24873 VON.n123 VON.n122 0.003
R24874 VON.n132 VON.n131 0.003
R24875 VON.n185 VON.n184 0.003
R24876 VON.n211 VON.n210 0.003
R24877 VON.n218 VON.n217 0.003
R24878 VON.n220 VON.n219 0.003
R24879 VON.n405 VON.n404 0.003
R24880 VON.n427 VON.n426 0.003
R24881 VON.n440 VON.n439 0.003
R24882 VON.n485 VON.n470 0.003
R24883 VON.n606 VON.n605 0.003
R24884 VON.n613 VON.n612 0.003
R24885 VON.n102 VON.n75 0.001
R24886 VON.n99 VON.n98 0.001
R24887 VON.n93 VON.n88 0.001
R24888 VON.n144 VON.n143 0.001
R24889 VON.n152 VON.n150 0.001
R24890 VON.n156 VON.n153 0.001
R24891 VON.n163 VON.n160 0.001
R24892 VON.n172 VON.n168 0.001
R24893 VON.n182 VON.n178 0.001
R24894 VON.n322 VON.n321 0.001
R24895 VON.n355 VON.n354 0.001
R24896 VON.n356 VON.n355 0.001
R24897 VON.n358 VON.n357 0.001
R24898 VON.n394 VON.n393 0.001
R24899 VON.n393 VON.n392 0.001
R24900 VON.n382 VON.n381 0.001
R24901 VON.n376 VON.n374 0.001
R24902 VON.n369 VON.n368 0.001
R24903 VON.n480 VON.n479 0.001
R24904 VON.n522 VON.n520 0.001
R24905 VON.n527 VON.n526 0.001
R24906 VON.n530 VON.n529 0.001
R24907 VON.n551 VON.n548 0.001
R24908 VON.n585 VON.n569 0.001
R24909 VON.n617 VON.n616 0.001
R24910 VON.n660 VON.n659 0.001
R24911 VON.n121 VON.n120 0.001
R24912 VON.n230 VON.n229 0.001
R24913 VON.n263 VON.n262 0.001
R24914 VON.n265 VON.n264 0.001
R24915 VON.n403 VON.n402 0.001
R24916 VON.n506 VON.n505 0.001
R24917 VON.n564 VON.n563 0.001
R24918 VON.n604 VON.n603 0.001
R24919 VON.n815 VON.n61 0.001
R24920 net3_ota.n510 net3_ota.t3 39.136
R24921 net3_ota.n38 net3_ota.t0 17.4
R24922 net3_ota.n108 net3_ota.n107 9.3
R24923 net3_ota.n204 net3_ota.n203 9.3
R24924 net3_ota.n340 net3_ota.n339 9.3
R24925 net3_ota.n436 net3_ota.n435 9.3
R24926 net3_ota.n225 net3_ota.n224 8.886
R24927 net3_ota.n460 net3_ota.n459 8.886
R24928 net3_ota.n39 net3_ota.n38 8.5
R24929 net3_ota.n3 net3_ota.n2 8.282
R24930 net3_ota.n224 net3_ota.t1 7.141
R24931 net3_ota.n459 net3_ota.t2 7.141
R24932 net3_ota.n54 net3_ota.n53 7.033
R24933 net3_ota.n286 net3_ota.n285 7.033
R24934 net3_ota.n263 net3_ota.n262 7.03
R24935 net3_ota.n495 net3_ota.n494 7.03
R24936 net3_ota.n510 net3_ota.n509 6.212
R24937 net3_ota.n4 net3_ota.n3 4.5
R24938 net3_ota.n34 net3_ota.n33 4.5
R24939 net3_ota.n41 net3_ota.n40 4.5
R24940 net3_ota.n10 net3_ota.n9 4.5
R24941 net3_ota.n91 net3_ota.n90 4.5
R24942 net3_ota.n207 net3_ota.n199 4.5
R24943 net3_ota.n232 net3_ota.n227 4.5
R24944 net3_ota.n186 net3_ota.n185 4.5
R24945 net3_ota.n160 net3_ota.n158 4.5
R24946 net3_ota.n171 net3_ota.n166 4.5
R24947 net3_ota.n150 net3_ota.n147 4.5
R24948 net3_ota.n129 net3_ota.n128 4.5
R24949 net3_ota.n140 net3_ota.n135 4.5
R24950 net3_ota.n114 net3_ota.n113 4.5
R24951 net3_ota.n73 net3_ota.n72 4.5
R24952 net3_ota.n251 net3_ota.n250 4.5
R24953 net3_ota.n323 net3_ota.n322 4.5
R24954 net3_ota.n439 net3_ota.n431 4.5
R24955 net3_ota.n418 net3_ota.n417 4.5
R24956 net3_ota.n392 net3_ota.n390 4.5
R24957 net3_ota.n403 net3_ota.n398 4.5
R24958 net3_ota.n382 net3_ota.n379 4.5
R24959 net3_ota.n361 net3_ota.n360 4.5
R24960 net3_ota.n372 net3_ota.n367 4.5
R24961 net3_ota.n346 net3_ota.n345 4.5
R24962 net3_ota.n305 net3_ota.n304 4.5
R24963 net3_ota.n463 net3_ota.n462 4.5
R24964 net3_ota.n482 net3_ota.n481 4.5
R24965 net3_ota.n40 net3_ota.n37 4.141
R24966 net3_ota.n227 net3_ota.n223 4.141
R24967 net3_ota.n166 net3_ota.n165 4.141
R24968 net3_ota.n128 net3_ota.n127 4.141
R24969 net3_ota.n72 net3_ota.n71 4.141
R24970 net3_ota.n462 net3_ota.n458 4.141
R24971 net3_ota.n398 net3_ota.n397 4.141
R24972 net3_ota.n360 net3_ota.n359 4.141
R24973 net3_ota.n304 net3_ota.n303 4.141
R24974 net3_ota.n9 net3_ota.n8 3.764
R24975 net3_ota.n3 net3_ota.n1 3.764
R24976 net3_ota.n185 net3_ota.n184 3.764
R24977 net3_ota.n113 net3_ota.n112 3.764
R24978 net3_ota.n417 net3_ota.n416 3.764
R24979 net3_ota.n345 net3_ota.n344 3.764
R24980 net3_ota.n33 net3_ota.n32 3.388
R24981 net3_ota.n250 net3_ota.n247 3.388
R24982 net3_ota.n199 net3_ota.n196 3.388
R24983 net3_ota.n135 net3_ota.n133 3.388
R24984 net3_ota.n90 net3_ota.n89 3.388
R24985 net3_ota.n481 net3_ota.n478 3.388
R24986 net3_ota.n431 net3_ota.n428 3.388
R24987 net3_ota.n367 net3_ota.n365 3.388
R24988 net3_ota.n322 net3_ota.n321 3.388
R24989 net3_ota.n250 net3_ota.n249 3.011
R24990 net3_ota.n199 net3_ota.n198 3.011
R24991 net3_ota.n203 net3_ota.n202 3.011
R24992 net3_ota.n158 net3_ota.n156 3.011
R24993 net3_ota.n135 net3_ota.n134 3.011
R24994 net3_ota.n90 net3_ota.n88 3.011
R24995 net3_ota.n481 net3_ota.n480 3.011
R24996 net3_ota.n431 net3_ota.n430 3.011
R24997 net3_ota.n435 net3_ota.n434 3.011
R24998 net3_ota.n390 net3_ota.n388 3.011
R24999 net3_ota.n367 net3_ota.n366 3.011
R25000 net3_ota.n322 net3_ota.n320 3.011
R25001 net3_ota.n9 net3_ota.n7 2.635
R25002 net3_ota.n185 net3_ota.n182 2.635
R25003 net3_ota.n147 net3_ota.n146 2.635
R25004 net3_ota.n107 net3_ota.n106 2.635
R25005 net3_ota.n113 net3_ota.n111 2.635
R25006 net3_ota.n417 net3_ota.n414 2.635
R25007 net3_ota.n379 net3_ota.n378 2.635
R25008 net3_ota.n339 net3_ota.n338 2.635
R25009 net3_ota.n345 net3_ota.n343 2.635
R25010 net3_ota net3_ota.n44 2.569
R25011 net3_ota.n40 net3_ota.n39 2.258
R25012 net3_ota.n227 net3_ota.n226 2.258
R25013 net3_ota.n72 net3_ota.n70 2.258
R25014 net3_ota.n462 net3_ota.n461 2.258
R25015 net3_ota.n304 net3_ota.n302 2.258
R25016 net3_ota net3_ota.n510 1.814
R25017 net3_ota.n98 net3_ota.n54 1.508
R25018 net3_ota.n330 net3_ota.n286 1.508
R25019 net3_ota.n158 net3_ota.n157 1.505
R25020 net3_ota.n390 net3_ota.n389 1.505
R25021 net3_ota.n92 net3_ota.n91 1.5
R25022 net3_ota.n269 net3_ota.n268 1.5
R25023 net3_ota.n233 net3_ota.n232 1.5
R25024 net3_ota.n208 net3_ota.n207 1.5
R25025 net3_ota.n187 net3_ota.n186 1.5
R25026 net3_ota.n161 net3_ota.n160 1.5
R25027 net3_ota.n172 net3_ota.n171 1.5
R25028 net3_ota.n151 net3_ota.n150 1.5
R25029 net3_ota.n130 net3_ota.n129 1.5
R25030 net3_ota.n141 net3_ota.n140 1.5
R25031 net3_ota.n115 net3_ota.n114 1.5
R25032 net3_ota.n74 net3_ota.n73 1.5
R25033 net3_ota.n252 net3_ota.n251 1.5
R25034 net3_ota.n324 net3_ota.n323 1.5
R25035 net3_ota.n501 net3_ota.n500 1.5
R25036 net3_ota.n440 net3_ota.n439 1.5
R25037 net3_ota.n419 net3_ota.n418 1.5
R25038 net3_ota.n393 net3_ota.n392 1.5
R25039 net3_ota.n404 net3_ota.n403 1.5
R25040 net3_ota.n383 net3_ota.n382 1.5
R25041 net3_ota.n362 net3_ota.n361 1.5
R25042 net3_ota.n373 net3_ota.n372 1.5
R25043 net3_ota.n347 net3_ota.n346 1.5
R25044 net3_ota.n306 net3_ota.n305 1.5
R25045 net3_ota.n464 net3_ota.n463 1.5
R25046 net3_ota.n483 net3_ota.n482 1.5
R25047 net3_ota.n509 net3_ota.n508 1.448
R25048 net3_ota.n43 net3_ota.n42 1.384
R25049 net3_ota.n12 net3_ota.n11 1.384
R25050 net3_ota.n509 net3_ota.n276 1.366
R25051 net3_ota.n13 net3_ota.n12 1.146
R25052 net3_ota.n44 net3_ota.n43 1.137
R25053 net3_ota.n23 net3_ota.n22 1.137
R25054 net3_ota.n19 net3_ota.n18 1.137
R25055 net3_ota.n117 net3_ota.n116 1.137
R25056 net3_ota.n124 net3_ota.n123 1.137
R25057 net3_ota.n216 net3_ota.n215 1.137
R25058 net3_ota.n274 net3_ota.n273 1.137
R25059 net3_ota.n237 net3_ota.n236 1.137
R25060 net3_ota.n191 net3_ota.n190 1.137
R25061 net3_ota.n212 net3_ota.n211 1.137
R25062 net3_ota.n174 net3_ota.n173 1.137
R25063 net3_ota.n155 net3_ota.n154 1.137
R25064 net3_ota.n258 net3_ota.n257 1.137
R25065 net3_ota.n490 net3_ota.n489 1.137
R25066 net3_ota.n349 net3_ota.n348 1.137
R25067 net3_ota.n356 net3_ota.n355 1.137
R25068 net3_ota.n448 net3_ota.n447 1.137
R25069 net3_ota.n506 net3_ota.n505 1.137
R25070 net3_ota.n423 net3_ota.n422 1.137
R25071 net3_ota.n444 net3_ota.n443 1.137
R25072 net3_ota.n406 net3_ota.n405 1.137
R25073 net3_ota.n387 net3_ota.n386 1.137
R25074 net3_ota.n468 net3_ota.n467 1.137
R25075 net3_ota.n147 net3_ota.n145 1.129
R25076 net3_ota.n379 net3_ota.n377 1.129
R25077 net3_ota.n99 net3_ota.n98 0.72
R25078 net3_ota.n331 net3_ota.n330 0.72
R25079 net3_ota.n262 net3_ota.n261 0.155
R25080 net3_ota.n53 net3_ota.n52 0.155
R25081 net3_ota.n494 net3_ota.n493 0.155
R25082 net3_ota.n285 net3_ota.n284 0.155
R25083 net3_ota.n249 net3_ota.n248 0.144
R25084 net3_ota.n480 net3_ota.n479 0.144
R25085 net3_ota.n88 net3_ota.n87 0.144
R25086 net3_ota.n320 net3_ota.n319 0.144
R25087 net3_ota.n226 net3_ota.n225 0.133
R25088 net3_ota.n461 net3_ota.n460 0.133
R25089 net3_ota.n70 net3_ota.n69 0.132
R25090 net3_ota.n302 net3_ota.n301 0.132
R25091 net3_ota.n230 net3_ota.n229 0.056
R25092 net3_ota.n456 net3_ota.n455 0.056
R25093 net3_ota.n84 net3_ota.n83 0.047
R25094 net3_ota.n316 net3_ota.n315 0.047
R25095 net3_ota.n233 net3_ota.n219 0.045
R25096 net3_ota.n189 net3_ota.n188 0.045
R25097 net3_ota.n173 net3_ota.n172 0.045
R25098 net3_ota.n421 net3_ota.n420 0.045
R25099 net3_ota.n405 net3_ota.n404 0.045
R25100 net3_ota.n204 net3_ota.n201 0.043
R25101 net3_ota.n154 net3_ota.n130 0.043
R25102 net3_ota.n436 net3_ota.n433 0.043
R25103 net3_ota.n386 net3_ota.n362 0.043
R25104 net3_ota.n252 net3_ota.n240 0.041
R25105 net3_ota.n75 net3_ota.n74 0.041
R25106 net3_ota.n483 net3_ota.n471 0.041
R25107 net3_ota.n307 net3_ota.n306 0.041
R25108 net3_ota.n160 net3_ota.n159 0.039
R25109 net3_ota.n273 net3_ota.n272 0.039
R25110 net3_ota.n93 net3_ota.n92 0.039
R25111 net3_ota.n392 net3_ota.n391 0.039
R25112 net3_ota.n505 net3_ota.n504 0.039
R25113 net3_ota.n325 net3_ota.n324 0.039
R25114 net3_ota.n150 net3_ota.n144 0.037
R25115 net3_ota.n66 net3_ota.n65 0.037
R25116 net3_ota.n97 net3_ota.n96 0.037
R25117 net3_ota.n274 net3_ota.n258 0.037
R25118 net3_ota.n174 net3_ota.n155 0.037
R25119 net3_ota.n382 net3_ota.n376 0.037
R25120 net3_ota.n298 net3_ota.n297 0.037
R25121 net3_ota.n329 net3_ota.n328 0.037
R25122 net3_ota.n506 net3_ota.n490 0.037
R25123 net3_ota.n406 net3_ota.n387 0.037
R25124 net3_ota.n30 net3_ota.n29 0.035
R25125 net3_ota.n31 net3_ota.n30 0.035
R25126 net3_ota.n22 net3_ota.n20 0.035
R25127 net3_ota.n138 net3_ota.n137 0.034
R25128 net3_ota.n48 net3_ota.n47 0.034
R25129 net3_ota.n271 net3_ota.n270 0.034
R25130 net3_ota.n164 net3_ota.n163 0.034
R25131 net3_ota.n95 net3_ota.n94 0.034
R25132 net3_ota.n370 net3_ota.n369 0.034
R25133 net3_ota.n280 net3_ota.n279 0.034
R25134 net3_ota.n503 net3_ota.n502 0.034
R25135 net3_ota.n396 net3_ota.n395 0.034
R25136 net3_ota.n327 net3_ota.n326 0.034
R25137 net3_ota.n260 net3_ota.n259 0.032
R25138 net3_ota.n152 net3_ota.n151 0.032
R25139 net3_ota.n142 net3_ota.n141 0.032
R25140 net3_ota.n492 net3_ota.n491 0.032
R25141 net3_ota.n384 net3_ota.n383 0.032
R25142 net3_ota.n374 net3_ota.n373 0.032
R25143 net3_ota.n50 net3_ota.n49 0.03
R25144 net3_ota.n254 net3_ota.n253 0.03
R25145 net3_ota.n187 net3_ota.n177 0.03
R25146 net3_ota.n162 net3_ota.n161 0.03
R25147 net3_ota.n282 net3_ota.n281 0.03
R25148 net3_ota.n486 net3_ota.n485 0.03
R25149 net3_ota.n419 net3_ota.n409 0.03
R25150 net3_ota.n394 net3_ota.n393 0.03
R25151 net3_ota.n266 net3_ota.n265 0.028
R25152 net3_ota.n77 net3_ota.n76 0.028
R25153 net3_ota.n498 net3_ota.n497 0.028
R25154 net3_ota.n309 net3_ota.n308 0.028
R25155 net3_ota.n23 net3_ota.n19 0.027
R25156 net3_ota.n64 net3_ota.n63 0.026
R25157 net3_ota.n85 net3_ota.n84 0.026
R25158 net3_ota.n256 net3_ota.n255 0.026
R25159 net3_ota.n56 net3_ota.n55 0.026
R25160 net3_ota.n296 net3_ota.n295 0.026
R25161 net3_ota.n317 net3_ota.n316 0.026
R25162 net3_ota.n488 net3_ota.n487 0.026
R25163 net3_ota.n288 net3_ota.n287 0.026
R25164 net3_ota.n243 net3_ota.n242 0.024
R25165 net3_ota.n245 net3_ota.n244 0.024
R25166 net3_ota.n222 net3_ota.n221 0.024
R25167 net3_ota.n236 net3_ota.n235 0.024
R25168 net3_ota.n214 net3_ota.n213 0.024
R25169 net3_ota.n211 net3_ota.n210 0.024
R25170 net3_ota.n123 net3_ota.n122 0.024
R25171 net3_ota.n58 net3_ota.n57 0.024
R25172 net3_ota.n61 net3_ota.n60 0.024
R25173 net3_ota.n79 net3_ota.n78 0.024
R25174 net3_ota.n474 net3_ota.n473 0.024
R25175 net3_ota.n476 net3_ota.n475 0.024
R25176 net3_ota.n453 net3_ota.n452 0.024
R25177 net3_ota.n467 net3_ota.n466 0.024
R25178 net3_ota.n446 net3_ota.n445 0.024
R25179 net3_ota.n443 net3_ota.n442 0.024
R25180 net3_ota.n355 net3_ota.n354 0.024
R25181 net3_ota.n290 net3_ota.n289 0.024
R25182 net3_ota.n293 net3_ota.n292 0.024
R25183 net3_ota.n311 net3_ota.n310 0.024
R25184 net3_ota.n198 net3_ota.n197 0.024
R25185 net3_ota.n111 net3_ota.n110 0.024
R25186 net3_ota.n430 net3_ota.n429 0.024
R25187 net3_ota.n343 net3_ota.n342 0.024
R25188 net3_ota.n238 net3_ota.n237 0.023
R25189 net3_ota.n191 net3_ota.n176 0.023
R25190 net3_ota.n125 net3_ota.n124 0.023
R25191 net3_ota.n102 net3_ota.n101 0.023
R25192 net3_ota.n469 net3_ota.n468 0.023
R25193 net3_ota.n423 net3_ota.n408 0.023
R25194 net3_ota.n357 net3_ota.n356 0.023
R25195 net3_ota.n334 net3_ota.n333 0.023
R25196 net3_ota.n67 net3_ota.n66 0.022
R25197 net3_ota.n46 net3_ota.n45 0.022
R25198 net3_ota.n299 net3_ota.n298 0.022
R25199 net3_ota.n278 net3_ota.n277 0.022
R25200 net3_ota.n41 net3_ota.n36 0.02
R25201 net3_ota.n232 net3_ota.n222 0.02
R25202 net3_ota.n82 net3_ota.n81 0.02
R25203 net3_ota.n216 net3_ota.n212 0.02
R25204 net3_ota.n117 net3_ota.n105 0.02
R25205 net3_ota.n463 net3_ota.n453 0.02
R25206 net3_ota.n314 net3_ota.n313 0.02
R25207 net3_ota.n448 net3_ota.n444 0.02
R25208 net3_ota.n349 net3_ota.n337 0.02
R25209 net3_ota.n10 net3_ota.n6 0.018
R25210 net3_ota.n5 net3_ota.n4 0.018
R25211 net3_ota.n17 net3_ota.n16 0.018
R25212 net3_ota.n186 net3_ota.n181 0.018
R25213 net3_ota.n109 net3_ota.n108 0.018
R25214 net3_ota.n78 net3_ota.n77 0.018
R25215 net3_ota.n418 net3_ota.n413 0.018
R25216 net3_ota.n341 net3_ota.n340 0.018
R25217 net3_ota.n310 net3_ota.n309 0.018
R25218 net3_ota.n35 net3_ota.n34 0.017
R25219 net3_ota.n251 net3_ota.n243 0.017
R25220 net3_ota.n207 net3_ota.n195 0.017
R25221 net3_ota.n205 net3_ota.n204 0.017
R25222 net3_ota.n170 net3_ota.n169 0.017
R25223 net3_ota.n255 net3_ota.n254 0.017
R25224 net3_ota.n482 net3_ota.n474 0.017
R25225 net3_ota.n439 net3_ota.n427 0.017
R25226 net3_ota.n437 net3_ota.n436 0.017
R25227 net3_ota.n402 net3_ota.n401 0.017
R25228 net3_ota.n487 net3_ota.n486 0.017
R25229 net3_ota.n12 net3_ota.n0 0.015
R25230 net3_ota.n16 net3_ota.n15 0.015
R25231 net3_ota.n27 net3_ota.n26 0.015
R25232 net3_ota.n168 net3_ota.n167 0.015
R25233 net3_ota.n235 net3_ota.n234 0.015
R25234 net3_ota.n210 net3_ota.n209 0.015
R25235 net3_ota.n122 net3_ota.n121 0.015
R25236 net3_ota.n400 net3_ota.n399 0.015
R25237 net3_ota.n466 net3_ota.n465 0.015
R25238 net3_ota.n442 net3_ota.n441 0.015
R25239 net3_ota.n354 net3_ota.n353 0.015
R25240 net3_ota.n11 net3_ota.n10 0.013
R25241 net3_ota.n43 net3_ota.n28 0.013
R25242 net3_ota.n150 net3_ota.n149 0.013
R25243 net3_ota.n149 net3_ota.n148 0.013
R25244 net3_ota.n139 net3_ota.n138 0.013
R25245 net3_ota.n114 net3_ota.n109 0.013
R25246 net3_ota.n116 net3_ota.n115 0.013
R25247 net3_ota.n59 net3_ota.n58 0.013
R25248 net3_ota.n382 net3_ota.n381 0.013
R25249 net3_ota.n381 net3_ota.n380 0.013
R25250 net3_ota.n371 net3_ota.n370 0.013
R25251 net3_ota.n346 net3_ota.n341 0.013
R25252 net3_ota.n348 net3_ota.n347 0.013
R25253 net3_ota.n291 net3_ota.n290 0.013
R25254 net3_ota.n184 net3_ota.n183 0.012
R25255 net3_ota.n133 net3_ota.n132 0.012
R25256 net3_ota.n416 net3_ota.n415 0.012
R25257 net3_ota.n365 net3_ota.n364 0.012
R25258 net3_ota.n276 net3_ota.n275 0.012
R25259 net3_ota.n239 net3_ota.n238 0.012
R25260 net3_ota.n176 net3_ota.n175 0.012
R25261 net3_ota.n126 net3_ota.n125 0.012
R25262 net3_ota.n101 net3_ota.n100 0.012
R25263 net3_ota.n508 net3_ota.n507 0.012
R25264 net3_ota.n470 net3_ota.n469 0.012
R25265 net3_ota.n408 net3_ota.n407 0.012
R25266 net3_ota.n358 net3_ota.n357 0.012
R25267 net3_ota.n333 net3_ota.n332 0.012
R25268 net3_ota.n42 net3_ota.n41 0.011
R25269 net3_ota.n28 net3_ota.n27 0.011
R25270 net3_ota.n267 net3_ota.n266 0.011
R25271 net3_ota.n246 net3_ota.n245 0.011
R25272 net3_ota.n229 net3_ota.n228 0.011
R25273 net3_ota.n207 net3_ota.n206 0.011
R25274 net3_ota.n49 net3_ota.n48 0.011
R25275 net3_ota.n54 net3_ota.n51 0.011
R25276 net3_ota.n215 net3_ota.n214 0.011
R25277 net3_ota.n211 net3_ota.n208 0.011
R25278 net3_ota.n151 net3_ota.n142 0.011
R25279 net3_ota.n96 net3_ota.n95 0.011
R25280 net3_ota.n499 net3_ota.n498 0.011
R25281 net3_ota.n477 net3_ota.n476 0.011
R25282 net3_ota.n455 net3_ota.n454 0.011
R25283 net3_ota.n439 net3_ota.n438 0.011
R25284 net3_ota.n281 net3_ota.n280 0.011
R25285 net3_ota.n286 net3_ota.n283 0.011
R25286 net3_ota.n447 net3_ota.n446 0.011
R25287 net3_ota.n443 net3_ota.n440 0.011
R25288 net3_ota.n383 net3_ota.n374 0.011
R25289 net3_ota.n328 net3_ota.n327 0.011
R25290 net3_ota.n19 net3_ota.n14 0.009
R25291 net3_ota.n24 net3_ota.n23 0.009
R25292 net3_ota.n44 net3_ota.n25 0.009
R25293 net3_ota.n265 net3_ota.n264 0.009
R25294 net3_ota.n179 net3_ota.n178 0.009
R25295 net3_ota.n181 net3_ota.n180 0.009
R25296 net3_ota.n65 net3_ota.n64 0.009
R25297 net3_ota.n272 net3_ota.n271 0.009
R25298 net3_ota.n257 net3_ota.n256 0.009
R25299 net3_ota.n173 net3_ota.n162 0.009
R25300 net3_ota.n57 net3_ota.n56 0.009
R25301 net3_ota.n80 net3_ota.n79 0.009
R25302 net3_ota.n497 net3_ota.n496 0.009
R25303 net3_ota.n411 net3_ota.n410 0.009
R25304 net3_ota.n413 net3_ota.n412 0.009
R25305 net3_ota.n297 net3_ota.n296 0.009
R25306 net3_ota.n504 net3_ota.n503 0.009
R25307 net3_ota.n489 net3_ota.n488 0.009
R25308 net3_ota.n405 net3_ota.n394 0.009
R25309 net3_ota.n289 net3_ota.n288 0.009
R25310 net3_ota.n312 net3_ota.n311 0.009
R25311 net3_ota.n34 net3_ota.n31 0.007
R25312 net3_ota.n22 net3_ota.n21 0.007
R25313 net3_ota.n268 net3_ota.n267 0.007
R25314 net3_ota.n231 net3_ota.n230 0.007
R25315 net3_ota.n195 net3_ota.n194 0.007
R25316 net3_ota.n73 net3_ota.n68 0.007
R25317 net3_ota.n86 net3_ota.n85 0.007
R25318 net3_ota.n91 net3_ota.n86 0.007
R25319 net3_ota.n51 net3_ota.n50 0.007
R25320 net3_ota.n273 net3_ota.n269 0.007
R25321 net3_ota.n74 net3_ota.n61 0.007
R25322 net3_ota.n92 net3_ota.n80 0.007
R25323 net3_ota.n237 net3_ota.n218 0.007
R25324 net3_ota.n217 net3_ota.n216 0.007
R25325 net3_ota.n212 net3_ota.n193 0.007
R25326 net3_ota.n192 net3_ota.n191 0.007
R25327 net3_ota.n124 net3_ota.n119 0.007
R25328 net3_ota.n118 net3_ota.n117 0.007
R25329 net3_ota.n105 net3_ota.n104 0.007
R25330 net3_ota.n103 net3_ota.n102 0.007
R25331 net3_ota.n500 net3_ota.n499 0.007
R25332 net3_ota.n457 net3_ota.n456 0.007
R25333 net3_ota.n427 net3_ota.n426 0.007
R25334 net3_ota.n305 net3_ota.n300 0.007
R25335 net3_ota.n318 net3_ota.n317 0.007
R25336 net3_ota.n323 net3_ota.n318 0.007
R25337 net3_ota.n283 net3_ota.n282 0.007
R25338 net3_ota.n505 net3_ota.n501 0.007
R25339 net3_ota.n306 net3_ota.n293 0.007
R25340 net3_ota.n324 net3_ota.n312 0.007
R25341 net3_ota.n468 net3_ota.n450 0.007
R25342 net3_ota.n449 net3_ota.n448 0.007
R25343 net3_ota.n444 net3_ota.n425 0.007
R25344 net3_ota.n424 net3_ota.n423 0.007
R25345 net3_ota.n356 net3_ota.n351 0.007
R25346 net3_ota.n350 net3_ota.n349 0.007
R25347 net3_ota.n337 net3_ota.n336 0.007
R25348 net3_ota.n335 net3_ota.n334 0.007
R25349 net3_ota.n6 net3_ota.n5 0.005
R25350 net3_ota.n36 net3_ota.n35 0.005
R25351 net3_ota.n18 net3_ota.n17 0.005
R25352 net3_ota.n14 net3_ota.n13 0.005
R25353 net3_ota.n25 net3_ota.n24 0.005
R25354 net3_ota.n83 net3_ota.n82 0.005
R25355 net3_ota.n153 net3_ota.n152 0.005
R25356 net3_ota.n76 net3_ota.n75 0.005
R25357 net3_ota.n315 net3_ota.n314 0.005
R25358 net3_ota.n385 net3_ota.n384 0.005
R25359 net3_ota.n308 net3_ota.n307 0.005
R25360 net3_ota.n98 net3_ota.n97 0.004
R25361 net3_ota.n330 net3_ota.n329 0.004
R25362 net3_ota.n268 net3_ota.n263 0.004
R25363 net3_ota.n500 net3_ota.n495 0.004
R25364 net3_ota.n218 net3_ota.n217 0.004
R25365 net3_ota.n193 net3_ota.n192 0.004
R25366 net3_ota.n119 net3_ota.n118 0.004
R25367 net3_ota.n104 net3_ota.n103 0.004
R25368 net3_ota.n450 net3_ota.n449 0.004
R25369 net3_ota.n425 net3_ota.n424 0.004
R25370 net3_ota.n351 net3_ota.n350 0.004
R25371 net3_ota.n336 net3_ota.n335 0.004
R25372 net3_ota.n242 net3_ota.n241 0.003
R25373 net3_ota.n251 net3_ota.n246 0.003
R25374 net3_ota.n221 net3_ota.n220 0.003
R25375 net3_ota.n232 net3_ota.n231 0.003
R25376 net3_ota.n206 net3_ota.n205 0.003
R25377 net3_ota.n201 net3_ota.n200 0.003
R25378 net3_ota.n186 net3_ota.n179 0.003
R25379 net3_ota.n171 net3_ota.n170 0.003
R25380 net3_ota.n144 net3_ota.n143 0.003
R25381 net3_ota.n63 net3_ota.n62 0.003
R25382 net3_ota.n68 net3_ota.n67 0.003
R25383 net3_ota.n257 net3_ota.n252 0.003
R25384 net3_ota.n236 net3_ota.n233 0.003
R25385 net3_ota.n190 net3_ota.n189 0.003
R25386 net3_ota.n188 net3_ota.n187 0.003
R25387 net3_ota.n172 net3_ota.n164 0.003
R25388 net3_ota.n154 net3_ota.n153 0.003
R25389 net3_ota.n473 net3_ota.n472 0.003
R25390 net3_ota.n482 net3_ota.n477 0.003
R25391 net3_ota.n452 net3_ota.n451 0.003
R25392 net3_ota.n463 net3_ota.n457 0.003
R25393 net3_ota.n438 net3_ota.n437 0.003
R25394 net3_ota.n433 net3_ota.n432 0.003
R25395 net3_ota.n418 net3_ota.n411 0.003
R25396 net3_ota.n403 net3_ota.n402 0.003
R25397 net3_ota.n376 net3_ota.n375 0.003
R25398 net3_ota.n295 net3_ota.n294 0.003
R25399 net3_ota.n300 net3_ota.n299 0.003
R25400 net3_ota.n489 net3_ota.n483 0.003
R25401 net3_ota.n485 net3_ota.n484 0.003
R25402 net3_ota.n467 net3_ota.n464 0.003
R25403 net3_ota.n422 net3_ota.n421 0.003
R25404 net3_ota.n420 net3_ota.n419 0.003
R25405 net3_ota.n404 net3_ota.n396 0.003
R25406 net3_ota.n386 net3_ota.n385 0.003
R25407 net3_ota.n275 net3_ota.n274 0.002
R25408 net3_ota.n258 net3_ota.n239 0.002
R25409 net3_ota.n175 net3_ota.n174 0.002
R25410 net3_ota.n155 net3_ota.n126 0.002
R25411 net3_ota.n100 net3_ota.n99 0.002
R25412 net3_ota.n507 net3_ota.n506 0.002
R25413 net3_ota.n490 net3_ota.n470 0.002
R25414 net3_ota.n407 net3_ota.n406 0.002
R25415 net3_ota.n387 net3_ota.n358 0.002
R25416 net3_ota.n332 net3_ota.n331 0.002
R25417 net3_ota.n169 net3_ota.n168 0.001
R25418 net3_ota.n140 net3_ota.n139 0.001
R25419 net3_ota.n137 net3_ota.n136 0.001
R25420 net3_ota.n47 net3_ota.n46 0.001
R25421 net3_ota.n269 net3_ota.n260 0.001
R25422 net3_ota.n141 net3_ota.n131 0.001
R25423 net3_ota.n123 net3_ota.n120 0.001
R25424 net3_ota.n60 net3_ota.n59 0.001
R25425 net3_ota.n94 net3_ota.n93 0.001
R25426 net3_ota.n401 net3_ota.n400 0.001
R25427 net3_ota.n372 net3_ota.n371 0.001
R25428 net3_ota.n369 net3_ota.n368 0.001
R25429 net3_ota.n279 net3_ota.n278 0.001
R25430 net3_ota.n501 net3_ota.n492 0.001
R25431 net3_ota.n373 net3_ota.n363 0.001
R25432 net3_ota.n355 net3_ota.n352 0.001
R25433 net3_ota.n292 net3_ota.n291 0.001
R25434 net3_ota.n326 net3_ota.n325 0.001
R25435 Nbais.n256 Nbais.n255 175.251
R25436 Nbais.n179 Nbais.n178 175.251
R25437 Nbais.n86 Nbais.n85 175.251
R25438 Nbais.n2 Nbais.t0 124.695
R25439 Nbais.n255 Nbais.t3 122.709
R25440 Nbais.n178 Nbais.t1 122.709
R25441 Nbais.n85 Nbais.t2 122.709
R25442 Nbais.n294 Nbais.t11 117.491
R25443 Nbais.n307 Nbais.t13 117.249
R25444 Nbais.n306 Nbais.t4 117.249
R25445 Nbais.n305 Nbais.t12 117.249
R25446 Nbais.n304 Nbais.t5 117.249
R25447 Nbais.n303 Nbais.t14 117.249
R25448 Nbais.n302 Nbais.t6 117.249
R25449 Nbais.n301 Nbais.t7 117.249
R25450 Nbais.n300 Nbais.t16 117.249
R25451 Nbais.n299 Nbais.t8 117.249
R25452 Nbais.n298 Nbais.t15 117.249
R25453 Nbais.n297 Nbais.t10 117.249
R25454 Nbais.n296 Nbais.t17 117.249
R25455 Nbais.n295 Nbais.t9 117.249
R25456 Nbais.n294 Nbais.t18 117.249
R25457 Nbais.n1 Nbais.n0 92.5
R25458 Nbais.n11 Nbais.n10 31.034
R25459 Nbais.n2 Nbais.n1 15.431
R25460 Nbais.n293 Nbais.n19 11.676
R25461 Nbais.n15 Nbais.n14 9.3
R25462 Nbais.n6 Nbais.n5 9.3
R25463 Nbais.n4 Nbais.n3 9.3
R25464 Nbais.n13 Nbais.n12 9.3
R25465 Nbais.n12 Nbais.n11 9.3
R25466 Nbais.n17 Nbais.n16 9.3
R25467 Nbais.n19 Nbais.n18 9.3
R25468 Nbais.n63 Nbais.n62 9.3
R25469 Nbais.n239 Nbais.n238 9.013
R25470 Nbais.n199 Nbais.n198 9.013
R25471 Nbais.n113 Nbais.n112 9.013
R25472 Nbais.n229 Nbais.n228 9.013
R25473 Nbais.n98 Nbais.n97 9.013
R25474 Nbais.n34 Nbais.n33 9.013
R25475 Nbais.n257 Nbais.n256 6.413
R25476 Nbais.n180 Nbais.n179 6.413
R25477 Nbais.n87 Nbais.n86 6.413
R25478 Nbais.n12 Nbais.n8 5.647
R25479 Nbais.n183 Nbais.n182 4.5
R25480 Nbais.n165 Nbais.n155 4.5
R25481 Nbais.n170 Nbais.n151 4.5
R25482 Nbais.n167 Nbais.n153 4.5
R25483 Nbais.n162 Nbais.n159 4.5
R25484 Nbais.n220 Nbais.n218 4.5
R25485 Nbais.n92 Nbais.n89 4.5
R25486 Nbais.n49 Nbais.n48 4.5
R25487 Nbais.n40 Nbais.n39 4.5
R25488 Nbais.n45 Nbais.n44 4.5
R25489 Nbais.n55 Nbais.n54 4.5
R25490 Nbais.n66 Nbais.n65 4.5
R25491 Nbais.n260 Nbais.n259 4.5
R25492 Nbais.n145 Nbais.n142 4.5
R25493 Nbais.n270 Nbais.n269 4.5
R25494 Nbais.n287 Nbais.n285 4.5
R25495 Nbais.n139 Nbais.n136 4.5
R25496 Nbais.n128 Nbais.n125 4.5
R25497 Nbais.n10 Nbais.n9 4.137
R25498 Nbais.n114 Nbais.n113 3.992
R25499 Nbais.n230 Nbais.n229 3.992
R25500 Nbais.n240 Nbais.n239 3.882
R25501 Nbais.n99 Nbais.n98 3.882
R25502 Nbais.n70 Nbais.n34 2.792
R25503 Nbais.n256 Nbais.n254 2.787
R25504 Nbais.n179 Nbais.n177 2.787
R25505 Nbais.n200 Nbais.n199 2.738
R25506 Nbais.n257 Nbais.n253 2.695
R25507 Nbais.n180 Nbais.n176 2.695
R25508 Nbais.n63 Nbais.n61 2.695
R25509 Nbais.n285 Nbais.n284 2.656
R25510 Nbais.n32 Nbais.n31 2.535
R25511 Nbais.n197 Nbais.n196 2.415
R25512 Nbais.n268 Nbais.n267 2.082
R25513 Nbais.n135 Nbais.n134 2.082
R25514 Nbais.n258 Nbais.n257 2.082
R25515 Nbais.n124 Nbais.n123 2.082
R25516 Nbais.n150 Nbais.n149 2.082
R25517 Nbais.n158 Nbais.n157 2.082
R25518 Nbais.n181 Nbais.n180 2.082
R25519 Nbais.n217 Nbais.n216 2.082
R25520 Nbais.n88 Nbais.n87 2.082
R25521 Nbais.n38 Nbais.n37 2.082
R25522 Nbais.n53 Nbais.n52 2.082
R25523 Nbais.n64 Nbais.n63 2.082
R25524 Nbais.n4 Nbais.n2 1.57
R25525 Nbais.n288 Nbais.n287 1.501
R25526 Nbais.n146 Nbais.n145 1.501
R25527 Nbais.n221 Nbais.n220 1.5
R25528 Nbais.n232 Nbais.n231 1.5
R25529 Nbais.n93 Nbais.n92 1.5
R25530 Nbais.n104 Nbais.n103 1.5
R25531 Nbais.n271 Nbais.n270 1.5
R25532 Nbais.n140 Nbais.n139 1.5
R25533 Nbais.n261 Nbais.n260 1.5
R25534 Nbais.n129 Nbais.n128 1.5
R25535 Nbais.n116 Nbais.n115 1.5
R25536 Nbais.n244 Nbais.n243 1.5
R25537 Nbais.n258 Nbais.n252 1.449
R25538 Nbais.n181 Nbais.n175 1.449
R25539 Nbais.n88 Nbais.n84 1.449
R25540 Nbais.n239 Nbais.n237 1.328
R25541 Nbais.n124 Nbais.n122 1.328
R25542 Nbais.n199 Nbais.n197 1.328
R25543 Nbais.n217 Nbais.n215 1.328
R25544 Nbais.n98 Nbais.n96 1.328
R25545 Nbais.n64 Nbais.n60 1.328
R25546 Nbais.n285 Nbais.n274 1.207
R25547 Nbais.n136 Nbais.n135 1.207
R25548 Nbais.n113 Nbais.n111 1.207
R25549 Nbais.n153 Nbais.n152 1.207
R25550 Nbais.n159 Nbais.n158 1.207
R25551 Nbais.n229 Nbais.n227 1.207
R25552 Nbais.n44 Nbais.n43 1.207
R25553 Nbais.n54 Nbais.n53 1.207
R25554 Nbais.n34 Nbais.n32 1.207
R25555 Nbais.n292 Nbais.n291 1.137
R25556 Nbais.n289 Nbais.n20 1.137
R25557 Nbais.n269 Nbais.n268 1.086
R25558 Nbais.n142 Nbais.n141 1.086
R25559 Nbais.n151 Nbais.n150 1.086
R25560 Nbais.n155 Nbais.n154 1.086
R25561 Nbais.n39 Nbais.n38 1.086
R25562 Nbais.n48 Nbais.n47 1.086
R25563 Nbais.n71 Nbais.n70 0.935
R25564 Nbais.n201 Nbais.n200 0.935
R25565 Nbais Nbais.n307 0.821
R25566 Nbais.n8 Nbais.n7 0.752
R25567 Nbais.n125 Nbais.n124 0.724
R25568 Nbais.n218 Nbais.n217 0.724
R25569 Nbais.n65 Nbais.n64 0.724
R25570 Nbais.n259 Nbais.n258 0.603
R25571 Nbais.n182 Nbais.n181 0.603
R25572 Nbais.n89 Nbais.n88 0.603
R25573 Nbais.n134 Nbais.n133 0.557
R25574 Nbais.n157 Nbais.n156 0.557
R25575 Nbais.n293 Nbais.n292 0.438
R25576 Nbais Nbais.n293 0.313
R25577 Nbais.n106 Nbais.n105 0.245
R25578 Nbais.n234 Nbais.n233 0.245
R25579 Nbais.n307 Nbais.n306 0.242
R25580 Nbais.n306 Nbais.n305 0.242
R25581 Nbais.n305 Nbais.n304 0.242
R25582 Nbais.n304 Nbais.n303 0.242
R25583 Nbais.n303 Nbais.n302 0.242
R25584 Nbais.n302 Nbais.n301 0.242
R25585 Nbais.n301 Nbais.n300 0.242
R25586 Nbais.n300 Nbais.n299 0.242
R25587 Nbais.n299 Nbais.n298 0.242
R25588 Nbais.n298 Nbais.n297 0.242
R25589 Nbais.n297 Nbais.n296 0.242
R25590 Nbais.n296 Nbais.n295 0.242
R25591 Nbais.n295 Nbais.n294 0.242
R25592 Nbais.n15 Nbais.n13 0.144
R25593 Nbais.n186 Nbais.n185 0.048
R25594 Nbais.n173 Nbais.n172 0.048
R25595 Nbais.n225 Nbais.n224 0.048
R25596 Nbais.n101 Nbais.n100 0.048
R25597 Nbais.n58 Nbais.n57 0.048
R25598 Nbais.n69 Nbais.n68 0.048
R25599 Nbais.n166 Nbais.n165 0.044
R25600 Nbais.n49 Nbais.n46 0.044
R25601 Nbais.n287 Nbais.n286 0.042
R25602 Nbais.n167 Nbais.n166 0.042
R25603 Nbais.n46 Nbais.n45 0.042
R25604 Nbais.n13 Nbais.n6 0.04
R25605 Nbais.n270 Nbais.n266 0.036
R25606 Nbais.n171 Nbais.n170 0.036
R25607 Nbais.n40 Nbais.n36 0.036
R25608 Nbais.n19 Nbais.n17 0.035
R25609 Nbais.n139 Nbais.n138 0.034
R25610 Nbais.n162 Nbais.n161 0.034
R25611 Nbais.n56 Nbais.n55 0.034
R25612 Nbais.n200 Nbais.n186 0.031
R25613 Nbais.n70 Nbais.n69 0.031
R25614 Nbais.n260 Nbais.n249 0.028
R25615 Nbais.n184 Nbais.n183 0.028
R25616 Nbais.n92 Nbais.n83 0.028
R25617 Nbais.n128 Nbais.n127 0.026
R25618 Nbais.n220 Nbais.n219 0.026
R25619 Nbais.n204 Nbais.n203 0.026
R25620 Nbais.n221 Nbais.n212 0.026
R25621 Nbais.n232 Nbais.n223 0.026
R25622 Nbais.n67 Nbais.n66 0.026
R25623 Nbais.n104 Nbais.n95 0.026
R25624 Nbais.n93 Nbais.n82 0.026
R25625 Nbais.n74 Nbais.n73 0.026
R25626 Nbais.n251 Nbais.n250 0.023
R25627 Nbais.n127 Nbais.n126 0.023
R25628 Nbais.n174 Nbais.n173 0.023
R25629 Nbais.n91 Nbais.n90 0.023
R25630 Nbais.n68 Nbais.n67 0.023
R25631 Nbais.n242 Nbais.n241 0.021
R25632 Nbais.n249 Nbais.n248 0.021
R25633 Nbais.n121 Nbais.n120 0.021
R25634 Nbais.n185 Nbais.n184 0.021
R25635 Nbais.n214 Nbais.n213 0.021
R25636 Nbais.n102 Nbais.n101 0.021
R25637 Nbais.n59 Nbais.n58 0.021
R25638 Nbais.n287 Nbais.n273 0.019
R25639 Nbais.n110 Nbais.n109 0.019
R25640 Nbais.n168 Nbais.n167 0.019
R25641 Nbais.n163 Nbais.n162 0.019
R25642 Nbais.n226 Nbais.n225 0.019
R25643 Nbais.n45 Nbais.n42 0.019
R25644 Nbais.n55 Nbais.n51 0.019
R25645 Nbais.n145 Nbais.n144 0.017
R25646 Nbais.n170 Nbais.n169 0.017
R25647 Nbais.n165 Nbais.n164 0.017
R25648 Nbais.n41 Nbais.n40 0.017
R25649 Nbais.n50 Nbais.n49 0.017
R25650 Nbais.n138 Nbais.n137 0.015
R25651 Nbais.n161 Nbais.n160 0.015
R25652 Nbais.n57 Nbais.n56 0.015
R25653 Nbais.n263 Nbais.n262 0.015
R25654 Nbais.n107 Nbais.n106 0.015
R25655 Nbais.n235 Nbais.n234 0.015
R25656 Nbais.n207 Nbais.n206 0.014
R25657 Nbais.n208 Nbais.n207 0.014
R25658 Nbais.n209 Nbais.n208 0.014
R25659 Nbais.n210 Nbais.n209 0.014
R25660 Nbais.n80 Nbais.n79 0.014
R25661 Nbais.n79 Nbais.n78 0.014
R25662 Nbais.n78 Nbais.n77 0.014
R25663 Nbais.n77 Nbais.n76 0.014
R25664 Nbais.n131 Nbais.n130 0.014
R25665 Nbais.n146 Nbais.n140 0.013
R25666 Nbais.n288 Nbais.n271 0.013
R25667 Nbais.n289 Nbais.n146 0.013
R25668 Nbais.n289 Nbais.n288 0.013
R25669 Nbais.n266 Nbais.n265 0.013
R25670 Nbais.n115 Nbais.n110 0.013
R25671 Nbais.n172 Nbais.n171 0.013
R25672 Nbais.n231 Nbais.n226 0.013
R25673 Nbais.n36 Nbais.n35 0.013
R25674 Nbais.n117 Nbais.n116 0.013
R25675 Nbais.n206 Nbais.n205 0.012
R25676 Nbais.n81 Nbais.n80 0.012
R25677 Nbais.n245 Nbais.n244 0.012
R25678 Nbais.n246 Nbais.n245 0.012
R25679 Nbais.n118 Nbais.n117 0.012
R25680 Nbais.n105 Nbais.n104 0.012
R25681 Nbais.n233 Nbais.n232 0.011
R25682 Nbais.n243 Nbais.n242 0.011
R25683 Nbais.n128 Nbais.n121 0.011
R25684 Nbais.n220 Nbais.n214 0.011
R25685 Nbais.n211 Nbais.n210 0.011
R25686 Nbais.n103 Nbais.n102 0.011
R25687 Nbais.n66 Nbais.n59 0.011
R25688 Nbais.n76 Nbais.n75 0.011
R25689 Nbais.n271 Nbais.n264 0.011
R25690 Nbais.n17 Nbais.n15 0.01
R25691 Nbais.n262 Nbais.n261 0.01
R25692 Nbais.n140 Nbais.n132 0.01
R25693 Nbais.n130 Nbais.n129 0.01
R25694 Nbais.n260 Nbais.n251 0.009
R25695 Nbais.n183 Nbais.n174 0.009
R25696 Nbais.n203 Nbais.n202 0.009
R25697 Nbais.n92 Nbais.n91 0.009
R25698 Nbais.n94 Nbais.n93 0.009
R25699 Nbais.n261 Nbais.n247 0.009
R25700 Nbais.n222 Nbais.n221 0.008
R25701 Nbais.n73 Nbais.n72 0.008
R25702 Nbais.n129 Nbais.n119 0.008
R25703 Nbais.n273 Nbais.n272 0.007
R25704 Nbais.n144 Nbais.n143 0.007
R25705 Nbais.n169 Nbais.n168 0.007
R25706 Nbais.n164 Nbais.n163 0.007
R25707 Nbais.n202 Nbais.n201 0.007
R25708 Nbais.n223 Nbais.n222 0.007
R25709 Nbais.n42 Nbais.n41 0.007
R25710 Nbais.n51 Nbais.n50 0.007
R25711 Nbais.n95 Nbais.n94 0.007
R25712 Nbais.n72 Nbais.n71 0.007
R25713 Nbais.n119 Nbais.n118 0.007
R25714 Nbais.n103 Nbais.n99 0.007
R25715 Nbais.n243 Nbais.n240 0.007
R25716 Nbais.n115 Nbais.n114 0.006
R25717 Nbais.n231 Nbais.n230 0.006
R25718 Nbais.n244 Nbais.n236 0.006
R25719 Nbais.n247 Nbais.n246 0.006
R25720 Nbais.n116 Nbais.n108 0.006
R25721 Nbais.n6 Nbais.n4 0.005
R25722 Nbais.n212 Nbais.n211 0.005
R25723 Nbais.n75 Nbais.n74 0.005
R25724 Nbais.n236 Nbais.n235 0.004
R25725 Nbais.n108 Nbais.n107 0.004
R25726 Nbais.n276 Nbais.n275 0.004
R25727 Nbais.n284 Nbais.n276 0.004
R25728 Nbais.n280 Nbais.n279 0.004
R25729 Nbais.n284 Nbais.n280 0.004
R25730 Nbais.n278 Nbais.n277 0.004
R25731 Nbais.n284 Nbais.n278 0.004
R25732 Nbais.n282 Nbais.n281 0.004
R25733 Nbais.n196 Nbais.n195 0.004
R25734 Nbais.n195 Nbais.n194 0.004
R25735 Nbais.n190 Nbais.n189 0.004
R25736 Nbais.n194 Nbais.n190 0.004
R25737 Nbais.n188 Nbais.n187 0.004
R25738 Nbais.n194 Nbais.n188 0.004
R25739 Nbais.n192 Nbais.n191 0.004
R25740 Nbais.n205 Nbais.n204 0.004
R25741 Nbais.n31 Nbais.n30 0.004
R25742 Nbais.n30 Nbais.n29 0.004
R25743 Nbais.n22 Nbais.n21 0.004
R25744 Nbais.n25 Nbais.n24 0.004
R25745 Nbais.n28 Nbais.n27 0.004
R25746 Nbais.n29 Nbais.n28 0.004
R25747 Nbais.n82 Nbais.n81 0.004
R25748 Nbais.n264 Nbais.n263 0.004
R25749 Nbais.n132 Nbais.n131 0.004
R25750 Nbais.n283 Nbais.n282 0.002
R25751 Nbais.n284 Nbais.n283 0.002
R25752 Nbais.n193 Nbais.n192 0.002
R25753 Nbais.n194 Nbais.n193 0.002
R25754 Nbais.n26 Nbais.n25 0.002
R25755 Nbais.n23 Nbais.n22 0.002
R25756 Nbais.n29 Nbais.n23 0.002
R25757 Nbais.n29 Nbais.n26 0.002
R25758 Nbais.n290 Nbais.n289 0.002
R25759 Nbais.n148 Nbais.n147 0.002
R25760 Nbais.n289 Nbais.n148 0.002
R25761 Nbais.n292 Nbais.n290 0.002
R25762 DN.n1 DN.t1 719.902
R25763 DN.n0 DN.t2 411.605
R25764 DN.n0 DN.t0 236.476
R25765 DN.n1 DN.n0 2.789
R25766 DN DN.n1 0.893
R25767 DNB DNB.t2 719.166
R25768 DNB.n1 DNB.t0 232.401
R25769 DNB.n7 DNB.n6 188.161
R25770 DNB.n18 DNB.t1 23.416
R25771 DNB.n1 DNB.n0 15.764
R25772 DNB.n3 DNB.n2 9.3
R25773 DNB.n9 DNB.n8 9.3
R25774 DNB.n5 DNB.n4 9.3
R25775 DNB DNB.n26 3.97
R25776 DNB.n26 DNB.n17 2.462
R25777 DNB.n26 DNB.n25 2.037
R25778 DNB.n3 DNB.n1 1.248
R25779 DNB.n23 DNB.n21 1.137
R25780 DNB.n19 DNB.n18 1.065
R25781 DNB.n11 DNB.n10 1.037
R25782 DNB.n15 DNB.n13 0.853
R25783 DNB.n8 DNB.n7 0.705
R25784 DNB.n25 DNB.n24 0.7
R25785 DNB.n17 DNB.n16 0.7
R25786 DNB.n10 DNB.n9 0.127
R25787 DNB.n13 DNB.n12 0.041
R25788 DNB.n9 DNB.n5 0.04
R25789 DNB.n21 DNB.n20 0.019
R25790 DNB.n15 DNB.n14 0.013
R25791 DNB.n13 DNB.n11 0.009
R25792 DNB.n5 DNB.n3 0.005
R25793 DNB.n21 DNB.n19 0.005
R25794 DNB.n16 DNB.n15 0.004
R25795 DNB.n24 DNB.n23 0.004
R25796 DNB.n23 DNB.n22 0.001
R25797 net1.n255 net1.t2 124.695
R25798 net1.n235 net1.t3 124.695
R25799 net1.n143 net1.n142 92.5
R25800 net1.n194 net1.n193 92.5
R25801 net1.n15 net1.n14 92.5
R25802 net1.n78 net1.n77 92.5
R25803 net1.n254 net1.n253 92.5
R25804 net1.n234 net1.n233 92.5
R25805 net1.n142 net1.t1 70.344
R25806 net1.n14 net1.t0 70.344
R25807 net1.n133 net1.n132 31.034
R25808 net1.n211 net1.n210 31.034
R25809 net1.n28 net1.n27 31.034
R25810 net1.n95 net1.n94 31.034
R25811 net1.n264 net1.n263 31.034
R25812 net1.n244 net1.n243 31.034
R25813 net1.n255 net1.n254 15.431
R25814 net1.n235 net1.n234 15.431
R25815 net1.n154 net1.n153 9.3
R25816 net1.n134 net1.n133 9.3
R25817 net1.n212 net1.n211 9.3
R25818 net1.n220 net1.n219 9.3
R25819 net1.n38 net1.n37 9.3
R25820 net1.n104 net1.n103 9.3
R25821 net1.n96 net1.n95 9.3
R25822 net1.n29 net1.n28 9.3
R25823 net1.n270 net1.n269 9.3
R25824 net1.n259 net1.n258 9.3
R25825 net1.n257 net1.n256 9.3
R25826 net1.n266 net1.n265 9.3
R25827 net1.n265 net1.n264 9.3
R25828 net1.n268 net1.n267 9.3
R25829 net1.n272 net1.n271 9.3
R25830 net1.n250 net1.n249 9.3
R25831 net1.n239 net1.n238 9.3
R25832 net1.n237 net1.n236 9.3
R25833 net1.n246 net1.n245 9.3
R25834 net1.n245 net1.n244 9.3
R25835 net1.n248 net1.n247 9.3
R25836 net1.n252 net1.n251 9.3
R25837 net1.n144 net1.n143 8.282
R25838 net1.n195 net1.n194 8.282
R25839 net1.n16 net1.n15 8.282
R25840 net1.n79 net1.n78 8.282
R25841 net1.n273 net1.n252 6.035
R25842 net1.n273 net1.n272 6.02
R25843 net1.n134 net1.n130 5.647
R25844 net1.n212 net1.n208 5.647
R25845 net1.n29 net1.n25 5.647
R25846 net1.n96 net1.n92 5.647
R25847 net1.n265 net1.n261 5.647
R25848 net1.n245 net1.n241 5.647
R25849 net1.n192 net1.n191 4.65
R25850 net1.n76 net1.n75 4.65
R25851 net1.n226 net1.n224 4.5
R25852 net1.n214 net1.n213 4.5
R25853 net1.n203 net1.n202 4.5
R25854 net1.n196 net1.n195 4.5
R25855 net1.n148 net1.n136 4.5
R25856 net1.n145 net1.n144 4.5
R25857 net1.n190 net1.n189 4.5
R25858 net1.n159 net1.n158 4.5
R25859 net1.n80 net1.n79 4.5
R25860 net1.n87 net1.n86 4.5
R25861 net1.n21 net1.n16 4.5
R25862 net1.n98 net1.n97 4.5
R25863 net1.n74 net1.n73 4.5
R25864 net1.n32 net1.n31 4.5
R25865 net1.n110 net1.n108 4.5
R25866 net1.n43 net1.n42 4.5
R25867 net1.n132 net1.n131 4.137
R25868 net1.n210 net1.n209 4.137
R25869 net1.n27 net1.n26 4.137
R25870 net1.n94 net1.n93 4.137
R25871 net1.n263 net1.n262 4.137
R25872 net1.n243 net1.n242 4.137
R25873 net1.n158 net1.n156 3.764
R25874 net1.n213 net1.n206 3.764
R25875 net1.n42 net1.n40 3.764
R25876 net1.n97 net1.n90 3.764
R25877 net1.n136 net1.n135 3.388
R25878 net1.n224 net1.n223 3.388
R25879 net1.n31 net1.n30 3.388
R25880 net1.n108 net1.n107 3.388
R25881 net1.n136 net1.n134 3.011
R25882 net1.n144 net1.n141 3.011
R25883 net1.n224 net1.n222 3.011
R25884 net1.n31 net1.n29 3.011
R25885 net1.n16 net1.n13 3.011
R25886 net1.n108 net1.n106 3.011
R25887 net1.n158 net1.n157 2.635
R25888 net1.n202 net1.n201 2.635
R25889 net1.n213 net1.n212 2.635
R25890 net1.n42 net1.n41 2.635
R25891 net1.n86 net1.n85 2.635
R25892 net1.n97 net1.n96 2.635
R25893 net1.n232 net1.n115 1.63
R25894 net1.n257 net1.n255 1.57
R25895 net1.n237 net1.n235 1.57
R25896 net1.n227 net1.n226 1.5
R25897 net1.n160 net1.n159 1.5
R25898 net1.n111 net1.n110 1.5
R25899 net1.n44 net1.n43 1.5
R25900 net1.n232 net1.n231 1.473
R25901 net1 net1.n273 1.46
R25902 net1.n230 net1.n229 0.853
R25903 net1.n114 net1.n113 0.853
R25904 net1.n130 net1.n129 0.752
R25905 net1.n208 net1.n207 0.752
R25906 net1.n25 net1.n24 0.752
R25907 net1.n92 net1.n91 0.752
R25908 net1.n261 net1.n260 0.752
R25909 net1.n241 net1.n240 0.752
R25910 net1.n46 net1.n45 0.704
R25911 net1.n162 net1.n161 0.702
R25912 net1 net1.n232 0.341
R25913 net1.n268 net1.n266 0.144
R25914 net1.n248 net1.n246 0.144
R25915 net1.n266 net1.n259 0.04
R25916 net1.n246 net1.n239 0.04
R25917 net1.n138 net1.n137 0.035
R25918 net1.n198 net1.n197 0.035
R25919 net1.n117 net1.n116 0.035
R25920 net1.n179 net1.n178 0.035
R25921 net1.n18 net1.n17 0.035
R25922 net1.n82 net1.n81 0.035
R25923 net1.n1 net1.n0 0.035
R25924 net1.n63 net1.n62 0.035
R25925 net1.n272 net1.n270 0.035
R25926 net1.n252 net1.n250 0.035
R25927 net1.n127 net1.n126 0.034
R25928 net1.n188 net1.n187 0.034
R25929 net1.n11 net1.n10 0.034
R25930 net1.n72 net1.n71 0.034
R25931 net1.n217 net1.n216 0.032
R25932 net1.n186 net1.n185 0.032
R25933 net1.n101 net1.n100 0.032
R25934 net1.n70 net1.n69 0.032
R25935 net1.n163 net1.n162 0.031
R25936 net1.n174 net1.n173 0.031
R25937 net1.n47 net1.n46 0.031
R25938 net1.n58 net1.n57 0.031
R25939 net1.n151 net1.n150 0.03
R25940 net1.n220 net1.n218 0.03
R25941 net1.n125 net1.n124 0.03
R25942 net1.n184 net1.n183 0.03
R25943 net1.n35 net1.n34 0.03
R25944 net1.n104 net1.n102 0.03
R25945 net1.n9 net1.n8 0.03
R25946 net1.n68 net1.n67 0.03
R25947 net1.n154 net1.n152 0.028
R25948 net1.n140 net1.n139 0.028
R25949 net1.n200 net1.n199 0.028
R25950 net1.n122 net1.n121 0.028
R25951 net1.n119 net1.n118 0.028
R25952 net1.n181 net1.n180 0.028
R25953 net1.n227 net1.n188 0.028
R25954 net1.n38 net1.n36 0.028
R25955 net1.n20 net1.n19 0.028
R25956 net1.n84 net1.n83 0.028
R25957 net1.n6 net1.n5 0.028
R25958 net1.n3 net1.n2 0.028
R25959 net1.n65 net1.n64 0.028
R25960 net1.n111 net1.n72 0.028
R25961 net1.n161 net1.n160 0.028
R25962 net1.n45 net1.n44 0.027
R25963 net1.n167 net1.n166 0.027
R25964 net1.n170 net1.n169 0.027
R25965 net1.n51 net1.n50 0.027
R25966 net1.n54 net1.n53 0.027
R25967 net1.n160 net1.n127 0.026
R25968 net1.n44 net1.n11 0.026
R25969 net1.n196 net1.n192 0.022
R25970 net1.n177 net1.n176 0.022
R25971 net1.n229 net1.n227 0.022
R25972 net1.n80 net1.n76 0.022
R25973 net1.n61 net1.n60 0.022
R25974 net1.n113 net1.n111 0.022
R25975 net1.n192 net1.n190 0.02
R25976 net1.n176 net1.n175 0.02
R25977 net1.n76 net1.n74 0.02
R25978 net1.n60 net1.n59 0.02
R25979 net1.n230 net1.n174 0.019
R25980 net1.n231 net1.n230 0.019
R25981 net1.n114 net1.n58 0.019
R25982 net1.n115 net1.n114 0.019
R25983 net1.n159 net1.n128 0.018
R25984 net1.n155 net1.n154 0.018
R25985 net1.n152 net1.n151 0.018
R25986 net1.n214 net1.n205 0.018
R25987 net1.n126 net1.n125 0.018
R25988 net1.n43 net1.n12 0.018
R25989 net1.n39 net1.n38 0.018
R25990 net1.n36 net1.n35 0.018
R25991 net1.n98 net1.n89 0.018
R25992 net1.n10 net1.n9 0.018
R25993 net1.n148 net1.n147 0.017
R25994 net1.n218 net1.n217 0.017
R25995 net1.n221 net1.n220 0.017
R25996 net1.n226 net1.n225 0.017
R25997 net1.n124 net1.n123 0.017
R25998 net1.n185 net1.n184 0.017
R25999 net1.n187 net1.n186 0.017
R26000 net1.n32 net1.n23 0.017
R26001 net1.n102 net1.n101 0.017
R26002 net1.n105 net1.n104 0.017
R26003 net1.n110 net1.n109 0.017
R26004 net1.n8 net1.n7 0.017
R26005 net1.n69 net1.n68 0.017
R26006 net1.n71 net1.n70 0.017
R26007 net1.n149 net1.n148 0.015
R26008 net1.n146 net1.n145 0.015
R26009 net1.n226 net1.n221 0.015
R26010 net1.n121 net1.n120 0.015
R26011 net1.n33 net1.n32 0.015
R26012 net1.n22 net1.n21 0.015
R26013 net1.n110 net1.n105 0.015
R26014 net1.n5 net1.n4 0.015
R26015 net1.n159 net1.n155 0.013
R26016 net1.n204 net1.n203 0.013
R26017 net1.n215 net1.n214 0.013
R26018 net1.n183 net1.n182 0.013
R26019 net1.n43 net1.n39 0.013
R26020 net1.n88 net1.n87 0.013
R26021 net1.n99 net1.n98 0.013
R26022 net1.n67 net1.n66 0.013
R26023 net1.n168 net1.n167 0.012
R26024 net1.n169 net1.n168 0.012
R26025 net1.n52 net1.n51 0.012
R26026 net1.n53 net1.n52 0.012
R26027 net1.n229 net1.n228 0.012
R26028 net1.n113 net1.n112 0.012
R26029 net1.n147 net1.n146 0.011
R26030 net1.n205 net1.n204 0.011
R26031 net1.n165 net1.n164 0.011
R26032 net1.n172 net1.n171 0.011
R26033 net1.n23 net1.n22 0.011
R26034 net1.n89 net1.n88 0.011
R26035 net1.n49 net1.n48 0.011
R26036 net1.n56 net1.n55 0.011
R26037 net1.n270 net1.n268 0.01
R26038 net1.n250 net1.n248 0.01
R26039 net1.n197 net1.n196 0.009
R26040 net1.n178 net1.n177 0.009
R26041 net1.n81 net1.n80 0.009
R26042 net1.n62 net1.n61 0.009
R26043 net1.n139 net1.n138 0.007
R26044 net1.n199 net1.n198 0.007
R26045 net1.n118 net1.n117 0.007
R26046 net1.n180 net1.n179 0.007
R26047 net1.n19 net1.n18 0.007
R26048 net1.n83 net1.n82 0.007
R26049 net1.n2 net1.n1 0.007
R26050 net1.n64 net1.n63 0.007
R26051 net1.n164 net1.n163 0.006
R26052 net1.n166 net1.n165 0.006
R26053 net1.n171 net1.n170 0.006
R26054 net1.n173 net1.n172 0.006
R26055 net1.n48 net1.n47 0.006
R26056 net1.n50 net1.n49 0.006
R26057 net1.n55 net1.n54 0.006
R26058 net1.n57 net1.n56 0.006
R26059 net1.n259 net1.n257 0.005
R26060 net1.n239 net1.n237 0.005
R26061 net1.n150 net1.n149 0.003
R26062 net1.n203 net1.n200 0.003
R26063 net1.n216 net1.n215 0.003
R26064 net1.n182 net1.n181 0.003
R26065 net1.n34 net1.n33 0.003
R26066 net1.n87 net1.n84 0.003
R26067 net1.n100 net1.n99 0.003
R26068 net1.n66 net1.n65 0.003
R26069 net1.n145 net1.n140 0.001
R26070 net1.n123 net1.n122 0.001
R26071 net1.n120 net1.n119 0.001
R26072 net1.n21 net1.n20 0.001
R26073 net1.n7 net1.n6 0.001
R26074 net1.n4 net1.n3 0.001
R26075 a_48058_n6837.n12 a_48058_n6837.t3 46.604
R26076 a_48058_n6837.n12 a_48058_n6837.t2 46.357
R26077 a_48058_n6837.n9 a_48058_n6837.t0 28.565
R26078 a_48058_n6837.t1 a_48058_n6837.n21 17.4
R26079 a_48058_n6837.n10 a_48058_n6837.n9 9.02
R26080 a_48058_n6837.n1 a_48058_n6837.n0 8.658
R26081 a_48058_n6837.n21 a_48058_n6837.n20 8.5
R26082 a_48058_n6837.n21 a_48058_n6837.n15 8.5
R26083 a_48058_n6837.n14 a_48058_n6837.n13 8.111
R26084 a_48058_n6837.n7 a_48058_n6837.n6 4.542
R26085 a_48058_n6837.n7 a_48058_n6837.n5 4.5
R26086 a_48058_n6837.n6 a_48058_n6837.n8 4.141
R26087 a_48058_n6837.n14 a_48058_n6837.n3 4.141
R26088 a_48058_n6837.n13 a_48058_n6837.n12 3.984
R26089 a_48058_n6837.n19 a_48058_n6837.n18 3.764
R26090 a_48058_n6837.n17 a_48058_n6837.n16 3.764
R26091 a_48058_n6837.n5 a_48058_n6837.n4 3.388
R26092 a_48058_n6837.n2 a_48058_n6837.n1 3.388
R26093 a_48058_n6837.n20 a_48058_n6837.n19 2.635
R26094 a_48058_n6837.n6 a_48058_n6837.n10 2.258
R26095 a_48058_n6837.n15 a_48058_n6837.n14 2.258
R26096 a_48058_n6837.n18 a_48058_n6837.n17 1.129
R26097 a_48058_n6837.n3 a_48058_n6837.n2 1.129
R26098 a_48058_n6837.n13 a_48058_n6837.n11 1.124
R26099 a_48058_n6837.n11 a_48058_n6837.n7 0.73
R26100 net5_ota.n64 net5_ota.t2 27.367
R26101 net5_ota.n18 net5_ota.t1 13.384
R26102 net5_ota.n127 net5_ota.n126 9.3
R26103 net5_ota.n229 net5_ota.n228 9.3
R26104 net5_ota.n193 net5_ota.n192 9.154
R26105 net5_ota.n19 net5_ota.n18 8.855
R26106 net5_ota.n192 net5_ota.t0 7.141
R26107 net5_ota.n36 net5_ota.n35 7.03
R26108 net5_ota.n287 net5_ota.n286 7.029
R26109 net5_ota.n71 net5_ota.n70 7.029
R26110 net5_ota.n59 net5_ota.n58 6.681
R26111 net5_ota.n20 net5_ota.n19 4.65
R26112 net5_ota.n194 net5_ota.n193 4.65
R26113 net5_ota.n30 net5_ota.n29 4.5
R26114 net5_ota.n53 net5_ota.n52 4.5
R26115 net5_ota.n17 net5_ota.n16 4.5
R26116 net5_ota.n22 net5_ota.n21 4.5
R26117 net5_ota.n93 net5_ota.n88 4.5
R26118 net5_ota.n232 net5_ota.n224 4.5
R26119 net5_ota.n256 net5_ota.n250 4.5
R26120 net5_ota.n211 net5_ota.n210 4.5
R26121 net5_ota.n181 net5_ota.n178 4.5
R26122 net5_ota.n196 net5_ota.n190 4.5
R26123 net5_ota.n170 net5_ota.n167 4.5
R26124 net5_ota.n186 net5_ota.n185 4.5
R26125 net5_ota.n160 net5_ota.n155 4.5
R26126 net5_ota.n138 net5_ota.n137 4.5
R26127 net5_ota.n112 net5_ota.n108 4.5
R26128 net5_ota.n275 net5_ota.n274 4.5
R26129 net5_ota.n64 net5_ota.n63 4.225
R26130 net5_ota.n250 net5_ota.n247 4.141
R26131 net5_ota.n108 net5_ota.n107 4.141
R26132 net5_ota.n224 net5_ota.n221 3.764
R26133 net5_ota.n155 net5_ota.n153 3.764
R26134 net5_ota.n274 net5_ota.n271 3.388
R26135 net5_ota.n210 net5_ota.n209 3.388
R26136 net5_ota.n137 net5_ota.n136 3.388
R26137 net5_ota.n88 net5_ota.n87 3.388
R26138 net5_ota.n52 net5_ota.n50 3.011
R26139 net5_ota.n274 net5_ota.n273 3.011
R26140 net5_ota.n210 net5_ota.n207 3.011
R26141 net5_ota.n178 net5_ota.n176 3.011
R26142 net5_ota.n126 net5_ota.n125 3.011
R26143 net5_ota.n137 net5_ota.n135 3.011
R26144 net5_ota.n88 net5_ota.n86 3.011
R26145 net5_ota.n29 net5_ota.n28 2.635
R26146 net5_ota.n224 net5_ota.n223 2.635
R26147 net5_ota.n228 net5_ota.n227 2.635
R26148 net5_ota.n167 net5_ota.n166 2.635
R26149 net5_ota.n155 net5_ota.n154 2.635
R26150 net5_ota.n250 net5_ota.n249 2.258
R26151 net5_ota.n108 net5_ota.n106 2.258
R26152 net5_ota net5_ota.n64 2.164
R26153 net5_ota net5_ota.n301 2.112
R26154 net5_ota.n29 net5_ota.n27 1.505
R26155 net5_ota.n167 net5_ota.n165 1.505
R26156 net5_ota.n74 net5_ota.n72 1.5
R26157 net5_ota.n94 net5_ota.n93 1.5
R26158 net5_ota.n257 net5_ota.n256 1.5
R26159 net5_ota.n293 net5_ota.n292 1.5
R26160 net5_ota.n233 net5_ota.n232 1.5
R26161 net5_ota.n212 net5_ota.n211 1.5
R26162 net5_ota.n182 net5_ota.n181 1.5
R26163 net5_ota.n197 net5_ota.n196 1.5
R26164 net5_ota.n171 net5_ota.n170 1.5
R26165 net5_ota.n187 net5_ota.n186 1.5
R26166 net5_ota.n161 net5_ota.n160 1.5
R26167 net5_ota.n139 net5_ota.n138 1.5
R26168 net5_ota.n113 net5_ota.n112 1.5
R26169 net5_ota.n276 net5_ota.n275 1.5
R26170 net5_ota.n37 net5_ota.n36 1.399
R26171 net5_ota.n62 net5_ota.n59 1.395
R26172 net5_ota.n63 net5_ota.n62 1.137
R26173 net5_ota.n46 net5_ota.n45 1.137
R26174 net5_ota.n76 net5_ota.n75 1.137
R26175 net5_ota.n96 net5_ota.n95 1.137
R26176 net5_ota.n115 net5_ota.n114 1.137
R26177 net5_ota.n123 net5_ota.n122 1.137
R26178 net5_ota.n141 net5_ota.n140 1.137
R26179 net5_ota.n148 net5_ota.n147 1.137
R26180 net5_ota.n241 net5_ota.n240 1.137
R26181 net5_ota.n299 net5_ota.n298 1.137
R26182 net5_ota.n262 net5_ota.n261 1.137
R26183 net5_ota.n216 net5_ota.n215 1.137
R26184 net5_ota.n237 net5_ota.n236 1.137
R26185 net5_ota.n199 net5_ota.n198 1.137
R26186 net5_ota.n175 net5_ota.n174 1.137
R26187 net5_ota.n283 net5_ota.n282 1.137
R26188 net5_ota.n52 net5_ota.n51 1.129
R26189 net5_ota.n178 net5_ota.n177 1.129
R26190 net5_ota.n38 net5_ota.n37 0.862
R26191 net5_ota.n286 net5_ota.n285 0.155
R26192 net5_ota.n70 net5_ota.n69 0.155
R26193 net5_ota.n273 net5_ota.n272 0.144
R26194 net5_ota.n86 net5_ota.n85 0.144
R26195 net5_ota.n249 net5_ota.n248 0.133
R26196 net5_ota.n106 net5_ota.n105 0.132
R26197 net5_ota.n229 net5_ota.n226 0.051
R26198 net5_ota.n170 net5_ota.n164 0.046
R26199 net5_ota.n214 net5_ota.n213 0.045
R26200 net5_ota.n198 net5_ota.n197 0.045
R26201 net5_ota.n299 net5_ota.n283 0.045
R26202 net5_ota.n199 net5_ota.n175 0.045
R26203 net5_ota.n96 net5_ota.n76 0.045
R26204 net5_ota.n181 net5_ota.n180 0.044
R26205 net5_ota.n113 net5_ota.n101 0.043
R26206 net5_ota.n253 net5_ota.n252 0.042
R26207 net5_ota.n158 net5_ota.n157 0.042
R26208 net5_ota.n94 net5_ota.n81 0.041
R26209 net5_ota.n90 net5_ota.n89 0.04
R26210 net5_ota.n298 net5_ota.n297 0.039
R26211 net5_ota.n75 net5_ota.n65 0.037
R26212 net5_ota.n58 net5_ota.n57 0.036
R26213 net5_ota.n35 net5_ota.n34 0.036
R26214 net5_ota.n15 net5_ota.n14 0.035
R26215 net5_ota.n24 net5_ota.n23 0.035
R26216 net5_ota.n2 net5_ota.n1 0.035
R26217 net5_ota.n7 net5_ota.n6 0.035
R26218 net5_ota.n290 net5_ota.n289 0.035
R26219 net5_ota.n296 net5_ota.n295 0.034
R26220 net5_ota.n189 net5_ota.n188 0.034
R26221 net5_ota.n80 net5_ota.n79 0.034
R26222 net5_ota.n67 net5_ota.n66 0.033
R26223 net5_ota.n293 net5_ota.n284 0.032
R26224 net5_ota.n172 net5_ota.n171 0.032
R26225 net5_ota.n162 net5_ota.n161 0.032
R26226 net5_ota.n269 net5_ota.n268 0.031
R26227 net5_ota.n132 net5_ota.n131 0.031
R26228 net5_ota.n12 net5_ota.n11 0.03
R26229 net5_ota.n279 net5_ota.n278 0.03
R26230 net5_ota.n212 net5_ota.n202 0.03
R26231 net5_ota.n183 net5_ota.n182 0.03
R26232 net5_ota.n83 net5_ota.n82 0.029
R26233 net5_ota.n92 net5_ota.n91 0.029
R26234 net5_ota.n26 net5_ota.n25 0.028
R26235 net5_ota.n9 net5_ota.n8 0.028
R26236 net5_ota.n100 net5_ota.n99 0.028
R26237 net5_ota.n263 net5_ota.n262 0.028
R26238 net5_ota.n216 net5_ota.n201 0.028
R26239 net5_ota.n149 net5_ota.n148 0.028
R26240 net5_ota.n115 net5_ota.n98 0.028
R26241 net5_ota.n267 net5_ota.n266 0.026
R26242 net5_ota.n246 net5_ota.n245 0.026
R26243 net5_ota.n254 net5_ota.n253 0.026
R26244 net5_ota.n111 net5_ota.n110 0.026
R26245 net5_ota.n281 net5_ota.n280 0.026
R26246 net5_ota.n256 net5_ota.n246 0.024
R26247 net5_ota.n103 net5_ota.n102 0.024
R26248 net5_ota.n112 net5_ota.n111 0.024
R26249 net5_ota.n261 net5_ota.n260 0.024
R26250 net5_ota.n239 net5_ota.n238 0.024
R26251 net5_ota.n236 net5_ota.n235 0.024
R26252 net5_ota.n147 net5_ota.n146 0.024
R26253 net5_ota.n122 net5_ota.n121 0.024
R26254 net5_ota.n78 net5_ota.n77 0.024
R26255 net5_ota.n241 net5_ota.n237 0.024
R26256 net5_ota.n141 net5_ota.n123 0.024
R26257 net5_ota.n223 net5_ota.n222 0.024
R26258 net5_ota.n135 net5_ota.n134 0.024
R26259 net5_ota.n22 net5_ota.n20 0.022
R26260 net5_ota.n5 net5_ota.n4 0.022
R26261 net5_ota.n46 net5_ota.n42 0.022
R26262 net5_ota.n40 net5_ota.n39 0.022
R26263 net5_ota.n232 net5_ota.n220 0.022
R26264 net5_ota.n230 net5_ota.n229 0.022
R26265 net5_ota.n139 net5_ota.n124 0.022
R26266 net5_ota.n20 net5_ota.n17 0.02
R26267 net5_ota.n4 net5_ota.n3 0.02
R26268 net5_ota.n275 net5_ota.n267 0.02
R26269 net5_ota.n211 net5_ota.n206 0.02
R26270 net5_ota.n195 net5_ota.n194 0.02
R26271 net5_ota.n194 net5_ota.n191 0.02
R26272 net5_ota.n128 net5_ota.n127 0.02
R26273 net5_ota.n138 net5_ota.n133 0.02
R26274 net5_ota.n93 net5_ota.n92 0.02
R26275 net5_ota.n33 net5_ota.n32 0.018
R26276 net5_ota.n74 net5_ota.n73 0.017
R26277 net5_ota.n56 net5_ota.n55 0.017
R26278 net5_ota.n62 net5_ota.n61 0.017
R26279 net5_ota.n280 net5_ota.n279 0.017
R26280 net5_ota.n54 net5_ota.n53 0.015
R26281 net5_ota.n44 net5_ota.n43 0.015
R26282 net5_ota.n170 net5_ota.n169 0.015
R26283 net5_ota.n138 net5_ota.n129 0.015
R26284 net5_ota.n235 net5_ota.n234 0.015
R26285 net5_ota.n146 net5_ota.n145 0.015
R26286 net5_ota.n301 net5_ota.n300 0.014
R26287 net5_ota.n264 net5_ota.n263 0.014
R26288 net5_ota.n201 net5_ota.n200 0.014
R26289 net5_ota.n150 net5_ota.n149 0.014
R26290 net5_ota.n98 net5_ota.n97 0.014
R26291 net5_ota.n37 net5_ota.n12 0.013
R26292 net5_ota.n31 net5_ota.n30 0.013
R26293 net5_ota.n11 net5_ota.n10 0.013
R26294 net5_ota.n252 net5_ota.n251 0.013
R26295 net5_ota.n232 net5_ota.n231 0.013
R26296 net5_ota.n204 net5_ota.n203 0.013
R26297 net5_ota.n206 net5_ota.n205 0.013
R26298 net5_ota.n169 net5_ota.n168 0.013
R26299 net5_ota.n159 net5_ota.n158 0.013
R26300 net5_ota.n140 net5_ota.n139 0.013
R26301 net5_ota.n121 net5_ota.n120 0.013
R26302 net5_ota.n209 net5_ota.n208 0.012
R26303 net5_ota.n153 net5_ota.n152 0.012
R26304 net5_ota.n55 net5_ota.n54 0.011
R26305 net5_ota.n17 net5_ota.n15 0.011
R26306 net5_ota.n32 net5_ota.n31 0.011
R26307 net5_ota.n3 net5_ota.n2 0.011
R26308 net5_ota.n292 net5_ota.n291 0.011
R26309 net5_ota.n291 net5_ota.n290 0.011
R26310 net5_ota.n289 net5_ota.n288 0.011
R26311 net5_ota.n270 net5_ota.n269 0.011
R26312 net5_ota.n131 net5_ota.n130 0.011
R26313 net5_ota.n84 net5_ota.n83 0.011
R26314 net5_ota.n68 net5_ota.n67 0.011
R26315 net5_ota.n72 net5_ota.n68 0.011
R26316 net5_ota.n259 net5_ota.n258 0.011
R26317 net5_ota.n240 net5_ota.n239 0.011
R26318 net5_ota.n236 net5_ota.n233 0.011
R26319 net5_ota.n171 net5_ota.n162 0.011
R26320 net5_ota.n23 net5_ota.n22 0.009
R26321 net5_ota.n6 net5_ota.n5 0.009
R26322 net5_ota.n48 net5_ota.n47 0.009
R26323 net5_ota.n42 net5_ota.n41 0.009
R26324 net5_ota.n41 net5_ota.n40 0.009
R26325 net5_ota.n298 net5_ota.n293 0.009
R26326 net5_ota.n297 net5_ota.n296 0.009
R26327 net5_ota.n282 net5_ota.n281 0.009
R26328 net5_ota.n122 net5_ota.n118 0.009
R26329 net5_ota.n95 net5_ota.n78 0.009
R26330 net5_ota.n75 net5_ota.n74 0.009
R26331 net5_ota.n262 net5_ota.n243 0.008
R26332 net5_ota.n242 net5_ota.n241 0.008
R26333 net5_ota.n237 net5_ota.n218 0.008
R26334 net5_ota.n217 net5_ota.n216 0.008
R26335 net5_ota.n148 net5_ota.n143 0.008
R26336 net5_ota.n142 net5_ota.n141 0.008
R26337 net5_ota.n123 net5_ota.n117 0.008
R26338 net5_ota.n116 net5_ota.n115 0.008
R26339 net5_ota.n14 net5_ota.n13 0.007
R26340 net5_ota.n25 net5_ota.n24 0.007
R26341 net5_ota.n1 net5_ota.n0 0.007
R26342 net5_ota.n8 net5_ota.n7 0.007
R26343 net5_ota.n184 net5_ota.n183 0.007
R26344 net5_ota.n173 net5_ota.n172 0.007
R26345 net5_ota.n275 net5_ota.n270 0.006
R26346 net5_ota.n256 net5_ota.n255 0.006
R26347 net5_ota.n255 net5_ota.n254 0.006
R26348 net5_ota.n220 net5_ota.n219 0.006
R26349 net5_ota.n133 net5_ota.n132 0.006
R26350 net5_ota.n104 net5_ota.n103 0.006
R26351 net5_ota.n112 net5_ota.n104 0.006
R26352 net5_ota.n110 net5_ota.n109 0.006
R26353 net5_ota.n93 net5_ota.n84 0.006
R26354 net5_ota.n63 net5_ota.n48 0.005
R26355 net5_ota.n47 net5_ota.n46 0.005
R26356 net5_ota.n39 net5_ota.n38 0.005
R26357 net5_ota.n282 net5_ota.n276 0.005
R26358 net5_ota.n261 net5_ota.n257 0.005
R26359 net5_ota.n188 net5_ota.n187 0.005
R26360 net5_ota.n114 net5_ota.n113 0.005
R26361 net5_ota.n101 net5_ota.n100 0.005
R26362 net5_ota.n95 net5_ota.n94 0.005
R26363 net5_ota.n243 net5_ota.n242 0.005
R26364 net5_ota.n218 net5_ota.n217 0.005
R26365 net5_ota.n143 net5_ota.n142 0.005
R26366 net5_ota.n117 net5_ota.n116 0.005
R26367 net5_ota.n292 net5_ota.n287 0.005
R26368 net5_ota.n72 net5_ota.n71 0.005
R26369 net5_ota.n59 net5_ota.n56 0.005
R26370 net5_ota.n36 net5_ota.n33 0.004
R26371 net5_ota.n266 net5_ota.n265 0.004
R26372 net5_ota.n245 net5_ota.n244 0.004
R26373 net5_ota.n226 net5_ota.n225 0.004
R26374 net5_ota.n211 net5_ota.n204 0.004
R26375 net5_ota.n196 net5_ota.n195 0.004
R26376 net5_ota.n30 net5_ota.n26 0.003
R26377 net5_ota.n10 net5_ota.n9 0.003
R26378 net5_ota.n295 net5_ota.n294 0.003
R26379 net5_ota.n278 net5_ota.n277 0.003
R26380 net5_ota.n260 net5_ota.n259 0.003
R26381 net5_ota.n215 net5_ota.n214 0.003
R26382 net5_ota.n213 net5_ota.n212 0.003
R26383 net5_ota.n197 net5_ota.n189 0.003
R26384 net5_ota.n300 net5_ota.n299 0.003
R26385 net5_ota.n283 net5_ota.n264 0.003
R26386 net5_ota.n200 net5_ota.n199 0.003
R26387 net5_ota.n175 net5_ota.n150 0.003
R26388 net5_ota.n97 net5_ota.n96 0.003
R26389 net5_ota.n231 net5_ota.n230 0.002
R26390 net5_ota.n180 net5_ota.n179 0.002
R26391 net5_ota.n164 net5_ota.n163 0.002
R26392 net5_ota.n160 net5_ota.n159 0.002
R26393 net5_ota.n157 net5_ota.n156 0.002
R26394 net5_ota.n129 net5_ota.n128 0.002
R26395 net5_ota.n91 net5_ota.n90 0.002
R26396 net5_ota.n53 net5_ota.n49 0.001
R26397 net5_ota.n61 net5_ota.n60 0.001
R26398 net5_ota.n45 net5_ota.n44 0.001
R26399 net5_ota.n198 net5_ota.n184 0.001
R26400 net5_ota.n174 net5_ota.n173 0.001
R26401 net5_ota.n161 net5_ota.n151 0.001
R26402 net5_ota.n147 net5_ota.n144 0.001
R26403 net5_ota.n120 net5_ota.n119 0.001
R26404 net5_ota.n81 net5_ota.n80 0.001
R26405 net7.n3378 net7.n3377 13.176
R26406 net7.n3016 net7.n3015 13.176
R26407 net7.n2654 net7.n2653 13.176
R26408 net7.n2292 net7.n2291 13.176
R26409 net7.n1930 net7.n1929 13.176
R26410 net7.n1568 net7.n1567 13.176
R26411 net7.n1206 net7.n1205 13.176
R26412 net7.n844 net7.n843 13.176
R26413 net7.n482 net7.n481 13.176
R26414 net7.n121 net7.n120 13.176
R26415 net7.n3817 net7.n3816 13.176
R26416 net7.n4178 net7.n4177 13.176
R26417 net7.n4540 net7.n4539 13.176
R26418 net7.n4902 net7.n4901 13.176
R26419 net7.n5264 net7.n5263 13.176
R26420 net7.n5626 net7.n5625 13.176
R26421 net7.n5988 net7.n5987 13.176
R26422 net7.n6350 net7.n6349 13.176
R26423 net7.n6712 net7.n6711 13.176
R26424 net7.n7074 net7.n7073 13.176
R26425 net7.n3412 net7.n3411 9.3
R26426 net7.n3538 net7.n3537 9.3
R26427 net7.n3541 net7.n3540 9.3
R26428 net7.n3549 net7.n3548 9.3
R26429 net7.n3588 net7.n3587 9.3
R26430 net7.n3599 net7.n3598 9.3
R26431 net7.n3590 net7.n3589 9.3
R26432 net7.n3578 net7.n3577 9.3
R26433 net7.n3580 net7.n3579 9.3
R26434 net7.n3552 net7.n3551 9.3
R26435 net7.n3528 net7.n3527 9.3
R26436 net7.n3383 net7.n3382 9.3
R26437 net7.n3414 net7.n3413 9.3
R26438 net7.n3299 net7.n3298 9.3
R26439 net7.n3287 net7.n3286 9.3
R26440 net7.n3285 net7.n3284 9.3
R26441 net7.n3050 net7.n3049 9.3
R26442 net7.n3176 net7.n3175 9.3
R26443 net7.n3179 net7.n3178 9.3
R26444 net7.n3187 net7.n3186 9.3
R26445 net7.n3226 net7.n3225 9.3
R26446 net7.n3237 net7.n3236 9.3
R26447 net7.n3228 net7.n3227 9.3
R26448 net7.n3216 net7.n3215 9.3
R26449 net7.n3218 net7.n3217 9.3
R26450 net7.n3190 net7.n3189 9.3
R26451 net7.n3166 net7.n3165 9.3
R26452 net7.n3021 net7.n3020 9.3
R26453 net7.n3052 net7.n3051 9.3
R26454 net7.n2937 net7.n2936 9.3
R26455 net7.n2925 net7.n2924 9.3
R26456 net7.n2923 net7.n2922 9.3
R26457 net7.n2688 net7.n2687 9.3
R26458 net7.n2814 net7.n2813 9.3
R26459 net7.n2817 net7.n2816 9.3
R26460 net7.n2825 net7.n2824 9.3
R26461 net7.n2864 net7.n2863 9.3
R26462 net7.n2875 net7.n2874 9.3
R26463 net7.n2866 net7.n2865 9.3
R26464 net7.n2854 net7.n2853 9.3
R26465 net7.n2856 net7.n2855 9.3
R26466 net7.n2828 net7.n2827 9.3
R26467 net7.n2804 net7.n2803 9.3
R26468 net7.n2659 net7.n2658 9.3
R26469 net7.n2690 net7.n2689 9.3
R26470 net7.n2575 net7.n2574 9.3
R26471 net7.n2563 net7.n2562 9.3
R26472 net7.n2561 net7.n2560 9.3
R26473 net7.n2326 net7.n2325 9.3
R26474 net7.n2452 net7.n2451 9.3
R26475 net7.n2455 net7.n2454 9.3
R26476 net7.n2463 net7.n2462 9.3
R26477 net7.n2502 net7.n2501 9.3
R26478 net7.n2513 net7.n2512 9.3
R26479 net7.n2504 net7.n2503 9.3
R26480 net7.n2492 net7.n2491 9.3
R26481 net7.n2494 net7.n2493 9.3
R26482 net7.n2466 net7.n2465 9.3
R26483 net7.n2442 net7.n2441 9.3
R26484 net7.n2297 net7.n2296 9.3
R26485 net7.n2328 net7.n2327 9.3
R26486 net7.n2213 net7.n2212 9.3
R26487 net7.n2201 net7.n2200 9.3
R26488 net7.n2199 net7.n2198 9.3
R26489 net7.n1964 net7.n1963 9.3
R26490 net7.n2090 net7.n2089 9.3
R26491 net7.n2093 net7.n2092 9.3
R26492 net7.n2101 net7.n2100 9.3
R26493 net7.n2140 net7.n2139 9.3
R26494 net7.n2151 net7.n2150 9.3
R26495 net7.n2142 net7.n2141 9.3
R26496 net7.n2130 net7.n2129 9.3
R26497 net7.n2132 net7.n2131 9.3
R26498 net7.n2104 net7.n2103 9.3
R26499 net7.n2080 net7.n2079 9.3
R26500 net7.n1935 net7.n1934 9.3
R26501 net7.n1966 net7.n1965 9.3
R26502 net7.n1851 net7.n1850 9.3
R26503 net7.n1839 net7.n1838 9.3
R26504 net7.n1837 net7.n1836 9.3
R26505 net7.n1602 net7.n1601 9.3
R26506 net7.n1728 net7.n1727 9.3
R26507 net7.n1731 net7.n1730 9.3
R26508 net7.n1739 net7.n1738 9.3
R26509 net7.n1778 net7.n1777 9.3
R26510 net7.n1789 net7.n1788 9.3
R26511 net7.n1780 net7.n1779 9.3
R26512 net7.n1768 net7.n1767 9.3
R26513 net7.n1770 net7.n1769 9.3
R26514 net7.n1742 net7.n1741 9.3
R26515 net7.n1718 net7.n1717 9.3
R26516 net7.n1573 net7.n1572 9.3
R26517 net7.n1604 net7.n1603 9.3
R26518 net7.n1489 net7.n1488 9.3
R26519 net7.n1477 net7.n1476 9.3
R26520 net7.n1475 net7.n1474 9.3
R26521 net7.n1240 net7.n1239 9.3
R26522 net7.n1366 net7.n1365 9.3
R26523 net7.n1369 net7.n1368 9.3
R26524 net7.n1377 net7.n1376 9.3
R26525 net7.n1416 net7.n1415 9.3
R26526 net7.n1427 net7.n1426 9.3
R26527 net7.n1418 net7.n1417 9.3
R26528 net7.n1406 net7.n1405 9.3
R26529 net7.n1408 net7.n1407 9.3
R26530 net7.n1380 net7.n1379 9.3
R26531 net7.n1356 net7.n1355 9.3
R26532 net7.n1211 net7.n1210 9.3
R26533 net7.n1242 net7.n1241 9.3
R26534 net7.n1127 net7.n1126 9.3
R26535 net7.n1115 net7.n1114 9.3
R26536 net7.n1113 net7.n1112 9.3
R26537 net7.n878 net7.n877 9.3
R26538 net7.n1004 net7.n1003 9.3
R26539 net7.n1007 net7.n1006 9.3
R26540 net7.n1015 net7.n1014 9.3
R26541 net7.n1054 net7.n1053 9.3
R26542 net7.n1065 net7.n1064 9.3
R26543 net7.n1056 net7.n1055 9.3
R26544 net7.n1044 net7.n1043 9.3
R26545 net7.n1046 net7.n1045 9.3
R26546 net7.n1018 net7.n1017 9.3
R26547 net7.n994 net7.n993 9.3
R26548 net7.n849 net7.n848 9.3
R26549 net7.n880 net7.n879 9.3
R26550 net7.n765 net7.n764 9.3
R26551 net7.n753 net7.n752 9.3
R26552 net7.n751 net7.n750 9.3
R26553 net7.n516 net7.n515 9.3
R26554 net7.n642 net7.n641 9.3
R26555 net7.n645 net7.n644 9.3
R26556 net7.n653 net7.n652 9.3
R26557 net7.n692 net7.n691 9.3
R26558 net7.n703 net7.n702 9.3
R26559 net7.n694 net7.n693 9.3
R26560 net7.n682 net7.n681 9.3
R26561 net7.n684 net7.n683 9.3
R26562 net7.n656 net7.n655 9.3
R26563 net7.n632 net7.n631 9.3
R26564 net7.n487 net7.n486 9.3
R26565 net7.n518 net7.n517 9.3
R26566 net7.n403 net7.n402 9.3
R26567 net7.n391 net7.n390 9.3
R26568 net7.n389 net7.n388 9.3
R26569 net7.n342 net7.n341 9.3
R26570 net7.n155 net7.n154 9.3
R26571 net7.n281 net7.n280 9.3
R26572 net7.n284 net7.n283 9.3
R26573 net7.n292 net7.n291 9.3
R26574 net7.n331 net7.n330 9.3
R26575 net7.n333 net7.n332 9.3
R26576 net7.n321 net7.n320 9.3
R26577 net7.n323 net7.n322 9.3
R26578 net7.n295 net7.n294 9.3
R26579 net7.n271 net7.n270 9.3
R26580 net7.n126 net7.n125 9.3
R26581 net7.n157 net7.n156 9.3
R26582 net7.n42 net7.n41 9.3
R26583 net7.n30 net7.n29 9.3
R26584 net7.n28 net7.n27 9.3
R26585 net7.n3793 net7.n3792 9.3
R26586 net7.n3674 net7.n3673 9.3
R26587 net7.n3676 net7.n3675 9.3
R26588 net7.n3685 net7.n3684 9.3
R26589 net7.n3667 net7.n3666 9.3
R26590 net7.n3669 net7.n3668 9.3
R26591 net7.n3780 net7.n3779 9.3
R26592 net7.n3822 net7.n3821 9.3
R26593 net7.n3806 net7.n3805 9.3
R26594 net7.n3795 net7.n3794 9.3
R26595 net7.n3782 net7.n3781 9.3
R26596 net7.n3836 net7.n3835 9.3
R26597 net7.n3838 net7.n3837 9.3
R26598 net7.n3966 net7.n3965 9.3
R26599 net7.n3954 net7.n3953 9.3
R26600 net7.n3952 net7.n3951 9.3
R26601 net7.n4154 net7.n4153 9.3
R26602 net7.n4035 net7.n4034 9.3
R26603 net7.n4037 net7.n4036 9.3
R26604 net7.n4046 net7.n4045 9.3
R26605 net7.n4028 net7.n4027 9.3
R26606 net7.n4030 net7.n4029 9.3
R26607 net7.n4141 net7.n4140 9.3
R26608 net7.n4183 net7.n4182 9.3
R26609 net7.n4167 net7.n4166 9.3
R26610 net7.n4156 net7.n4155 9.3
R26611 net7.n4143 net7.n4142 9.3
R26612 net7.n4197 net7.n4196 9.3
R26613 net7.n4199 net7.n4198 9.3
R26614 net7.n4327 net7.n4326 9.3
R26615 net7.n4315 net7.n4314 9.3
R26616 net7.n4313 net7.n4312 9.3
R26617 net7.n4516 net7.n4515 9.3
R26618 net7.n4397 net7.n4396 9.3
R26619 net7.n4399 net7.n4398 9.3
R26620 net7.n4408 net7.n4407 9.3
R26621 net7.n4390 net7.n4389 9.3
R26622 net7.n4392 net7.n4391 9.3
R26623 net7.n4503 net7.n4502 9.3
R26624 net7.n4545 net7.n4544 9.3
R26625 net7.n4529 net7.n4528 9.3
R26626 net7.n4518 net7.n4517 9.3
R26627 net7.n4505 net7.n4504 9.3
R26628 net7.n4559 net7.n4558 9.3
R26629 net7.n4561 net7.n4560 9.3
R26630 net7.n4689 net7.n4688 9.3
R26631 net7.n4677 net7.n4676 9.3
R26632 net7.n4675 net7.n4674 9.3
R26633 net7.n4878 net7.n4877 9.3
R26634 net7.n4759 net7.n4758 9.3
R26635 net7.n4761 net7.n4760 9.3
R26636 net7.n4770 net7.n4769 9.3
R26637 net7.n4752 net7.n4751 9.3
R26638 net7.n4754 net7.n4753 9.3
R26639 net7.n4865 net7.n4864 9.3
R26640 net7.n4907 net7.n4906 9.3
R26641 net7.n4891 net7.n4890 9.3
R26642 net7.n4880 net7.n4879 9.3
R26643 net7.n4867 net7.n4866 9.3
R26644 net7.n4921 net7.n4920 9.3
R26645 net7.n4923 net7.n4922 9.3
R26646 net7.n5051 net7.n5050 9.3
R26647 net7.n5039 net7.n5038 9.3
R26648 net7.n5037 net7.n5036 9.3
R26649 net7.n5240 net7.n5239 9.3
R26650 net7.n5121 net7.n5120 9.3
R26651 net7.n5123 net7.n5122 9.3
R26652 net7.n5132 net7.n5131 9.3
R26653 net7.n5114 net7.n5113 9.3
R26654 net7.n5116 net7.n5115 9.3
R26655 net7.n5227 net7.n5226 9.3
R26656 net7.n5269 net7.n5268 9.3
R26657 net7.n5253 net7.n5252 9.3
R26658 net7.n5242 net7.n5241 9.3
R26659 net7.n5229 net7.n5228 9.3
R26660 net7.n5283 net7.n5282 9.3
R26661 net7.n5285 net7.n5284 9.3
R26662 net7.n5413 net7.n5412 9.3
R26663 net7.n5401 net7.n5400 9.3
R26664 net7.n5399 net7.n5398 9.3
R26665 net7.n5602 net7.n5601 9.3
R26666 net7.n5483 net7.n5482 9.3
R26667 net7.n5485 net7.n5484 9.3
R26668 net7.n5494 net7.n5493 9.3
R26669 net7.n5476 net7.n5475 9.3
R26670 net7.n5478 net7.n5477 9.3
R26671 net7.n5589 net7.n5588 9.3
R26672 net7.n5631 net7.n5630 9.3
R26673 net7.n5615 net7.n5614 9.3
R26674 net7.n5604 net7.n5603 9.3
R26675 net7.n5591 net7.n5590 9.3
R26676 net7.n5645 net7.n5644 9.3
R26677 net7.n5647 net7.n5646 9.3
R26678 net7.n5775 net7.n5774 9.3
R26679 net7.n5763 net7.n5762 9.3
R26680 net7.n5761 net7.n5760 9.3
R26681 net7.n5964 net7.n5963 9.3
R26682 net7.n5845 net7.n5844 9.3
R26683 net7.n5847 net7.n5846 9.3
R26684 net7.n5856 net7.n5855 9.3
R26685 net7.n5838 net7.n5837 9.3
R26686 net7.n5840 net7.n5839 9.3
R26687 net7.n5951 net7.n5950 9.3
R26688 net7.n5993 net7.n5992 9.3
R26689 net7.n5977 net7.n5976 9.3
R26690 net7.n5966 net7.n5965 9.3
R26691 net7.n5953 net7.n5952 9.3
R26692 net7.n6007 net7.n6006 9.3
R26693 net7.n6009 net7.n6008 9.3
R26694 net7.n6137 net7.n6136 9.3
R26695 net7.n6125 net7.n6124 9.3
R26696 net7.n6123 net7.n6122 9.3
R26697 net7.n6326 net7.n6325 9.3
R26698 net7.n6207 net7.n6206 9.3
R26699 net7.n6209 net7.n6208 9.3
R26700 net7.n6218 net7.n6217 9.3
R26701 net7.n6200 net7.n6199 9.3
R26702 net7.n6202 net7.n6201 9.3
R26703 net7.n6313 net7.n6312 9.3
R26704 net7.n6355 net7.n6354 9.3
R26705 net7.n6339 net7.n6338 9.3
R26706 net7.n6328 net7.n6327 9.3
R26707 net7.n6315 net7.n6314 9.3
R26708 net7.n6369 net7.n6368 9.3
R26709 net7.n6371 net7.n6370 9.3
R26710 net7.n6499 net7.n6498 9.3
R26711 net7.n6487 net7.n6486 9.3
R26712 net7.n6485 net7.n6484 9.3
R26713 net7.n6688 net7.n6687 9.3
R26714 net7.n6569 net7.n6568 9.3
R26715 net7.n6571 net7.n6570 9.3
R26716 net7.n6580 net7.n6579 9.3
R26717 net7.n6562 net7.n6561 9.3
R26718 net7.n6564 net7.n6563 9.3
R26719 net7.n6675 net7.n6674 9.3
R26720 net7.n6717 net7.n6716 9.3
R26721 net7.n6701 net7.n6700 9.3
R26722 net7.n6690 net7.n6689 9.3
R26723 net7.n6677 net7.n6676 9.3
R26724 net7.n6731 net7.n6730 9.3
R26725 net7.n6733 net7.n6732 9.3
R26726 net7.n6861 net7.n6860 9.3
R26727 net7.n6849 net7.n6848 9.3
R26728 net7.n6847 net7.n6846 9.3
R26729 net7.n7050 net7.n7049 9.3
R26730 net7.n6931 net7.n6930 9.3
R26731 net7.n6933 net7.n6932 9.3
R26732 net7.n6942 net7.n6941 9.3
R26733 net7.n6924 net7.n6923 9.3
R26734 net7.n6926 net7.n6925 9.3
R26735 net7.n7037 net7.n7036 9.3
R26736 net7.n7079 net7.n7078 9.3
R26737 net7.n7063 net7.n7062 9.3
R26738 net7.n7052 net7.n7051 9.3
R26739 net7.n7039 net7.n7038 9.3
R26740 net7.n7093 net7.n7092 9.3
R26741 net7.n7095 net7.n7094 9.3
R26742 net7.n7223 net7.n7222 9.3
R26743 net7.n7211 net7.n7210 9.3
R26744 net7.n7209 net7.n7208 9.3
R26745 net7.n3693 net7.n3692 8.454
R26746 net7.n4054 net7.n4053 8.454
R26747 net7.n4416 net7.n4415 8.454
R26748 net7.n4778 net7.n4777 8.454
R26749 net7.n5140 net7.n5139 8.454
R26750 net7.n5502 net7.n5501 8.454
R26751 net7.n5864 net7.n5863 8.454
R26752 net7.n6226 net7.n6225 8.454
R26753 net7.n6588 net7.n6587 8.454
R26754 net7.n6950 net7.n6949 8.454
R26755 net7.n3309 net7.n3308 8.454
R26756 net7.n2947 net7.n2946 8.454
R26757 net7.n2585 net7.n2584 8.454
R26758 net7.n2223 net7.n2222 8.454
R26759 net7.n1861 net7.n1860 8.454
R26760 net7.n1499 net7.n1498 8.454
R26761 net7.n1137 net7.n1136 8.454
R26762 net7.n775 net7.n774 8.454
R26763 net7.n413 net7.n412 8.454
R26764 net7.n52 net7.n51 8.454
R26765 net7.n3610 net7.n3609 8.454
R26766 net7.n3248 net7.n3247 8.454
R26767 net7.n2886 net7.n2885 8.454
R26768 net7.n2524 net7.n2523 8.454
R26769 net7.n2162 net7.n2161 8.454
R26770 net7.n1800 net7.n1799 8.454
R26771 net7.n1438 net7.n1437 8.454
R26772 net7.n1076 net7.n1075 8.454
R26773 net7.n714 net7.n713 8.454
R26774 net7.n353 net7.n352 8.454
R26775 net7.n3977 net7.n3976 8.453
R26776 net7.n4338 net7.n4337 8.453
R26777 net7.n4700 net7.n4699 8.453
R26778 net7.n5062 net7.n5061 8.453
R26779 net7.n5424 net7.n5423 8.453
R26780 net7.n5786 net7.n5785 8.453
R26781 net7.n6148 net7.n6147 8.453
R26782 net7.n6510 net7.n6509 8.453
R26783 net7.n6872 net7.n6871 8.453
R26784 net7.n7234 net7.n7233 8.453
R26785 net7.n3540 net7.n3539 5.458
R26786 net7.n3178 net7.n3177 5.458
R26787 net7.n2816 net7.n2815 5.458
R26788 net7.n2454 net7.n2453 5.458
R26789 net7.n2092 net7.n2091 5.458
R26790 net7.n1730 net7.n1729 5.458
R26791 net7.n1368 net7.n1367 5.458
R26792 net7.n1006 net7.n1005 5.458
R26793 net7.n644 net7.n643 5.458
R26794 net7.n283 net7.n282 5.458
R26795 net7.n3792 net7.n3791 5.458
R26796 net7.n4153 net7.n4152 5.458
R26797 net7.n4515 net7.n4514 5.458
R26798 net7.n4877 net7.n4876 5.458
R26799 net7.n5239 net7.n5238 5.458
R26800 net7.n5601 net7.n5600 5.458
R26801 net7.n5963 net7.n5962 5.458
R26802 net7.n6325 net7.n6324 5.458
R26803 net7.n6687 net7.n6686 5.458
R26804 net7.n7049 net7.n7048 5.458
R26805 net7.n3411 net7.n3410 5.081
R26806 net7.n3049 net7.n3048 5.081
R26807 net7.n2687 net7.n2686 5.081
R26808 net7.n2325 net7.n2324 5.081
R26809 net7.n1963 net7.n1962 5.081
R26810 net7.n1601 net7.n1600 5.081
R26811 net7.n1239 net7.n1238 5.081
R26812 net7.n877 net7.n876 5.081
R26813 net7.n515 net7.n514 5.081
R26814 net7.n154 net7.n153 5.081
R26815 net7.n3835 net7.n3834 5.081
R26816 net7.n4196 net7.n4195 5.081
R26817 net7.n4558 net7.n4557 5.081
R26818 net7.n4920 net7.n4919 5.081
R26819 net7.n5282 net7.n5281 5.081
R26820 net7.n5644 net7.n5643 5.081
R26821 net7.n6006 net7.n6005 5.081
R26822 net7.n6368 net7.n6367 5.081
R26823 net7.n6730 net7.n6729 5.081
R26824 net7.n7092 net7.n7091 5.081
R26825 net7.n3277 net7.n3276 4.65
R26826 net7.n3404 net7.n3403 4.65
R26827 net7.n2915 net7.n2914 4.65
R26828 net7.n3042 net7.n3041 4.65
R26829 net7.n2553 net7.n2552 4.65
R26830 net7.n2680 net7.n2679 4.65
R26831 net7.n2191 net7.n2190 4.65
R26832 net7.n2318 net7.n2317 4.65
R26833 net7.n1829 net7.n1828 4.65
R26834 net7.n1956 net7.n1955 4.65
R26835 net7.n1467 net7.n1466 4.65
R26836 net7.n1594 net7.n1593 4.65
R26837 net7.n1105 net7.n1104 4.65
R26838 net7.n1232 net7.n1231 4.65
R26839 net7.n743 net7.n742 4.65
R26840 net7.n870 net7.n869 4.65
R26841 net7.n381 net7.n380 4.65
R26842 net7.n508 net7.n507 4.65
R26843 net7.n20 net7.n19 4.65
R26844 net7.n147 net7.n146 4.65
R26845 net7.n3944 net7.n3943 4.65
R26846 net7.n3912 net7.n3911 4.65
R26847 net7.n4305 net7.n4304 4.65
R26848 net7.n4273 net7.n4272 4.65
R26849 net7.n4667 net7.n4666 4.65
R26850 net7.n4635 net7.n4634 4.65
R26851 net7.n5029 net7.n5028 4.65
R26852 net7.n4997 net7.n4996 4.65
R26853 net7.n5391 net7.n5390 4.65
R26854 net7.n5359 net7.n5358 4.65
R26855 net7.n5753 net7.n5752 4.65
R26856 net7.n5721 net7.n5720 4.65
R26857 net7.n6115 net7.n6114 4.65
R26858 net7.n6083 net7.n6082 4.65
R26859 net7.n6477 net7.n6476 4.65
R26860 net7.n6445 net7.n6444 4.65
R26861 net7.n6839 net7.n6838 4.65
R26862 net7.n6807 net7.n6806 4.65
R26863 net7.n7201 net7.n7200 4.65
R26864 net7.n7169 net7.n7168 4.65
R26865 net7.n3292 net7.n3291 4.5
R26866 net7.n3568 net7.n3567 4.5
R26867 net7.n3562 net7.n3519 4.5
R26868 net7.n3574 net7.n3515 4.5
R26869 net7.n3584 net7.n3583 4.5
R26870 net7.n3603 net7.n3602 4.5
R26871 net7.n3592 net7.n3512 4.5
R26872 net7.n3558 net7.n3557 4.5
R26873 net7.n3545 net7.n3521 4.5
R26874 net7.n3535 net7.n3534 4.5
R26875 net7.n3525 net7.n3523 4.5
R26876 net7.n3380 net7.n3379 4.5
R26877 net7.n3417 net7.n3416 4.5
R26878 net7.n3398 net7.n3389 4.5
R26879 net7.n3346 net7.n3343 4.5
R26880 net7.n3394 net7.n3393 4.5
R26881 net7.n3273 net7.n3272 4.5
R26882 net7.n3303 net7.n3302 4.5
R26883 net7.n2930 net7.n2929 4.5
R26884 net7.n3206 net7.n3205 4.5
R26885 net7.n3200 net7.n3157 4.5
R26886 net7.n3212 net7.n3153 4.5
R26887 net7.n3222 net7.n3221 4.5
R26888 net7.n3241 net7.n3240 4.5
R26889 net7.n3230 net7.n3150 4.5
R26890 net7.n3196 net7.n3195 4.5
R26891 net7.n3183 net7.n3159 4.5
R26892 net7.n3173 net7.n3172 4.5
R26893 net7.n3163 net7.n3161 4.5
R26894 net7.n3018 net7.n3017 4.5
R26895 net7.n3055 net7.n3054 4.5
R26896 net7.n3036 net7.n3027 4.5
R26897 net7.n2984 net7.n2981 4.5
R26898 net7.n3032 net7.n3031 4.5
R26899 net7.n2911 net7.n2910 4.5
R26900 net7.n2941 net7.n2940 4.5
R26901 net7.n2568 net7.n2567 4.5
R26902 net7.n2844 net7.n2843 4.5
R26903 net7.n2838 net7.n2795 4.5
R26904 net7.n2850 net7.n2791 4.5
R26905 net7.n2860 net7.n2859 4.5
R26906 net7.n2879 net7.n2878 4.5
R26907 net7.n2868 net7.n2788 4.5
R26908 net7.n2834 net7.n2833 4.5
R26909 net7.n2821 net7.n2797 4.5
R26910 net7.n2811 net7.n2810 4.5
R26911 net7.n2801 net7.n2799 4.5
R26912 net7.n2656 net7.n2655 4.5
R26913 net7.n2693 net7.n2692 4.5
R26914 net7.n2674 net7.n2665 4.5
R26915 net7.n2622 net7.n2619 4.5
R26916 net7.n2670 net7.n2669 4.5
R26917 net7.n2549 net7.n2548 4.5
R26918 net7.n2579 net7.n2578 4.5
R26919 net7.n2206 net7.n2205 4.5
R26920 net7.n2482 net7.n2481 4.5
R26921 net7.n2476 net7.n2433 4.5
R26922 net7.n2488 net7.n2429 4.5
R26923 net7.n2498 net7.n2497 4.5
R26924 net7.n2517 net7.n2516 4.5
R26925 net7.n2506 net7.n2426 4.5
R26926 net7.n2472 net7.n2471 4.5
R26927 net7.n2459 net7.n2435 4.5
R26928 net7.n2449 net7.n2448 4.5
R26929 net7.n2439 net7.n2437 4.5
R26930 net7.n2294 net7.n2293 4.5
R26931 net7.n2331 net7.n2330 4.5
R26932 net7.n2312 net7.n2303 4.5
R26933 net7.n2260 net7.n2257 4.5
R26934 net7.n2308 net7.n2307 4.5
R26935 net7.n2187 net7.n2186 4.5
R26936 net7.n2217 net7.n2216 4.5
R26937 net7.n1844 net7.n1843 4.5
R26938 net7.n2120 net7.n2119 4.5
R26939 net7.n2114 net7.n2071 4.5
R26940 net7.n2126 net7.n2067 4.5
R26941 net7.n2136 net7.n2135 4.5
R26942 net7.n2155 net7.n2154 4.5
R26943 net7.n2144 net7.n2064 4.5
R26944 net7.n2110 net7.n2109 4.5
R26945 net7.n2097 net7.n2073 4.5
R26946 net7.n2087 net7.n2086 4.5
R26947 net7.n2077 net7.n2075 4.5
R26948 net7.n1932 net7.n1931 4.5
R26949 net7.n1969 net7.n1968 4.5
R26950 net7.n1950 net7.n1941 4.5
R26951 net7.n1898 net7.n1895 4.5
R26952 net7.n1946 net7.n1945 4.5
R26953 net7.n1825 net7.n1824 4.5
R26954 net7.n1855 net7.n1854 4.5
R26955 net7.n1482 net7.n1481 4.5
R26956 net7.n1758 net7.n1757 4.5
R26957 net7.n1752 net7.n1709 4.5
R26958 net7.n1764 net7.n1705 4.5
R26959 net7.n1774 net7.n1773 4.5
R26960 net7.n1793 net7.n1792 4.5
R26961 net7.n1782 net7.n1702 4.5
R26962 net7.n1748 net7.n1747 4.5
R26963 net7.n1735 net7.n1711 4.5
R26964 net7.n1725 net7.n1724 4.5
R26965 net7.n1715 net7.n1713 4.5
R26966 net7.n1570 net7.n1569 4.5
R26967 net7.n1607 net7.n1606 4.5
R26968 net7.n1588 net7.n1579 4.5
R26969 net7.n1536 net7.n1533 4.5
R26970 net7.n1584 net7.n1583 4.5
R26971 net7.n1463 net7.n1462 4.5
R26972 net7.n1493 net7.n1492 4.5
R26973 net7.n1120 net7.n1119 4.5
R26974 net7.n1396 net7.n1395 4.5
R26975 net7.n1390 net7.n1347 4.5
R26976 net7.n1402 net7.n1343 4.5
R26977 net7.n1412 net7.n1411 4.5
R26978 net7.n1431 net7.n1430 4.5
R26979 net7.n1420 net7.n1340 4.5
R26980 net7.n1386 net7.n1385 4.5
R26981 net7.n1373 net7.n1349 4.5
R26982 net7.n1363 net7.n1362 4.5
R26983 net7.n1353 net7.n1351 4.5
R26984 net7.n1208 net7.n1207 4.5
R26985 net7.n1245 net7.n1244 4.5
R26986 net7.n1226 net7.n1217 4.5
R26987 net7.n1174 net7.n1171 4.5
R26988 net7.n1222 net7.n1221 4.5
R26989 net7.n1101 net7.n1100 4.5
R26990 net7.n1131 net7.n1130 4.5
R26991 net7.n758 net7.n757 4.5
R26992 net7.n1034 net7.n1033 4.5
R26993 net7.n1028 net7.n985 4.5
R26994 net7.n1040 net7.n981 4.5
R26995 net7.n1050 net7.n1049 4.5
R26996 net7.n1069 net7.n1068 4.5
R26997 net7.n1058 net7.n978 4.5
R26998 net7.n1024 net7.n1023 4.5
R26999 net7.n1011 net7.n987 4.5
R27000 net7.n1001 net7.n1000 4.5
R27001 net7.n991 net7.n989 4.5
R27002 net7.n846 net7.n845 4.5
R27003 net7.n883 net7.n882 4.5
R27004 net7.n864 net7.n855 4.5
R27005 net7.n812 net7.n809 4.5
R27006 net7.n860 net7.n859 4.5
R27007 net7.n739 net7.n738 4.5
R27008 net7.n769 net7.n768 4.5
R27009 net7.n396 net7.n395 4.5
R27010 net7.n672 net7.n671 4.5
R27011 net7.n666 net7.n623 4.5
R27012 net7.n678 net7.n619 4.5
R27013 net7.n688 net7.n687 4.5
R27014 net7.n707 net7.n706 4.5
R27015 net7.n696 net7.n616 4.5
R27016 net7.n662 net7.n661 4.5
R27017 net7.n649 net7.n625 4.5
R27018 net7.n639 net7.n638 4.5
R27019 net7.n629 net7.n627 4.5
R27020 net7.n484 net7.n483 4.5
R27021 net7.n521 net7.n520 4.5
R27022 net7.n502 net7.n493 4.5
R27023 net7.n450 net7.n447 4.5
R27024 net7.n498 net7.n497 4.5
R27025 net7.n377 net7.n376 4.5
R27026 net7.n407 net7.n406 4.5
R27027 net7.n35 net7.n34 4.5
R27028 net7.n311 net7.n310 4.5
R27029 net7.n305 net7.n262 4.5
R27030 net7.n317 net7.n258 4.5
R27031 net7.n327 net7.n326 4.5
R27032 net7.n335 net7.n255 4.5
R27033 net7.n301 net7.n300 4.5
R27034 net7.n288 net7.n264 4.5
R27035 net7.n278 net7.n277 4.5
R27036 net7.n268 net7.n266 4.5
R27037 net7.n123 net7.n122 4.5
R27038 net7.n160 net7.n159 4.5
R27039 net7.n141 net7.n132 4.5
R27040 net7.n89 net7.n86 4.5
R27041 net7.n137 net7.n136 4.5
R27042 net7.n16 net7.n15 4.5
R27043 net7.n46 net7.n45 4.5
R27044 net7.n346 net7.n345 4.5
R27045 net7.n3959 net7.n3958 4.5
R27046 net7.n3940 net7.n3939 4.5
R27047 net7.n3932 net7.n3931 4.5
R27048 net7.n3918 net7.n3917 4.5
R27049 net7.n3839 net7.n3827 4.5
R27050 net7.n3819 net7.n3818 4.5
R27051 net7.n3809 net7.n3808 4.5
R27052 net7.n3799 net7.n3798 4.5
R27053 net7.n3787 net7.n3786 4.5
R27054 net7.n3670 net7.n3636 4.5
R27055 net7.n3663 net7.n3639 4.5
R27056 net7.n3678 net7.n3633 4.5
R27057 net7.n3687 net7.n3630 4.5
R27058 net7.n3657 net7.n3642 4.5
R27059 net7.n3654 net7.n3646 4.5
R27060 net7.n3650 net7.n3649 4.5
R27061 net7.n3926 net7.n3925 4.5
R27062 net7.n3970 net7.n3969 4.5
R27063 net7.n4320 net7.n4319 4.5
R27064 net7.n4301 net7.n4300 4.5
R27065 net7.n4293 net7.n4292 4.5
R27066 net7.n4279 net7.n4278 4.5
R27067 net7.n4200 net7.n4188 4.5
R27068 net7.n4180 net7.n4179 4.5
R27069 net7.n4170 net7.n4169 4.5
R27070 net7.n4160 net7.n4159 4.5
R27071 net7.n4148 net7.n4147 4.5
R27072 net7.n4031 net7.n3997 4.5
R27073 net7.n4024 net7.n4000 4.5
R27074 net7.n4039 net7.n3994 4.5
R27075 net7.n4048 net7.n3991 4.5
R27076 net7.n4018 net7.n4003 4.5
R27077 net7.n4015 net7.n4007 4.5
R27078 net7.n4011 net7.n4010 4.5
R27079 net7.n4287 net7.n4286 4.5
R27080 net7.n4331 net7.n4330 4.5
R27081 net7.n4682 net7.n4681 4.5
R27082 net7.n4663 net7.n4662 4.5
R27083 net7.n4655 net7.n4654 4.5
R27084 net7.n4641 net7.n4640 4.5
R27085 net7.n4562 net7.n4550 4.5
R27086 net7.n4542 net7.n4541 4.5
R27087 net7.n4532 net7.n4531 4.5
R27088 net7.n4522 net7.n4521 4.5
R27089 net7.n4510 net7.n4509 4.5
R27090 net7.n4393 net7.n4359 4.5
R27091 net7.n4386 net7.n4362 4.5
R27092 net7.n4401 net7.n4356 4.5
R27093 net7.n4410 net7.n4353 4.5
R27094 net7.n4380 net7.n4365 4.5
R27095 net7.n4377 net7.n4369 4.5
R27096 net7.n4373 net7.n4372 4.5
R27097 net7.n4649 net7.n4648 4.5
R27098 net7.n4693 net7.n4692 4.5
R27099 net7.n5044 net7.n5043 4.5
R27100 net7.n5025 net7.n5024 4.5
R27101 net7.n5017 net7.n5016 4.5
R27102 net7.n5003 net7.n5002 4.5
R27103 net7.n4924 net7.n4912 4.5
R27104 net7.n4904 net7.n4903 4.5
R27105 net7.n4894 net7.n4893 4.5
R27106 net7.n4884 net7.n4883 4.5
R27107 net7.n4872 net7.n4871 4.5
R27108 net7.n4755 net7.n4721 4.5
R27109 net7.n4748 net7.n4724 4.5
R27110 net7.n4763 net7.n4718 4.5
R27111 net7.n4772 net7.n4715 4.5
R27112 net7.n4742 net7.n4727 4.5
R27113 net7.n4739 net7.n4731 4.5
R27114 net7.n4735 net7.n4734 4.5
R27115 net7.n5011 net7.n5010 4.5
R27116 net7.n5055 net7.n5054 4.5
R27117 net7.n5406 net7.n5405 4.5
R27118 net7.n5387 net7.n5386 4.5
R27119 net7.n5379 net7.n5378 4.5
R27120 net7.n5365 net7.n5364 4.5
R27121 net7.n5286 net7.n5274 4.5
R27122 net7.n5266 net7.n5265 4.5
R27123 net7.n5256 net7.n5255 4.5
R27124 net7.n5246 net7.n5245 4.5
R27125 net7.n5234 net7.n5233 4.5
R27126 net7.n5117 net7.n5083 4.5
R27127 net7.n5110 net7.n5086 4.5
R27128 net7.n5125 net7.n5080 4.5
R27129 net7.n5134 net7.n5077 4.5
R27130 net7.n5104 net7.n5089 4.5
R27131 net7.n5101 net7.n5093 4.5
R27132 net7.n5097 net7.n5096 4.5
R27133 net7.n5373 net7.n5372 4.5
R27134 net7.n5417 net7.n5416 4.5
R27135 net7.n5768 net7.n5767 4.5
R27136 net7.n5749 net7.n5748 4.5
R27137 net7.n5741 net7.n5740 4.5
R27138 net7.n5727 net7.n5726 4.5
R27139 net7.n5648 net7.n5636 4.5
R27140 net7.n5628 net7.n5627 4.5
R27141 net7.n5618 net7.n5617 4.5
R27142 net7.n5608 net7.n5607 4.5
R27143 net7.n5596 net7.n5595 4.5
R27144 net7.n5479 net7.n5445 4.5
R27145 net7.n5472 net7.n5448 4.5
R27146 net7.n5487 net7.n5442 4.5
R27147 net7.n5496 net7.n5439 4.5
R27148 net7.n5466 net7.n5451 4.5
R27149 net7.n5463 net7.n5455 4.5
R27150 net7.n5459 net7.n5458 4.5
R27151 net7.n5735 net7.n5734 4.5
R27152 net7.n5779 net7.n5778 4.5
R27153 net7.n6130 net7.n6129 4.5
R27154 net7.n6111 net7.n6110 4.5
R27155 net7.n6103 net7.n6102 4.5
R27156 net7.n6089 net7.n6088 4.5
R27157 net7.n6010 net7.n5998 4.5
R27158 net7.n5990 net7.n5989 4.5
R27159 net7.n5980 net7.n5979 4.5
R27160 net7.n5970 net7.n5969 4.5
R27161 net7.n5958 net7.n5957 4.5
R27162 net7.n5841 net7.n5807 4.5
R27163 net7.n5834 net7.n5810 4.5
R27164 net7.n5849 net7.n5804 4.5
R27165 net7.n5858 net7.n5801 4.5
R27166 net7.n5828 net7.n5813 4.5
R27167 net7.n5825 net7.n5817 4.5
R27168 net7.n5821 net7.n5820 4.5
R27169 net7.n6097 net7.n6096 4.5
R27170 net7.n6141 net7.n6140 4.5
R27171 net7.n6492 net7.n6491 4.5
R27172 net7.n6473 net7.n6472 4.5
R27173 net7.n6465 net7.n6464 4.5
R27174 net7.n6451 net7.n6450 4.5
R27175 net7.n6372 net7.n6360 4.5
R27176 net7.n6352 net7.n6351 4.5
R27177 net7.n6342 net7.n6341 4.5
R27178 net7.n6332 net7.n6331 4.5
R27179 net7.n6320 net7.n6319 4.5
R27180 net7.n6203 net7.n6169 4.5
R27181 net7.n6196 net7.n6172 4.5
R27182 net7.n6211 net7.n6166 4.5
R27183 net7.n6220 net7.n6163 4.5
R27184 net7.n6190 net7.n6175 4.5
R27185 net7.n6187 net7.n6179 4.5
R27186 net7.n6183 net7.n6182 4.5
R27187 net7.n6459 net7.n6458 4.5
R27188 net7.n6503 net7.n6502 4.5
R27189 net7.n6854 net7.n6853 4.5
R27190 net7.n6835 net7.n6834 4.5
R27191 net7.n6827 net7.n6826 4.5
R27192 net7.n6813 net7.n6812 4.5
R27193 net7.n6734 net7.n6722 4.5
R27194 net7.n6714 net7.n6713 4.5
R27195 net7.n6704 net7.n6703 4.5
R27196 net7.n6694 net7.n6693 4.5
R27197 net7.n6682 net7.n6681 4.5
R27198 net7.n6565 net7.n6531 4.5
R27199 net7.n6558 net7.n6534 4.5
R27200 net7.n6573 net7.n6528 4.5
R27201 net7.n6582 net7.n6525 4.5
R27202 net7.n6552 net7.n6537 4.5
R27203 net7.n6549 net7.n6541 4.5
R27204 net7.n6545 net7.n6544 4.5
R27205 net7.n6821 net7.n6820 4.5
R27206 net7.n6865 net7.n6864 4.5
R27207 net7.n7216 net7.n7215 4.5
R27208 net7.n7197 net7.n7196 4.5
R27209 net7.n7189 net7.n7188 4.5
R27210 net7.n7175 net7.n7174 4.5
R27211 net7.n7096 net7.n7084 4.5
R27212 net7.n7076 net7.n7075 4.5
R27213 net7.n7066 net7.n7065 4.5
R27214 net7.n7056 net7.n7055 4.5
R27215 net7.n7044 net7.n7043 4.5
R27216 net7.n6927 net7.n6893 4.5
R27217 net7.n6920 net7.n6896 4.5
R27218 net7.n6935 net7.n6890 4.5
R27219 net7.n6944 net7.n6887 4.5
R27220 net7.n6914 net7.n6899 4.5
R27221 net7.n6911 net7.n6903 4.5
R27222 net7.n6907 net7.n6906 4.5
R27223 net7.n7183 net7.n7182 4.5
R27224 net7.n7227 net7.n7226 4.5
R27225 net7.n3515 net7.n3513 4.325
R27226 net7.n3153 net7.n3151 4.325
R27227 net7.n2791 net7.n2789 4.325
R27228 net7.n2429 net7.n2427 4.325
R27229 net7.n2067 net7.n2065 4.325
R27230 net7.n1705 net7.n1703 4.325
R27231 net7.n1343 net7.n1341 4.325
R27232 net7.n981 net7.n979 4.325
R27233 net7.n619 net7.n617 4.325
R27234 net7.n258 net7.n256 4.325
R27235 net7.n3639 net7.n3637 4.325
R27236 net7.n4000 net7.n3998 4.325
R27237 net7.n4362 net7.n4360 4.325
R27238 net7.n4724 net7.n4722 4.325
R27239 net7.n5086 net7.n5084 4.325
R27240 net7.n5448 net7.n5446 4.325
R27241 net7.n5810 net7.n5808 4.325
R27242 net7.n6172 net7.n6170 4.325
R27243 net7.n6534 net7.n6532 4.325
R27244 net7.n6896 net7.n6894 4.325
R27245 net7.n3608 net7.t9 4.289
R27246 net7.n3246 net7.t6 4.289
R27247 net7.n2884 net7.t8 4.289
R27248 net7.n2522 net7.t7 4.289
R27249 net7.n2160 net7.t4 4.289
R27250 net7.n1798 net7.t2 4.289
R27251 net7.n1436 net7.t5 4.289
R27252 net7.n1074 net7.t3 4.289
R27253 net7.n712 net7.t0 4.289
R27254 net7.n351 net7.t1 4.289
R27255 net7.n3975 net7.t10 4.289
R27256 net7.n4336 net7.t16 4.289
R27257 net7.n4698 net7.t11 4.289
R27258 net7.n5060 net7.t12 4.289
R27259 net7.n5422 net7.t17 4.289
R27260 net7.n5784 net7.t18 4.289
R27261 net7.n6146 net7.t13 4.289
R27262 net7.n6508 net7.t14 4.289
R27263 net7.n6870 net7.t19 4.289
R27264 net7.n7232 net7.t15 4.289
R27265 net7.n3519 net7.n3516 3.95
R27266 net7.n3157 net7.n3154 3.95
R27267 net7.n2795 net7.n2792 3.95
R27268 net7.n2433 net7.n2430 3.95
R27269 net7.n2071 net7.n2068 3.95
R27270 net7.n1709 net7.n1706 3.95
R27271 net7.n1347 net7.n1344 3.95
R27272 net7.n985 net7.n982 3.95
R27273 net7.n623 net7.n620 3.95
R27274 net7.n262 net7.n259 3.95
R27275 net7.n3646 net7.n3643 3.95
R27276 net7.n4007 net7.n4004 3.95
R27277 net7.n4369 net7.n4366 3.95
R27278 net7.n4731 net7.n4728 3.95
R27279 net7.n5093 net7.n5090 3.95
R27280 net7.n5455 net7.n5452 3.95
R27281 net7.n5817 net7.n5814 3.95
R27282 net7.n6179 net7.n6176 3.95
R27283 net7.n6541 net7.n6538 3.95
R27284 net7.n6903 net7.n6900 3.95
R27285 net7.n3272 net7.n3271 3.948
R27286 net7.n2910 net7.n2909 3.948
R27287 net7.n2548 net7.n2547 3.948
R27288 net7.n2186 net7.n2185 3.948
R27289 net7.n1824 net7.n1823 3.948
R27290 net7.n1462 net7.n1461 3.948
R27291 net7.n1100 net7.n1099 3.948
R27292 net7.n738 net7.n737 3.948
R27293 net7.n376 net7.n375 3.948
R27294 net7.n15 net7.n14 3.948
R27295 net7.n3939 net7.n3938 3.948
R27296 net7.n4300 net7.n4299 3.948
R27297 net7.n4662 net7.n4661 3.948
R27298 net7.n5024 net7.n5023 3.948
R27299 net7.n5386 net7.n5385 3.948
R27300 net7.n5748 net7.n5747 3.948
R27301 net7.n6110 net7.n6109 3.948
R27302 net7.n6472 net7.n6471 3.948
R27303 net7.n6834 net7.n6833 3.948
R27304 net7.n7196 net7.n7195 3.948
R27305 net7.n3393 net7.n3392 3.573
R27306 net7.n3031 net7.n3030 3.573
R27307 net7.n2669 net7.n2668 3.573
R27308 net7.n2307 net7.n2306 3.573
R27309 net7.n1945 net7.n1944 3.573
R27310 net7.n1583 net7.n1582 3.573
R27311 net7.n1221 net7.n1220 3.573
R27312 net7.n859 net7.n858 3.573
R27313 net7.n497 net7.n496 3.573
R27314 net7.n136 net7.n135 3.573
R27315 net7.n3925 net7.n3924 3.573
R27316 net7.n4286 net7.n4285 3.573
R27317 net7.n4648 net7.n4647 3.573
R27318 net7.n5010 net7.n5009 3.573
R27319 net7.n5372 net7.n5371 3.573
R27320 net7.n5734 net7.n5733 3.573
R27321 net7.n6096 net7.n6095 3.573
R27322 net7.n6458 net7.n6457 3.573
R27323 net7.n6820 net7.n6819 3.573
R27324 net7.n7182 net7.n7181 3.573
R27325 net7.n3406 net7.n3387 3.033
R27326 net7.n3281 net7.n3280 3.033
R27327 net7.n3044 net7.n3025 3.033
R27328 net7.n2919 net7.n2918 3.033
R27329 net7.n2682 net7.n2663 3.033
R27330 net7.n2557 net7.n2556 3.033
R27331 net7.n2320 net7.n2301 3.033
R27332 net7.n2195 net7.n2194 3.033
R27333 net7.n1958 net7.n1939 3.033
R27334 net7.n1833 net7.n1832 3.033
R27335 net7.n1596 net7.n1577 3.033
R27336 net7.n1471 net7.n1470 3.033
R27337 net7.n1234 net7.n1215 3.033
R27338 net7.n1109 net7.n1108 3.033
R27339 net7.n872 net7.n853 3.033
R27340 net7.n747 net7.n746 3.033
R27341 net7.n510 net7.n491 3.033
R27342 net7.n385 net7.n384 3.033
R27343 net7.n149 net7.n130 3.033
R27344 net7.n24 net7.n23 3.033
R27345 net7.n3830 net7.n3828 3.033
R27346 net7.n3948 net7.n3947 3.033
R27347 net7.n4191 net7.n4189 3.033
R27348 net7.n4309 net7.n4308 3.033
R27349 net7.n4553 net7.n4551 3.033
R27350 net7.n4671 net7.n4670 3.033
R27351 net7.n4915 net7.n4913 3.033
R27352 net7.n5033 net7.n5032 3.033
R27353 net7.n5277 net7.n5275 3.033
R27354 net7.n5395 net7.n5394 3.033
R27355 net7.n5639 net7.n5637 3.033
R27356 net7.n5757 net7.n5756 3.033
R27357 net7.n6001 net7.n5999 3.033
R27358 net7.n6119 net7.n6118 3.033
R27359 net7.n6363 net7.n6361 3.033
R27360 net7.n6481 net7.n6480 3.033
R27361 net7.n6725 net7.n6723 3.033
R27362 net7.n6843 net7.n6842 3.033
R27363 net7.n7087 net7.n7085 3.033
R27364 net7.n7205 net7.n7204 3.033
R27365 net7.n3518 net7.n3517 2.258
R27366 net7.n3391 net7.n3390 2.258
R27367 net7.n3156 net7.n3155 2.258
R27368 net7.n3029 net7.n3028 2.258
R27369 net7.n2794 net7.n2793 2.258
R27370 net7.n2667 net7.n2666 2.258
R27371 net7.n2432 net7.n2431 2.258
R27372 net7.n2305 net7.n2304 2.258
R27373 net7.n2070 net7.n2069 2.258
R27374 net7.n1943 net7.n1942 2.258
R27375 net7.n1708 net7.n1707 2.258
R27376 net7.n1581 net7.n1580 2.258
R27377 net7.n1346 net7.n1345 2.258
R27378 net7.n1219 net7.n1218 2.258
R27379 net7.n984 net7.n983 2.258
R27380 net7.n857 net7.n856 2.258
R27381 net7.n622 net7.n621 2.258
R27382 net7.n495 net7.n494 2.258
R27383 net7.n261 net7.n260 2.258
R27384 net7.n134 net7.n133 2.258
R27385 net7.n3645 net7.n3644 2.258
R27386 net7.n3923 net7.n3922 2.258
R27387 net7.n4006 net7.n4005 2.258
R27388 net7.n4284 net7.n4283 2.258
R27389 net7.n4368 net7.n4367 2.258
R27390 net7.n4646 net7.n4645 2.258
R27391 net7.n4730 net7.n4729 2.258
R27392 net7.n5008 net7.n5007 2.258
R27393 net7.n5092 net7.n5091 2.258
R27394 net7.n5370 net7.n5369 2.258
R27395 net7.n5454 net7.n5453 2.258
R27396 net7.n5732 net7.n5731 2.258
R27397 net7.n5816 net7.n5815 2.258
R27398 net7.n6094 net7.n6093 2.258
R27399 net7.n6178 net7.n6177 2.258
R27400 net7.n6456 net7.n6455 2.258
R27401 net7.n6540 net7.n6539 2.258
R27402 net7.n6818 net7.n6817 2.258
R27403 net7.n6902 net7.n6901 2.258
R27404 net7.n7180 net7.n7179 2.258
R27405 net7.n722 net7.n360 2.089
R27406 net7.n3618 net7.n3617 2.031
R27407 net7.n2894 net7.n2893 2.031
R27408 net7.n2170 net7.n2169 2.031
R27409 net7.n1446 net7.n1445 2.031
R27410 net7.n722 net7.n721 2.031
R27411 net7.n3256 net7.n3255 2.03
R27412 net7.n2532 net7.n2531 2.03
R27413 net7.n1808 net7.n1807 2.03
R27414 net7.n1084 net7.n1083 2.03
R27415 net7.n3566 net7.n3565 1.882
R27416 net7.n3567 net7.n3566 1.882
R27417 net7.n3342 net7.n3341 1.882
R27418 net7.n3204 net7.n3203 1.882
R27419 net7.n3205 net7.n3204 1.882
R27420 net7.n2980 net7.n2979 1.882
R27421 net7.n2842 net7.n2841 1.882
R27422 net7.n2843 net7.n2842 1.882
R27423 net7.n2618 net7.n2617 1.882
R27424 net7.n2480 net7.n2479 1.882
R27425 net7.n2481 net7.n2480 1.882
R27426 net7.n2256 net7.n2255 1.882
R27427 net7.n2118 net7.n2117 1.882
R27428 net7.n2119 net7.n2118 1.882
R27429 net7.n1894 net7.n1893 1.882
R27430 net7.n1756 net7.n1755 1.882
R27431 net7.n1757 net7.n1756 1.882
R27432 net7.n1532 net7.n1531 1.882
R27433 net7.n1394 net7.n1393 1.882
R27434 net7.n1395 net7.n1394 1.882
R27435 net7.n1170 net7.n1169 1.882
R27436 net7.n1032 net7.n1031 1.882
R27437 net7.n1033 net7.n1032 1.882
R27438 net7.n808 net7.n807 1.882
R27439 net7.n670 net7.n669 1.882
R27440 net7.n671 net7.n670 1.882
R27441 net7.n446 net7.n445 1.882
R27442 net7.n309 net7.n308 1.882
R27443 net7.n310 net7.n309 1.882
R27444 net7.n85 net7.n84 1.882
R27445 net7.n3641 net7.n3640 1.882
R27446 net7.n3642 net7.n3641 1.882
R27447 net7.n3930 net7.n3929 1.882
R27448 net7.n4002 net7.n4001 1.882
R27449 net7.n4003 net7.n4002 1.882
R27450 net7.n4291 net7.n4290 1.882
R27451 net7.n4364 net7.n4363 1.882
R27452 net7.n4365 net7.n4364 1.882
R27453 net7.n4653 net7.n4652 1.882
R27454 net7.n4726 net7.n4725 1.882
R27455 net7.n4727 net7.n4726 1.882
R27456 net7.n5015 net7.n5014 1.882
R27457 net7.n5088 net7.n5087 1.882
R27458 net7.n5089 net7.n5088 1.882
R27459 net7.n5377 net7.n5376 1.882
R27460 net7.n5450 net7.n5449 1.882
R27461 net7.n5451 net7.n5450 1.882
R27462 net7.n5739 net7.n5738 1.882
R27463 net7.n5812 net7.n5811 1.882
R27464 net7.n5813 net7.n5812 1.882
R27465 net7.n6101 net7.n6100 1.882
R27466 net7.n6174 net7.n6173 1.882
R27467 net7.n6175 net7.n6174 1.882
R27468 net7.n6463 net7.n6462 1.882
R27469 net7.n6536 net7.n6535 1.882
R27470 net7.n6537 net7.n6536 1.882
R27471 net7.n6825 net7.n6824 1.882
R27472 net7.n6898 net7.n6897 1.882
R27473 net7.n6899 net7.n6898 1.882
R27474 net7.n7187 net7.n7186 1.882
R27475 net7.n3609 net7.n3608 1.844
R27476 net7.n3247 net7.n3246 1.844
R27477 net7.n2885 net7.n2884 1.844
R27478 net7.n2523 net7.n2522 1.844
R27479 net7.n2161 net7.n2160 1.844
R27480 net7.n1799 net7.n1798 1.844
R27481 net7.n1437 net7.n1436 1.844
R27482 net7.n1075 net7.n1074 1.844
R27483 net7.n713 net7.n712 1.844
R27484 net7.n352 net7.n351 1.844
R27485 net7.n3976 net7.n3975 1.844
R27486 net7.n4337 net7.n4336 1.844
R27487 net7.n4699 net7.n4698 1.844
R27488 net7.n5061 net7.n5060 1.844
R27489 net7.n5423 net7.n5422 1.844
R27490 net7.n5785 net7.n5784 1.844
R27491 net7.n6147 net7.n6146 1.844
R27492 net7.n6509 net7.n6508 1.844
R27493 net7.n6871 net7.n6870 1.844
R27494 net7.n7233 net7.n7232 1.844
R27495 net7.n3393 net7.n3391 1.505
R27496 net7.n3343 net7.n3342 1.505
R27497 net7.n3031 net7.n3029 1.505
R27498 net7.n2981 net7.n2980 1.505
R27499 net7.n2669 net7.n2667 1.505
R27500 net7.n2619 net7.n2618 1.505
R27501 net7.n2307 net7.n2305 1.505
R27502 net7.n2257 net7.n2256 1.505
R27503 net7.n1945 net7.n1943 1.505
R27504 net7.n1895 net7.n1894 1.505
R27505 net7.n1583 net7.n1581 1.505
R27506 net7.n1533 net7.n1532 1.505
R27507 net7.n1221 net7.n1219 1.505
R27508 net7.n1171 net7.n1170 1.505
R27509 net7.n859 net7.n857 1.505
R27510 net7.n809 net7.n808 1.505
R27511 net7.n497 net7.n495 1.505
R27512 net7.n447 net7.n446 1.505
R27513 net7.n136 net7.n134 1.505
R27514 net7.n86 net7.n85 1.505
R27515 net7.n3925 net7.n3923 1.505
R27516 net7.n3931 net7.n3930 1.505
R27517 net7.n4286 net7.n4284 1.505
R27518 net7.n4292 net7.n4291 1.505
R27519 net7.n4648 net7.n4646 1.505
R27520 net7.n4654 net7.n4653 1.505
R27521 net7.n5010 net7.n5008 1.505
R27522 net7.n5016 net7.n5015 1.505
R27523 net7.n5372 net7.n5370 1.505
R27524 net7.n5378 net7.n5377 1.505
R27525 net7.n5734 net7.n5732 1.505
R27526 net7.n5740 net7.n5739 1.505
R27527 net7.n6096 net7.n6094 1.505
R27528 net7.n6102 net7.n6101 1.505
R27529 net7.n6458 net7.n6456 1.505
R27530 net7.n6464 net7.n6463 1.505
R27531 net7.n6820 net7.n6818 1.505
R27532 net7.n6826 net7.n6825 1.505
R27533 net7.n7182 net7.n7180 1.505
R27534 net7.n7188 net7.n7187 1.505
R27535 net7.n4341 net7.n3979 1.182
R27536 net7 net7.n7237 1.159
R27537 net7.n3369 net7.n3368 1.137
R27538 net7.n3447 net7.n3446 1.137
R27539 net7.n3454 net7.n3453 1.137
R27540 net7.n3458 net7.n3457 1.137
R27541 net7.n3465 net7.n3464 1.137
R27542 net7.n3483 net7.n3482 1.137
R27543 net7.n3500 net7.n3499 1.137
R27544 net7.n3507 net7.n3506 1.137
R27545 net7.n3496 net7.n3495 1.137
R27546 net7.n3489 net7.n3488 1.137
R27547 net7.n3475 net7.n3474 1.137
R27548 net7.n3439 net7.n3438 1.137
R27549 net7.n3430 net7.n3429 1.137
R27550 net7.n3421 net7.n3420 1.137
R27551 net7.n3358 net7.n3357 1.137
R27552 net7.n3365 net7.n3364 1.137
R27553 net7.n3350 net7.n3349 1.137
R27554 net7.n3335 net7.n3334 1.137
R27555 net7.n3319 net7.n3318 1.137
R27556 net7.n3326 net7.n3325 1.137
R27557 net7.n3617 net7.n3616 1.137
R27558 net7.n3007 net7.n3006 1.137
R27559 net7.n3085 net7.n3084 1.137
R27560 net7.n3092 net7.n3091 1.137
R27561 net7.n3096 net7.n3095 1.137
R27562 net7.n3103 net7.n3102 1.137
R27563 net7.n3121 net7.n3120 1.137
R27564 net7.n3138 net7.n3137 1.137
R27565 net7.n3145 net7.n3144 1.137
R27566 net7.n3134 net7.n3133 1.137
R27567 net7.n3127 net7.n3126 1.137
R27568 net7.n3113 net7.n3112 1.137
R27569 net7.n3077 net7.n3076 1.137
R27570 net7.n3068 net7.n3067 1.137
R27571 net7.n3059 net7.n3058 1.137
R27572 net7.n2996 net7.n2995 1.137
R27573 net7.n3003 net7.n3002 1.137
R27574 net7.n2988 net7.n2987 1.137
R27575 net7.n2973 net7.n2972 1.137
R27576 net7.n2957 net7.n2956 1.137
R27577 net7.n2964 net7.n2963 1.137
R27578 net7.n3255 net7.n3254 1.137
R27579 net7.n2645 net7.n2644 1.137
R27580 net7.n2723 net7.n2722 1.137
R27581 net7.n2730 net7.n2729 1.137
R27582 net7.n2734 net7.n2733 1.137
R27583 net7.n2741 net7.n2740 1.137
R27584 net7.n2759 net7.n2758 1.137
R27585 net7.n2776 net7.n2775 1.137
R27586 net7.n2783 net7.n2782 1.137
R27587 net7.n2772 net7.n2771 1.137
R27588 net7.n2765 net7.n2764 1.137
R27589 net7.n2751 net7.n2750 1.137
R27590 net7.n2715 net7.n2714 1.137
R27591 net7.n2706 net7.n2705 1.137
R27592 net7.n2697 net7.n2696 1.137
R27593 net7.n2634 net7.n2633 1.137
R27594 net7.n2641 net7.n2640 1.137
R27595 net7.n2626 net7.n2625 1.137
R27596 net7.n2611 net7.n2610 1.137
R27597 net7.n2595 net7.n2594 1.137
R27598 net7.n2602 net7.n2601 1.137
R27599 net7.n2893 net7.n2892 1.137
R27600 net7.n2283 net7.n2282 1.137
R27601 net7.n2361 net7.n2360 1.137
R27602 net7.n2368 net7.n2367 1.137
R27603 net7.n2372 net7.n2371 1.137
R27604 net7.n2379 net7.n2378 1.137
R27605 net7.n2397 net7.n2396 1.137
R27606 net7.n2414 net7.n2413 1.137
R27607 net7.n2421 net7.n2420 1.137
R27608 net7.n2410 net7.n2409 1.137
R27609 net7.n2403 net7.n2402 1.137
R27610 net7.n2389 net7.n2388 1.137
R27611 net7.n2353 net7.n2352 1.137
R27612 net7.n2344 net7.n2343 1.137
R27613 net7.n2335 net7.n2334 1.137
R27614 net7.n2272 net7.n2271 1.137
R27615 net7.n2279 net7.n2278 1.137
R27616 net7.n2264 net7.n2263 1.137
R27617 net7.n2249 net7.n2248 1.137
R27618 net7.n2233 net7.n2232 1.137
R27619 net7.n2240 net7.n2239 1.137
R27620 net7.n2531 net7.n2530 1.137
R27621 net7.n1921 net7.n1920 1.137
R27622 net7.n1999 net7.n1998 1.137
R27623 net7.n2006 net7.n2005 1.137
R27624 net7.n2010 net7.n2009 1.137
R27625 net7.n2017 net7.n2016 1.137
R27626 net7.n2035 net7.n2034 1.137
R27627 net7.n2052 net7.n2051 1.137
R27628 net7.n2059 net7.n2058 1.137
R27629 net7.n2048 net7.n2047 1.137
R27630 net7.n2041 net7.n2040 1.137
R27631 net7.n2027 net7.n2026 1.137
R27632 net7.n1991 net7.n1990 1.137
R27633 net7.n1982 net7.n1981 1.137
R27634 net7.n1973 net7.n1972 1.137
R27635 net7.n1910 net7.n1909 1.137
R27636 net7.n1917 net7.n1916 1.137
R27637 net7.n1902 net7.n1901 1.137
R27638 net7.n1887 net7.n1886 1.137
R27639 net7.n1871 net7.n1870 1.137
R27640 net7.n1878 net7.n1877 1.137
R27641 net7.n2169 net7.n2168 1.137
R27642 net7.n1559 net7.n1558 1.137
R27643 net7.n1637 net7.n1636 1.137
R27644 net7.n1644 net7.n1643 1.137
R27645 net7.n1648 net7.n1647 1.137
R27646 net7.n1655 net7.n1654 1.137
R27647 net7.n1673 net7.n1672 1.137
R27648 net7.n1690 net7.n1689 1.137
R27649 net7.n1697 net7.n1696 1.137
R27650 net7.n1686 net7.n1685 1.137
R27651 net7.n1679 net7.n1678 1.137
R27652 net7.n1665 net7.n1664 1.137
R27653 net7.n1629 net7.n1628 1.137
R27654 net7.n1620 net7.n1619 1.137
R27655 net7.n1611 net7.n1610 1.137
R27656 net7.n1548 net7.n1547 1.137
R27657 net7.n1555 net7.n1554 1.137
R27658 net7.n1540 net7.n1539 1.137
R27659 net7.n1525 net7.n1524 1.137
R27660 net7.n1509 net7.n1508 1.137
R27661 net7.n1516 net7.n1515 1.137
R27662 net7.n1807 net7.n1806 1.137
R27663 net7.n1197 net7.n1196 1.137
R27664 net7.n1275 net7.n1274 1.137
R27665 net7.n1282 net7.n1281 1.137
R27666 net7.n1286 net7.n1285 1.137
R27667 net7.n1293 net7.n1292 1.137
R27668 net7.n1311 net7.n1310 1.137
R27669 net7.n1328 net7.n1327 1.137
R27670 net7.n1335 net7.n1334 1.137
R27671 net7.n1324 net7.n1323 1.137
R27672 net7.n1317 net7.n1316 1.137
R27673 net7.n1303 net7.n1302 1.137
R27674 net7.n1267 net7.n1266 1.137
R27675 net7.n1258 net7.n1257 1.137
R27676 net7.n1249 net7.n1248 1.137
R27677 net7.n1186 net7.n1185 1.137
R27678 net7.n1193 net7.n1192 1.137
R27679 net7.n1178 net7.n1177 1.137
R27680 net7.n1163 net7.n1162 1.137
R27681 net7.n1147 net7.n1146 1.137
R27682 net7.n1154 net7.n1153 1.137
R27683 net7.n1445 net7.n1444 1.137
R27684 net7.n835 net7.n834 1.137
R27685 net7.n913 net7.n912 1.137
R27686 net7.n920 net7.n919 1.137
R27687 net7.n924 net7.n923 1.137
R27688 net7.n931 net7.n930 1.137
R27689 net7.n949 net7.n948 1.137
R27690 net7.n966 net7.n965 1.137
R27691 net7.n973 net7.n972 1.137
R27692 net7.n962 net7.n961 1.137
R27693 net7.n955 net7.n954 1.137
R27694 net7.n941 net7.n940 1.137
R27695 net7.n905 net7.n904 1.137
R27696 net7.n896 net7.n895 1.137
R27697 net7.n887 net7.n886 1.137
R27698 net7.n824 net7.n823 1.137
R27699 net7.n831 net7.n830 1.137
R27700 net7.n816 net7.n815 1.137
R27701 net7.n801 net7.n800 1.137
R27702 net7.n785 net7.n784 1.137
R27703 net7.n792 net7.n791 1.137
R27704 net7.n1083 net7.n1082 1.137
R27705 net7.n473 net7.n472 1.137
R27706 net7.n551 net7.n550 1.137
R27707 net7.n558 net7.n557 1.137
R27708 net7.n562 net7.n561 1.137
R27709 net7.n569 net7.n568 1.137
R27710 net7.n587 net7.n586 1.137
R27711 net7.n604 net7.n603 1.137
R27712 net7.n611 net7.n610 1.137
R27713 net7.n600 net7.n599 1.137
R27714 net7.n593 net7.n592 1.137
R27715 net7.n579 net7.n578 1.137
R27716 net7.n543 net7.n542 1.137
R27717 net7.n534 net7.n533 1.137
R27718 net7.n525 net7.n524 1.137
R27719 net7.n462 net7.n461 1.137
R27720 net7.n469 net7.n468 1.137
R27721 net7.n454 net7.n453 1.137
R27722 net7.n439 net7.n438 1.137
R27723 net7.n423 net7.n422 1.137
R27724 net7.n430 net7.n429 1.137
R27725 net7.n721 net7.n720 1.137
R27726 net7.n360 net7.n359 1.137
R27727 net7.n112 net7.n111 1.137
R27728 net7.n190 net7.n189 1.137
R27729 net7.n197 net7.n196 1.137
R27730 net7.n201 net7.n200 1.137
R27731 net7.n208 net7.n207 1.137
R27732 net7.n226 net7.n225 1.137
R27733 net7.n243 net7.n242 1.137
R27734 net7.n239 net7.n238 1.137
R27735 net7.n232 net7.n231 1.137
R27736 net7.n218 net7.n217 1.137
R27737 net7.n182 net7.n181 1.137
R27738 net7.n173 net7.n172 1.137
R27739 net7.n164 net7.n163 1.137
R27740 net7.n101 net7.n100 1.137
R27741 net7.n108 net7.n107 1.137
R27742 net7.n93 net7.n92 1.137
R27743 net7.n78 net7.n77 1.137
R27744 net7.n62 net7.n61 1.137
R27745 net7.n69 net7.n68 1.137
R27746 net7.n250 net7.n249 1.137
R27747 net7.n3894 net7.n3893 1.137
R27748 net7.n3902 net7.n3901 1.137
R27749 net7.n3852 net7.n3851 1.137
R27750 net7.n3745 net7.n3744 1.137
R27751 net7.n3717 net7.n3716 1.137
R27752 net7.n3703 net7.n3702 1.137
R27753 net7.n3709 net7.n3708 1.137
R27754 net7.n3726 net7.n3725 1.137
R27755 net7.n3741 net7.n3740 1.137
R27756 net7.n3734 net7.n3733 1.137
R27757 net7.n3752 net7.n3751 1.137
R27758 net7.n3762 net7.n3761 1.137
R27759 net7.n3848 net7.n3847 1.137
R27760 net7.n3771 net7.n3770 1.137
R27761 net7.n3841 net7.n3840 1.137
R27762 net7.n3859 net7.n3858 1.137
R27763 net7.n3869 net7.n3868 1.137
R27764 net7.n3875 net7.n3874 1.137
R27765 net7.n3890 net7.n3889 1.137
R27766 net7.n3883 net7.n3882 1.137
R27767 net7.n3979 net7.n3978 1.137
R27768 net7.n4255 net7.n4254 1.137
R27769 net7.n4263 net7.n4262 1.137
R27770 net7.n4213 net7.n4212 1.137
R27771 net7.n4106 net7.n4105 1.137
R27772 net7.n4078 net7.n4077 1.137
R27773 net7.n4064 net7.n4063 1.137
R27774 net7.n4070 net7.n4069 1.137
R27775 net7.n4087 net7.n4086 1.137
R27776 net7.n4102 net7.n4101 1.137
R27777 net7.n4095 net7.n4094 1.137
R27778 net7.n4113 net7.n4112 1.137
R27779 net7.n4123 net7.n4122 1.137
R27780 net7.n4209 net7.n4208 1.137
R27781 net7.n4132 net7.n4131 1.137
R27782 net7.n4202 net7.n4201 1.137
R27783 net7.n4220 net7.n4219 1.137
R27784 net7.n4230 net7.n4229 1.137
R27785 net7.n4236 net7.n4235 1.137
R27786 net7.n4251 net7.n4250 1.137
R27787 net7.n4244 net7.n4243 1.137
R27788 net7.n4340 net7.n4339 1.137
R27789 net7.n4617 net7.n4616 1.137
R27790 net7.n4625 net7.n4624 1.137
R27791 net7.n4575 net7.n4574 1.137
R27792 net7.n4468 net7.n4467 1.137
R27793 net7.n4440 net7.n4439 1.137
R27794 net7.n4426 net7.n4425 1.137
R27795 net7.n4432 net7.n4431 1.137
R27796 net7.n4449 net7.n4448 1.137
R27797 net7.n4464 net7.n4463 1.137
R27798 net7.n4457 net7.n4456 1.137
R27799 net7.n4475 net7.n4474 1.137
R27800 net7.n4485 net7.n4484 1.137
R27801 net7.n4571 net7.n4570 1.137
R27802 net7.n4494 net7.n4493 1.137
R27803 net7.n4564 net7.n4563 1.137
R27804 net7.n4582 net7.n4581 1.137
R27805 net7.n4592 net7.n4591 1.137
R27806 net7.n4598 net7.n4597 1.137
R27807 net7.n4613 net7.n4612 1.137
R27808 net7.n4606 net7.n4605 1.137
R27809 net7.n4702 net7.n4701 1.137
R27810 net7.n4979 net7.n4978 1.137
R27811 net7.n4987 net7.n4986 1.137
R27812 net7.n4937 net7.n4936 1.137
R27813 net7.n4830 net7.n4829 1.137
R27814 net7.n4802 net7.n4801 1.137
R27815 net7.n4788 net7.n4787 1.137
R27816 net7.n4794 net7.n4793 1.137
R27817 net7.n4811 net7.n4810 1.137
R27818 net7.n4826 net7.n4825 1.137
R27819 net7.n4819 net7.n4818 1.137
R27820 net7.n4837 net7.n4836 1.137
R27821 net7.n4847 net7.n4846 1.137
R27822 net7.n4933 net7.n4932 1.137
R27823 net7.n4856 net7.n4855 1.137
R27824 net7.n4926 net7.n4925 1.137
R27825 net7.n4944 net7.n4943 1.137
R27826 net7.n4954 net7.n4953 1.137
R27827 net7.n4960 net7.n4959 1.137
R27828 net7.n4975 net7.n4974 1.137
R27829 net7.n4968 net7.n4967 1.137
R27830 net7.n5064 net7.n5063 1.137
R27831 net7.n5341 net7.n5340 1.137
R27832 net7.n5349 net7.n5348 1.137
R27833 net7.n5299 net7.n5298 1.137
R27834 net7.n5192 net7.n5191 1.137
R27835 net7.n5164 net7.n5163 1.137
R27836 net7.n5150 net7.n5149 1.137
R27837 net7.n5156 net7.n5155 1.137
R27838 net7.n5173 net7.n5172 1.137
R27839 net7.n5188 net7.n5187 1.137
R27840 net7.n5181 net7.n5180 1.137
R27841 net7.n5199 net7.n5198 1.137
R27842 net7.n5209 net7.n5208 1.137
R27843 net7.n5295 net7.n5294 1.137
R27844 net7.n5218 net7.n5217 1.137
R27845 net7.n5288 net7.n5287 1.137
R27846 net7.n5306 net7.n5305 1.137
R27847 net7.n5316 net7.n5315 1.137
R27848 net7.n5322 net7.n5321 1.137
R27849 net7.n5337 net7.n5336 1.137
R27850 net7.n5330 net7.n5329 1.137
R27851 net7.n5426 net7.n5425 1.137
R27852 net7.n5703 net7.n5702 1.137
R27853 net7.n5711 net7.n5710 1.137
R27854 net7.n5661 net7.n5660 1.137
R27855 net7.n5554 net7.n5553 1.137
R27856 net7.n5526 net7.n5525 1.137
R27857 net7.n5512 net7.n5511 1.137
R27858 net7.n5518 net7.n5517 1.137
R27859 net7.n5535 net7.n5534 1.137
R27860 net7.n5550 net7.n5549 1.137
R27861 net7.n5543 net7.n5542 1.137
R27862 net7.n5561 net7.n5560 1.137
R27863 net7.n5571 net7.n5570 1.137
R27864 net7.n5657 net7.n5656 1.137
R27865 net7.n5580 net7.n5579 1.137
R27866 net7.n5650 net7.n5649 1.137
R27867 net7.n5668 net7.n5667 1.137
R27868 net7.n5678 net7.n5677 1.137
R27869 net7.n5684 net7.n5683 1.137
R27870 net7.n5699 net7.n5698 1.137
R27871 net7.n5692 net7.n5691 1.137
R27872 net7.n5788 net7.n5787 1.137
R27873 net7.n6065 net7.n6064 1.137
R27874 net7.n6073 net7.n6072 1.137
R27875 net7.n6023 net7.n6022 1.137
R27876 net7.n5916 net7.n5915 1.137
R27877 net7.n5888 net7.n5887 1.137
R27878 net7.n5874 net7.n5873 1.137
R27879 net7.n5880 net7.n5879 1.137
R27880 net7.n5897 net7.n5896 1.137
R27881 net7.n5912 net7.n5911 1.137
R27882 net7.n5905 net7.n5904 1.137
R27883 net7.n5923 net7.n5922 1.137
R27884 net7.n5933 net7.n5932 1.137
R27885 net7.n6019 net7.n6018 1.137
R27886 net7.n5942 net7.n5941 1.137
R27887 net7.n6012 net7.n6011 1.137
R27888 net7.n6030 net7.n6029 1.137
R27889 net7.n6040 net7.n6039 1.137
R27890 net7.n6046 net7.n6045 1.137
R27891 net7.n6061 net7.n6060 1.137
R27892 net7.n6054 net7.n6053 1.137
R27893 net7.n6150 net7.n6149 1.137
R27894 net7.n6427 net7.n6426 1.137
R27895 net7.n6435 net7.n6434 1.137
R27896 net7.n6385 net7.n6384 1.137
R27897 net7.n6278 net7.n6277 1.137
R27898 net7.n6250 net7.n6249 1.137
R27899 net7.n6236 net7.n6235 1.137
R27900 net7.n6242 net7.n6241 1.137
R27901 net7.n6259 net7.n6258 1.137
R27902 net7.n6274 net7.n6273 1.137
R27903 net7.n6267 net7.n6266 1.137
R27904 net7.n6285 net7.n6284 1.137
R27905 net7.n6295 net7.n6294 1.137
R27906 net7.n6381 net7.n6380 1.137
R27907 net7.n6304 net7.n6303 1.137
R27908 net7.n6374 net7.n6373 1.137
R27909 net7.n6392 net7.n6391 1.137
R27910 net7.n6402 net7.n6401 1.137
R27911 net7.n6408 net7.n6407 1.137
R27912 net7.n6423 net7.n6422 1.137
R27913 net7.n6416 net7.n6415 1.137
R27914 net7.n6512 net7.n6511 1.137
R27915 net7.n6789 net7.n6788 1.137
R27916 net7.n6797 net7.n6796 1.137
R27917 net7.n6747 net7.n6746 1.137
R27918 net7.n6640 net7.n6639 1.137
R27919 net7.n6612 net7.n6611 1.137
R27920 net7.n6598 net7.n6597 1.137
R27921 net7.n6604 net7.n6603 1.137
R27922 net7.n6621 net7.n6620 1.137
R27923 net7.n6636 net7.n6635 1.137
R27924 net7.n6629 net7.n6628 1.137
R27925 net7.n6647 net7.n6646 1.137
R27926 net7.n6657 net7.n6656 1.137
R27927 net7.n6743 net7.n6742 1.137
R27928 net7.n6666 net7.n6665 1.137
R27929 net7.n6736 net7.n6735 1.137
R27930 net7.n6754 net7.n6753 1.137
R27931 net7.n6764 net7.n6763 1.137
R27932 net7.n6770 net7.n6769 1.137
R27933 net7.n6785 net7.n6784 1.137
R27934 net7.n6778 net7.n6777 1.137
R27935 net7.n6874 net7.n6873 1.137
R27936 net7.n7151 net7.n7150 1.137
R27937 net7.n7159 net7.n7158 1.137
R27938 net7.n7109 net7.n7108 1.137
R27939 net7.n7002 net7.n7001 1.137
R27940 net7.n6974 net7.n6973 1.137
R27941 net7.n6960 net7.n6959 1.137
R27942 net7.n6966 net7.n6965 1.137
R27943 net7.n6983 net7.n6982 1.137
R27944 net7.n6998 net7.n6997 1.137
R27945 net7.n6991 net7.n6990 1.137
R27946 net7.n7009 net7.n7008 1.137
R27947 net7.n7019 net7.n7018 1.137
R27948 net7.n7105 net7.n7104 1.137
R27949 net7.n7028 net7.n7027 1.137
R27950 net7.n7098 net7.n7097 1.137
R27951 net7.n7116 net7.n7115 1.137
R27952 net7.n7126 net7.n7125 1.137
R27953 net7.n7132 net7.n7131 1.137
R27954 net7.n7147 net7.n7146 1.137
R27955 net7.n7140 net7.n7139 1.137
R27956 net7.n7236 net7.n7235 1.137
R27957 net7.n3512 net7.n3511 1.129
R27958 net7.n3519 net7.n3518 1.129
R27959 net7.n3557 net7.n3556 1.129
R27960 net7.n3150 net7.n3149 1.129
R27961 net7.n3157 net7.n3156 1.129
R27962 net7.n3195 net7.n3194 1.129
R27963 net7.n2788 net7.n2787 1.129
R27964 net7.n2795 net7.n2794 1.129
R27965 net7.n2833 net7.n2832 1.129
R27966 net7.n2426 net7.n2425 1.129
R27967 net7.n2433 net7.n2432 1.129
R27968 net7.n2471 net7.n2470 1.129
R27969 net7.n2064 net7.n2063 1.129
R27970 net7.n2071 net7.n2070 1.129
R27971 net7.n2109 net7.n2108 1.129
R27972 net7.n1702 net7.n1701 1.129
R27973 net7.n1709 net7.n1708 1.129
R27974 net7.n1747 net7.n1746 1.129
R27975 net7.n1340 net7.n1339 1.129
R27976 net7.n1347 net7.n1346 1.129
R27977 net7.n1385 net7.n1384 1.129
R27978 net7.n978 net7.n977 1.129
R27979 net7.n985 net7.n984 1.129
R27980 net7.n1023 net7.n1022 1.129
R27981 net7.n616 net7.n615 1.129
R27982 net7.n623 net7.n622 1.129
R27983 net7.n661 net7.n660 1.129
R27984 net7.n255 net7.n254 1.129
R27985 net7.n262 net7.n261 1.129
R27986 net7.n300 net7.n299 1.129
R27987 net7.n3633 net7.n3632 1.129
R27988 net7.n3646 net7.n3645 1.129
R27989 net7.n3649 net7.n3648 1.129
R27990 net7.n3994 net7.n3993 1.129
R27991 net7.n4007 net7.n4006 1.129
R27992 net7.n4010 net7.n4009 1.129
R27993 net7.n4356 net7.n4355 1.129
R27994 net7.n4369 net7.n4368 1.129
R27995 net7.n4372 net7.n4371 1.129
R27996 net7.n4718 net7.n4717 1.129
R27997 net7.n4731 net7.n4730 1.129
R27998 net7.n4734 net7.n4733 1.129
R27999 net7.n5080 net7.n5079 1.129
R28000 net7.n5093 net7.n5092 1.129
R28001 net7.n5096 net7.n5095 1.129
R28002 net7.n5442 net7.n5441 1.129
R28003 net7.n5455 net7.n5454 1.129
R28004 net7.n5458 net7.n5457 1.129
R28005 net7.n5804 net7.n5803 1.129
R28006 net7.n5817 net7.n5816 1.129
R28007 net7.n5820 net7.n5819 1.129
R28008 net7.n6166 net7.n6165 1.129
R28009 net7.n6179 net7.n6178 1.129
R28010 net7.n6182 net7.n6181 1.129
R28011 net7.n6528 net7.n6527 1.129
R28012 net7.n6541 net7.n6540 1.129
R28013 net7.n6544 net7.n6543 1.129
R28014 net7.n6890 net7.n6889 1.129
R28015 net7.n6903 net7.n6902 1.129
R28016 net7.n6906 net7.n6905 1.129
R28017 net7.n3347 net7.n3346 1.125
R28018 net7.n2985 net7.n2984 1.125
R28019 net7.n2623 net7.n2622 1.125
R28020 net7.n2261 net7.n2260 1.125
R28021 net7.n1899 net7.n1898 1.125
R28022 net7.n1537 net7.n1536 1.125
R28023 net7.n1175 net7.n1174 1.125
R28024 net7.n813 net7.n812 1.125
R28025 net7.n451 net7.n450 1.125
R28026 net7.n90 net7.n89 1.125
R28027 net7.n4341 net7.n4340 1.089
R28028 net7.n4703 net7.n4702 1.089
R28029 net7.n5065 net7.n5064 1.089
R28030 net7.n5427 net7.n5426 1.089
R28031 net7.n5789 net7.n5788 1.089
R28032 net7.n6151 net7.n6150 1.089
R28033 net7.n6513 net7.n6512 1.089
R28034 net7.n6875 net7.n6874 1.089
R28035 net7.n7237 net7.n7236 1.089
R28036 net7.n3420 net7.n3417 1.042
R28037 net7.n3058 net7.n3055 1.042
R28038 net7.n2696 net7.n2693 1.042
R28039 net7.n2334 net7.n2331 1.042
R28040 net7.n1972 net7.n1969 1.042
R28041 net7.n1610 net7.n1607 1.042
R28042 net7.n1248 net7.n1245 1.042
R28043 net7.n886 net7.n883 1.042
R28044 net7.n524 net7.n521 1.042
R28045 net7.n163 net7.n160 1.042
R28046 net7.n3840 net7.n3839 1.042
R28047 net7.n4201 net7.n4200 1.042
R28048 net7.n4563 net7.n4562 1.042
R28049 net7.n4925 net7.n4924 1.042
R28050 net7.n5287 net7.n5286 1.042
R28051 net7.n5649 net7.n5648 1.042
R28052 net7.n6011 net7.n6010 1.042
R28053 net7.n6373 net7.n6372 1.042
R28054 net7.n6735 net7.n6734 1.042
R28055 net7.n7097 net7.n7096 1.042
R28056 net7.n3311 net7.n3310 0.869
R28057 net7.n2949 net7.n2948 0.869
R28058 net7.n2587 net7.n2586 0.869
R28059 net7.n2225 net7.n2224 0.869
R28060 net7.n1863 net7.n1862 0.869
R28061 net7.n1501 net7.n1500 0.869
R28062 net7.n1139 net7.n1138 0.869
R28063 net7.n777 net7.n776 0.869
R28064 net7.n415 net7.n414 0.869
R28065 net7.n54 net7.n53 0.869
R28066 net7.n3695 net7.n3694 0.869
R28067 net7.n4056 net7.n4055 0.869
R28068 net7.n4418 net7.n4417 0.869
R28069 net7.n4780 net7.n4779 0.869
R28070 net7.n5142 net7.n5141 0.869
R28071 net7.n5504 net7.n5503 0.869
R28072 net7.n5866 net7.n5865 0.869
R28073 net7.n6228 net7.n6227 0.869
R28074 net7.n6590 net7.n6589 0.869
R28075 net7.n6952 net7.n6951 0.869
R28076 net7.n3602 net7.n3601 0.752
R28077 net7.n3416 net7.n3415 0.752
R28078 net7.n3389 net7.n3388 0.752
R28079 net7.n3272 net7.n3270 0.752
R28080 net7.n3291 net7.n3290 0.752
R28081 net7.n3302 net7.n3301 0.752
R28082 net7.n3240 net7.n3239 0.752
R28083 net7.n3054 net7.n3053 0.752
R28084 net7.n3027 net7.n3026 0.752
R28085 net7.n2910 net7.n2908 0.752
R28086 net7.n2929 net7.n2928 0.752
R28087 net7.n2940 net7.n2939 0.752
R28088 net7.n2878 net7.n2877 0.752
R28089 net7.n2692 net7.n2691 0.752
R28090 net7.n2665 net7.n2664 0.752
R28091 net7.n2548 net7.n2546 0.752
R28092 net7.n2567 net7.n2566 0.752
R28093 net7.n2578 net7.n2577 0.752
R28094 net7.n2516 net7.n2515 0.752
R28095 net7.n2330 net7.n2329 0.752
R28096 net7.n2303 net7.n2302 0.752
R28097 net7.n2186 net7.n2184 0.752
R28098 net7.n2205 net7.n2204 0.752
R28099 net7.n2216 net7.n2215 0.752
R28100 net7.n2154 net7.n2153 0.752
R28101 net7.n1968 net7.n1967 0.752
R28102 net7.n1941 net7.n1940 0.752
R28103 net7.n1824 net7.n1822 0.752
R28104 net7.n1843 net7.n1842 0.752
R28105 net7.n1854 net7.n1853 0.752
R28106 net7.n1792 net7.n1791 0.752
R28107 net7.n1606 net7.n1605 0.752
R28108 net7.n1579 net7.n1578 0.752
R28109 net7.n1462 net7.n1460 0.752
R28110 net7.n1481 net7.n1480 0.752
R28111 net7.n1492 net7.n1491 0.752
R28112 net7.n1430 net7.n1429 0.752
R28113 net7.n1244 net7.n1243 0.752
R28114 net7.n1217 net7.n1216 0.752
R28115 net7.n1100 net7.n1098 0.752
R28116 net7.n1119 net7.n1118 0.752
R28117 net7.n1130 net7.n1129 0.752
R28118 net7.n1068 net7.n1067 0.752
R28119 net7.n882 net7.n881 0.752
R28120 net7.n855 net7.n854 0.752
R28121 net7.n738 net7.n736 0.752
R28122 net7.n757 net7.n756 0.752
R28123 net7.n768 net7.n767 0.752
R28124 net7.n706 net7.n705 0.752
R28125 net7.n520 net7.n519 0.752
R28126 net7.n493 net7.n492 0.752
R28127 net7.n376 net7.n374 0.752
R28128 net7.n395 net7.n394 0.752
R28129 net7.n406 net7.n405 0.752
R28130 net7.n345 net7.n344 0.752
R28131 net7.n159 net7.n158 0.752
R28132 net7.n132 net7.n131 0.752
R28133 net7.n15 net7.n13 0.752
R28134 net7.n34 net7.n33 0.752
R28135 net7.n45 net7.n44 0.752
R28136 net7.n3630 net7.n3629 0.752
R28137 net7.n3827 net7.n3826 0.752
R28138 net7.n3917 net7.n3916 0.752
R28139 net7.n3939 net7.n3937 0.752
R28140 net7.n3958 net7.n3957 0.752
R28141 net7.n3969 net7.n3968 0.752
R28142 net7.n3991 net7.n3990 0.752
R28143 net7.n4188 net7.n4187 0.752
R28144 net7.n4278 net7.n4277 0.752
R28145 net7.n4300 net7.n4298 0.752
R28146 net7.n4319 net7.n4318 0.752
R28147 net7.n4330 net7.n4329 0.752
R28148 net7.n4353 net7.n4352 0.752
R28149 net7.n4550 net7.n4549 0.752
R28150 net7.n4640 net7.n4639 0.752
R28151 net7.n4662 net7.n4660 0.752
R28152 net7.n4681 net7.n4680 0.752
R28153 net7.n4692 net7.n4691 0.752
R28154 net7.n4715 net7.n4714 0.752
R28155 net7.n4912 net7.n4911 0.752
R28156 net7.n5002 net7.n5001 0.752
R28157 net7.n5024 net7.n5022 0.752
R28158 net7.n5043 net7.n5042 0.752
R28159 net7.n5054 net7.n5053 0.752
R28160 net7.n5077 net7.n5076 0.752
R28161 net7.n5274 net7.n5273 0.752
R28162 net7.n5364 net7.n5363 0.752
R28163 net7.n5386 net7.n5384 0.752
R28164 net7.n5405 net7.n5404 0.752
R28165 net7.n5416 net7.n5415 0.752
R28166 net7.n5439 net7.n5438 0.752
R28167 net7.n5636 net7.n5635 0.752
R28168 net7.n5726 net7.n5725 0.752
R28169 net7.n5748 net7.n5746 0.752
R28170 net7.n5767 net7.n5766 0.752
R28171 net7.n5778 net7.n5777 0.752
R28172 net7.n5801 net7.n5800 0.752
R28173 net7.n5998 net7.n5997 0.752
R28174 net7.n6088 net7.n6087 0.752
R28175 net7.n6110 net7.n6108 0.752
R28176 net7.n6129 net7.n6128 0.752
R28177 net7.n6140 net7.n6139 0.752
R28178 net7.n6163 net7.n6162 0.752
R28179 net7.n6360 net7.n6359 0.752
R28180 net7.n6450 net7.n6449 0.752
R28181 net7.n6472 net7.n6470 0.752
R28182 net7.n6491 net7.n6490 0.752
R28183 net7.n6502 net7.n6501 0.752
R28184 net7.n6525 net7.n6524 0.752
R28185 net7.n6722 net7.n6721 0.752
R28186 net7.n6812 net7.n6811 0.752
R28187 net7.n6834 net7.n6832 0.752
R28188 net7.n6853 net7.n6852 0.752
R28189 net7.n6864 net7.n6863 0.752
R28190 net7.n6887 net7.n6886 0.752
R28191 net7.n7084 net7.n7083 0.752
R28192 net7.n7174 net7.n7173 0.752
R28193 net7.n7196 net7.n7194 0.752
R28194 net7.n7215 net7.n7214 0.752
R28195 net7.n7226 net7.n7225 0.752
R28196 net7 net7.n3618 0.743
R28197 net7.n3694 net7.n3693 0.729
R28198 net7.n4055 net7.n4054 0.729
R28199 net7.n4417 net7.n4416 0.729
R28200 net7.n4779 net7.n4778 0.729
R28201 net7.n5141 net7.n5140 0.729
R28202 net7.n5503 net7.n5502 0.729
R28203 net7.n5865 net7.n5864 0.729
R28204 net7.n6227 net7.n6226 0.729
R28205 net7.n6589 net7.n6588 0.729
R28206 net7.n6951 net7.n6950 0.729
R28207 net7.n3310 net7.n3309 0.728
R28208 net7.n2948 net7.n2947 0.728
R28209 net7.n2586 net7.n2585 0.728
R28210 net7.n2224 net7.n2223 0.728
R28211 net7.n1862 net7.n1861 0.728
R28212 net7.n1500 net7.n1499 0.728
R28213 net7.n1138 net7.n1137 0.728
R28214 net7.n776 net7.n775 0.728
R28215 net7.n414 net7.n413 0.728
R28216 net7.n53 net7.n52 0.728
R28217 net7.n3978 net7.n3977 0.725
R28218 net7.n4339 net7.n4338 0.725
R28219 net7.n4701 net7.n4700 0.725
R28220 net7.n5063 net7.n5062 0.725
R28221 net7.n5425 net7.n5424 0.725
R28222 net7.n5787 net7.n5786 0.725
R28223 net7.n6149 net7.n6148 0.725
R28224 net7.n6511 net7.n6510 0.725
R28225 net7.n6873 net7.n6872 0.725
R28226 net7.n7235 net7.n7234 0.725
R28227 net7.n3616 net7.n3610 0.725
R28228 net7.n3254 net7.n3248 0.725
R28229 net7.n2892 net7.n2886 0.725
R28230 net7.n2530 net7.n2524 0.725
R28231 net7.n2168 net7.n2162 0.725
R28232 net7.n1806 net7.n1800 0.725
R28233 net7.n1444 net7.n1438 0.725
R28234 net7.n1082 net7.n1076 0.725
R28235 net7.n720 net7.n714 0.725
R28236 net7.n359 net7.n353 0.725
R28237 net7.n3583 net7.n3582 0.376
R28238 net7.n3515 net7.n3514 0.376
R28239 net7.n3521 net7.n3520 0.376
R28240 net7.n3534 net7.n3533 0.376
R28241 net7.n3523 net7.n3522 0.376
R28242 net7.n3379 net7.n3378 0.376
R28243 net7.n3221 net7.n3220 0.376
R28244 net7.n3153 net7.n3152 0.376
R28245 net7.n3159 net7.n3158 0.376
R28246 net7.n3172 net7.n3171 0.376
R28247 net7.n3161 net7.n3160 0.376
R28248 net7.n3017 net7.n3016 0.376
R28249 net7.n2859 net7.n2858 0.376
R28250 net7.n2791 net7.n2790 0.376
R28251 net7.n2797 net7.n2796 0.376
R28252 net7.n2810 net7.n2809 0.376
R28253 net7.n2799 net7.n2798 0.376
R28254 net7.n2655 net7.n2654 0.376
R28255 net7.n2497 net7.n2496 0.376
R28256 net7.n2429 net7.n2428 0.376
R28257 net7.n2435 net7.n2434 0.376
R28258 net7.n2448 net7.n2447 0.376
R28259 net7.n2437 net7.n2436 0.376
R28260 net7.n2293 net7.n2292 0.376
R28261 net7.n2135 net7.n2134 0.376
R28262 net7.n2067 net7.n2066 0.376
R28263 net7.n2073 net7.n2072 0.376
R28264 net7.n2086 net7.n2085 0.376
R28265 net7.n2075 net7.n2074 0.376
R28266 net7.n1931 net7.n1930 0.376
R28267 net7.n1773 net7.n1772 0.376
R28268 net7.n1705 net7.n1704 0.376
R28269 net7.n1711 net7.n1710 0.376
R28270 net7.n1724 net7.n1723 0.376
R28271 net7.n1713 net7.n1712 0.376
R28272 net7.n1569 net7.n1568 0.376
R28273 net7.n1411 net7.n1410 0.376
R28274 net7.n1343 net7.n1342 0.376
R28275 net7.n1349 net7.n1348 0.376
R28276 net7.n1362 net7.n1361 0.376
R28277 net7.n1351 net7.n1350 0.376
R28278 net7.n1207 net7.n1206 0.376
R28279 net7.n1049 net7.n1048 0.376
R28280 net7.n981 net7.n980 0.376
R28281 net7.n987 net7.n986 0.376
R28282 net7.n1000 net7.n999 0.376
R28283 net7.n989 net7.n988 0.376
R28284 net7.n845 net7.n844 0.376
R28285 net7.n687 net7.n686 0.376
R28286 net7.n619 net7.n618 0.376
R28287 net7.n625 net7.n624 0.376
R28288 net7.n638 net7.n637 0.376
R28289 net7.n627 net7.n626 0.376
R28290 net7.n483 net7.n482 0.376
R28291 net7.n326 net7.n325 0.376
R28292 net7.n258 net7.n257 0.376
R28293 net7.n264 net7.n263 0.376
R28294 net7.n277 net7.n276 0.376
R28295 net7.n266 net7.n265 0.376
R28296 net7.n122 net7.n121 0.376
R28297 net7.n3636 net7.n3635 0.376
R28298 net7.n3639 net7.n3638 0.376
R28299 net7.n3786 net7.n3785 0.376
R28300 net7.n3798 net7.n3797 0.376
R28301 net7.n3808 net7.n3807 0.376
R28302 net7.n3818 net7.n3817 0.376
R28303 net7.n3997 net7.n3996 0.376
R28304 net7.n4000 net7.n3999 0.376
R28305 net7.n4147 net7.n4146 0.376
R28306 net7.n4159 net7.n4158 0.376
R28307 net7.n4169 net7.n4168 0.376
R28308 net7.n4179 net7.n4178 0.376
R28309 net7.n4359 net7.n4358 0.376
R28310 net7.n4362 net7.n4361 0.376
R28311 net7.n4509 net7.n4508 0.376
R28312 net7.n4521 net7.n4520 0.376
R28313 net7.n4531 net7.n4530 0.376
R28314 net7.n4541 net7.n4540 0.376
R28315 net7.n4721 net7.n4720 0.376
R28316 net7.n4724 net7.n4723 0.376
R28317 net7.n4871 net7.n4870 0.376
R28318 net7.n4883 net7.n4882 0.376
R28319 net7.n4893 net7.n4892 0.376
R28320 net7.n4903 net7.n4902 0.376
R28321 net7.n5083 net7.n5082 0.376
R28322 net7.n5086 net7.n5085 0.376
R28323 net7.n5233 net7.n5232 0.376
R28324 net7.n5245 net7.n5244 0.376
R28325 net7.n5255 net7.n5254 0.376
R28326 net7.n5265 net7.n5264 0.376
R28327 net7.n5445 net7.n5444 0.376
R28328 net7.n5448 net7.n5447 0.376
R28329 net7.n5595 net7.n5594 0.376
R28330 net7.n5607 net7.n5606 0.376
R28331 net7.n5617 net7.n5616 0.376
R28332 net7.n5627 net7.n5626 0.376
R28333 net7.n5807 net7.n5806 0.376
R28334 net7.n5810 net7.n5809 0.376
R28335 net7.n5957 net7.n5956 0.376
R28336 net7.n5969 net7.n5968 0.376
R28337 net7.n5979 net7.n5978 0.376
R28338 net7.n5989 net7.n5988 0.376
R28339 net7.n6169 net7.n6168 0.376
R28340 net7.n6172 net7.n6171 0.376
R28341 net7.n6319 net7.n6318 0.376
R28342 net7.n6331 net7.n6330 0.376
R28343 net7.n6341 net7.n6340 0.376
R28344 net7.n6351 net7.n6350 0.376
R28345 net7.n6531 net7.n6530 0.376
R28346 net7.n6534 net7.n6533 0.376
R28347 net7.n6681 net7.n6680 0.376
R28348 net7.n6693 net7.n6692 0.376
R28349 net7.n6703 net7.n6702 0.376
R28350 net7.n6713 net7.n6712 0.376
R28351 net7.n6893 net7.n6892 0.376
R28352 net7.n6896 net7.n6895 0.376
R28353 net7.n7043 net7.n7042 0.376
R28354 net7.n7055 net7.n7054 0.376
R28355 net7.n7065 net7.n7064 0.376
R28356 net7.n7075 net7.n7074 0.376
R28357 net7.n3382 net7.n3381 0.189
R28358 net7.n3020 net7.n3019 0.189
R28359 net7.n2658 net7.n2657 0.189
R28360 net7.n2296 net7.n2295 0.189
R28361 net7.n1934 net7.n1933 0.189
R28362 net7.n1572 net7.n1571 0.189
R28363 net7.n1210 net7.n1209 0.189
R28364 net7.n848 net7.n847 0.189
R28365 net7.n486 net7.n485 0.189
R28366 net7.n125 net7.n124 0.189
R28367 net7.n3805 net7.n3804 0.189
R28368 net7.n3821 net7.n3820 0.189
R28369 net7.n4166 net7.n4165 0.189
R28370 net7.n4182 net7.n4181 0.189
R28371 net7.n4528 net7.n4527 0.189
R28372 net7.n4544 net7.n4543 0.189
R28373 net7.n4890 net7.n4889 0.189
R28374 net7.n4906 net7.n4905 0.189
R28375 net7.n5252 net7.n5251 0.189
R28376 net7.n5268 net7.n5267 0.189
R28377 net7.n5614 net7.n5613 0.189
R28378 net7.n5630 net7.n5629 0.189
R28379 net7.n5976 net7.n5975 0.189
R28380 net7.n5992 net7.n5991 0.189
R28381 net7.n6338 net7.n6337 0.189
R28382 net7.n6354 net7.n6353 0.189
R28383 net7.n6700 net7.n6699 0.189
R28384 net7.n6716 net7.n6715 0.189
R28385 net7.n7062 net7.n7061 0.189
R28386 net7.n7078 net7.n7077 0.189
R28387 net7.n3527 net7.n3526 0.188
R28388 net7.n3165 net7.n3164 0.188
R28389 net7.n2803 net7.n2802 0.188
R28390 net7.n2441 net7.n2440 0.188
R28391 net7.n2079 net7.n2078 0.188
R28392 net7.n1717 net7.n1716 0.188
R28393 net7.n1355 net7.n1354 0.188
R28394 net7.n993 net7.n992 0.188
R28395 net7.n631 net7.n630 0.188
R28396 net7.n270 net7.n269 0.188
R28397 net7.n6513 net7.n6151 0.182
R28398 net7.n5789 net7.n5427 0.182
R28399 net7.n5065 net7.n4703 0.182
R28400 net7.n3403 net7.n3402 0.166
R28401 net7.n3041 net7.n3040 0.166
R28402 net7.n2679 net7.n2678 0.166
R28403 net7.n2317 net7.n2316 0.166
R28404 net7.n1955 net7.n1954 0.166
R28405 net7.n1593 net7.n1592 0.166
R28406 net7.n1231 net7.n1230 0.166
R28407 net7.n869 net7.n868 0.166
R28408 net7.n507 net7.n506 0.166
R28409 net7.n146 net7.n145 0.166
R28410 net7.n3779 net7.n3778 0.166
R28411 net7.n3911 net7.n3910 0.166
R28412 net7.n4140 net7.n4139 0.166
R28413 net7.n4272 net7.n4271 0.166
R28414 net7.n4502 net7.n4501 0.166
R28415 net7.n4634 net7.n4633 0.166
R28416 net7.n4864 net7.n4863 0.166
R28417 net7.n4996 net7.n4995 0.166
R28418 net7.n5226 net7.n5225 0.166
R28419 net7.n5358 net7.n5357 0.166
R28420 net7.n5588 net7.n5587 0.166
R28421 net7.n5720 net7.n5719 0.166
R28422 net7.n5950 net7.n5949 0.166
R28423 net7.n6082 net7.n6081 0.166
R28424 net7.n6312 net7.n6311 0.166
R28425 net7.n6444 net7.n6443 0.166
R28426 net7.n6674 net7.n6673 0.166
R28427 net7.n6806 net7.n6805 0.166
R28428 net7.n7036 net7.n7035 0.166
R28429 net7.n7168 net7.n7167 0.166
R28430 net7.n3551 net7.n3550 0.166
R28431 net7.n3189 net7.n3188 0.166
R28432 net7.n2827 net7.n2826 0.166
R28433 net7.n2465 net7.n2464 0.166
R28434 net7.n2103 net7.n2102 0.166
R28435 net7.n1741 net7.n1740 0.166
R28436 net7.n1379 net7.n1378 0.166
R28437 net7.n1017 net7.n1016 0.166
R28438 net7.n655 net7.n654 0.166
R28439 net7.n294 net7.n293 0.166
R28440 net7.n3280 net7.n3279 0.133
R28441 net7.n2918 net7.n2917 0.133
R28442 net7.n2556 net7.n2555 0.133
R28443 net7.n2194 net7.n2193 0.133
R28444 net7.n1832 net7.n1831 0.133
R28445 net7.n1470 net7.n1469 0.133
R28446 net7.n1108 net7.n1107 0.133
R28447 net7.n746 net7.n745 0.133
R28448 net7.n384 net7.n383 0.133
R28449 net7.n23 net7.n22 0.133
R28450 net7.n3582 net7.n3581 0.132
R28451 net7.n3220 net7.n3219 0.132
R28452 net7.n2858 net7.n2857 0.132
R28453 net7.n2496 net7.n2495 0.132
R28454 net7.n2134 net7.n2133 0.132
R28455 net7.n1772 net7.n1771 0.132
R28456 net7.n1410 net7.n1409 0.132
R28457 net7.n1048 net7.n1047 0.132
R28458 net7.n686 net7.n685 0.132
R28459 net7.n325 net7.n324 0.132
R28460 net7.n3635 net7.n3634 0.132
R28461 net7.n3947 net7.n3946 0.132
R28462 net7.n3996 net7.n3995 0.132
R28463 net7.n4308 net7.n4307 0.132
R28464 net7.n4358 net7.n4357 0.132
R28465 net7.n4670 net7.n4669 0.132
R28466 net7.n4720 net7.n4719 0.132
R28467 net7.n5032 net7.n5031 0.132
R28468 net7.n5082 net7.n5081 0.132
R28469 net7.n5394 net7.n5393 0.132
R28470 net7.n5444 net7.n5443 0.132
R28471 net7.n5756 net7.n5755 0.132
R28472 net7.n5806 net7.n5805 0.132
R28473 net7.n6118 net7.n6117 0.132
R28474 net7.n6168 net7.n6167 0.132
R28475 net7.n6480 net7.n6479 0.132
R28476 net7.n6530 net7.n6529 0.132
R28477 net7.n6842 net7.n6841 0.132
R28478 net7.n6892 net7.n6891 0.132
R28479 net7.n7204 net7.n7203 0.132
R28480 net7.n3290 net7.n3289 0.121
R28481 net7.n2928 net7.n2927 0.121
R28482 net7.n2566 net7.n2565 0.121
R28483 net7.n2204 net7.n2203 0.121
R28484 net7.n1842 net7.n1841 0.121
R28485 net7.n1480 net7.n1479 0.121
R28486 net7.n1118 net7.n1117 0.121
R28487 net7.n756 net7.n755 0.121
R28488 net7.n394 net7.n393 0.121
R28489 net7.n33 net7.n32 0.121
R28490 net7.n3632 net7.n3631 0.121
R28491 net7.n3957 net7.n3956 0.121
R28492 net7.n3993 net7.n3992 0.121
R28493 net7.n4318 net7.n4317 0.121
R28494 net7.n4355 net7.n4354 0.121
R28495 net7.n4680 net7.n4679 0.121
R28496 net7.n4717 net7.n4716 0.121
R28497 net7.n5042 net7.n5041 0.121
R28498 net7.n5079 net7.n5078 0.121
R28499 net7.n5404 net7.n5403 0.121
R28500 net7.n5441 net7.n5440 0.121
R28501 net7.n5766 net7.n5765 0.121
R28502 net7.n5803 net7.n5802 0.121
R28503 net7.n6128 net7.n6127 0.121
R28504 net7.n6165 net7.n6164 0.121
R28505 net7.n6490 net7.n6489 0.121
R28506 net7.n6527 net7.n6526 0.121
R28507 net7.n6852 net7.n6851 0.121
R28508 net7.n6889 net7.n6888 0.121
R28509 net7.n7214 net7.n7213 0.121
R28510 net7.n3511 net7.n3510 0.121
R28511 net7.n3149 net7.n3148 0.121
R28512 net7.n2787 net7.n2786 0.121
R28513 net7.n2425 net7.n2424 0.121
R28514 net7.n2063 net7.n2062 0.121
R28515 net7.n1701 net7.n1700 0.121
R28516 net7.n1339 net7.n1338 0.121
R28517 net7.n977 net7.n976 0.121
R28518 net7.n615 net7.n614 0.121
R28519 net7.n254 net7.n253 0.121
R28520 net7.n2894 net7.n2532 0.116
R28521 net7.n2170 net7.n1808 0.116
R28522 net7.n1446 net7.n1084 0.116
R28523 net7.n7237 net7.n6875 0.091
R28524 net7.n6875 net7.n6513 0.091
R28525 net7.n6151 net7.n5789 0.091
R28526 net7.n5427 net7.n5065 0.091
R28527 net7.n4703 net7.n4341 0.091
R28528 net7.n3618 net7.n3256 0.058
R28529 net7.n3256 net7.n2894 0.058
R28530 net7.n2532 net7.n2170 0.058
R28531 net7.n1808 net7.n1446 0.058
R28532 net7.n1084 net7.n722 0.058
R28533 net7.n3488 net7.n3487 0.049
R28534 net7.n3483 net7.n3475 0.049
R28535 net7.n3439 net7.n3430 0.049
R28536 net7.n3350 net7.n3335 0.049
R28537 net7.n3126 net7.n3125 0.049
R28538 net7.n3121 net7.n3113 0.049
R28539 net7.n3077 net7.n3068 0.049
R28540 net7.n2988 net7.n2973 0.049
R28541 net7.n2764 net7.n2763 0.049
R28542 net7.n2759 net7.n2751 0.049
R28543 net7.n2715 net7.n2706 0.049
R28544 net7.n2626 net7.n2611 0.049
R28545 net7.n2402 net7.n2401 0.049
R28546 net7.n2397 net7.n2389 0.049
R28547 net7.n2353 net7.n2344 0.049
R28548 net7.n2264 net7.n2249 0.049
R28549 net7.n2040 net7.n2039 0.049
R28550 net7.n2035 net7.n2027 0.049
R28551 net7.n1991 net7.n1982 0.049
R28552 net7.n1902 net7.n1887 0.049
R28553 net7.n1678 net7.n1677 0.049
R28554 net7.n1673 net7.n1665 0.049
R28555 net7.n1629 net7.n1620 0.049
R28556 net7.n1540 net7.n1525 0.049
R28557 net7.n1316 net7.n1315 0.049
R28558 net7.n1311 net7.n1303 0.049
R28559 net7.n1267 net7.n1258 0.049
R28560 net7.n1178 net7.n1163 0.049
R28561 net7.n954 net7.n953 0.049
R28562 net7.n949 net7.n941 0.049
R28563 net7.n905 net7.n896 0.049
R28564 net7.n816 net7.n801 0.049
R28565 net7.n592 net7.n591 0.049
R28566 net7.n587 net7.n579 0.049
R28567 net7.n543 net7.n534 0.049
R28568 net7.n454 net7.n439 0.049
R28569 net7.n231 net7.n230 0.049
R28570 net7.n226 net7.n218 0.049
R28571 net7.n182 net7.n173 0.049
R28572 net7.n93 net7.n78 0.049
R28573 net7.n3840 net7.n3775 0.049
R28574 net7.n3726 net7.n3717 0.049
R28575 net7.n3771 net7.n3762 0.049
R28576 net7.n3875 net7.n3869 0.049
R28577 net7.n4201 net7.n4136 0.049
R28578 net7.n4087 net7.n4078 0.049
R28579 net7.n4132 net7.n4123 0.049
R28580 net7.n4236 net7.n4230 0.049
R28581 net7.n4563 net7.n4498 0.049
R28582 net7.n4449 net7.n4440 0.049
R28583 net7.n4494 net7.n4485 0.049
R28584 net7.n4598 net7.n4592 0.049
R28585 net7.n4925 net7.n4860 0.049
R28586 net7.n4811 net7.n4802 0.049
R28587 net7.n4856 net7.n4847 0.049
R28588 net7.n4960 net7.n4954 0.049
R28589 net7.n5287 net7.n5222 0.049
R28590 net7.n5173 net7.n5164 0.049
R28591 net7.n5218 net7.n5209 0.049
R28592 net7.n5322 net7.n5316 0.049
R28593 net7.n5649 net7.n5584 0.049
R28594 net7.n5535 net7.n5526 0.049
R28595 net7.n5580 net7.n5571 0.049
R28596 net7.n5684 net7.n5678 0.049
R28597 net7.n6011 net7.n5946 0.049
R28598 net7.n5897 net7.n5888 0.049
R28599 net7.n5942 net7.n5933 0.049
R28600 net7.n6046 net7.n6040 0.049
R28601 net7.n6373 net7.n6308 0.049
R28602 net7.n6259 net7.n6250 0.049
R28603 net7.n6304 net7.n6295 0.049
R28604 net7.n6408 net7.n6402 0.049
R28605 net7.n6735 net7.n6670 0.049
R28606 net7.n6621 net7.n6612 0.049
R28607 net7.n6666 net7.n6657 0.049
R28608 net7.n6770 net7.n6764 0.049
R28609 net7.n7097 net7.n7032 0.049
R28610 net7.n6983 net7.n6974 0.049
R28611 net7.n7028 net7.n7019 0.049
R28612 net7.n7132 net7.n7126 0.049
R28613 net7.n3607 net7.n3606 0.047
R28614 net7.n3588 net7.n3586 0.047
R28615 net7.n3586 net7.n3585 0.047
R28616 net7.n3578 net7.n3576 0.047
R28617 net7.n3530 net7.n3529 0.047
R28618 net7.n3385 net7.n3384 0.047
R28619 net7.n3277 net7.n3275 0.047
R28620 net7.n3282 net7.n3281 0.047
R28621 net7.n3285 net7.n3283 0.047
R28622 net7.n3307 net7.n3306 0.047
R28623 net7.n3445 net7.n3444 0.047
R28624 net7.n3245 net7.n3244 0.047
R28625 net7.n3226 net7.n3224 0.047
R28626 net7.n3224 net7.n3223 0.047
R28627 net7.n3216 net7.n3214 0.047
R28628 net7.n3168 net7.n3167 0.047
R28629 net7.n3023 net7.n3022 0.047
R28630 net7.n2915 net7.n2913 0.047
R28631 net7.n2920 net7.n2919 0.047
R28632 net7.n2923 net7.n2921 0.047
R28633 net7.n2945 net7.n2944 0.047
R28634 net7.n3083 net7.n3082 0.047
R28635 net7.n2883 net7.n2882 0.047
R28636 net7.n2864 net7.n2862 0.047
R28637 net7.n2862 net7.n2861 0.047
R28638 net7.n2854 net7.n2852 0.047
R28639 net7.n2806 net7.n2805 0.047
R28640 net7.n2661 net7.n2660 0.047
R28641 net7.n2553 net7.n2551 0.047
R28642 net7.n2558 net7.n2557 0.047
R28643 net7.n2561 net7.n2559 0.047
R28644 net7.n2583 net7.n2582 0.047
R28645 net7.n2721 net7.n2720 0.047
R28646 net7.n2521 net7.n2520 0.047
R28647 net7.n2502 net7.n2500 0.047
R28648 net7.n2500 net7.n2499 0.047
R28649 net7.n2492 net7.n2490 0.047
R28650 net7.n2444 net7.n2443 0.047
R28651 net7.n2299 net7.n2298 0.047
R28652 net7.n2191 net7.n2189 0.047
R28653 net7.n2196 net7.n2195 0.047
R28654 net7.n2199 net7.n2197 0.047
R28655 net7.n2221 net7.n2220 0.047
R28656 net7.n2359 net7.n2358 0.047
R28657 net7.n2159 net7.n2158 0.047
R28658 net7.n2140 net7.n2138 0.047
R28659 net7.n2138 net7.n2137 0.047
R28660 net7.n2130 net7.n2128 0.047
R28661 net7.n2082 net7.n2081 0.047
R28662 net7.n1937 net7.n1936 0.047
R28663 net7.n1829 net7.n1827 0.047
R28664 net7.n1834 net7.n1833 0.047
R28665 net7.n1837 net7.n1835 0.047
R28666 net7.n1859 net7.n1858 0.047
R28667 net7.n1997 net7.n1996 0.047
R28668 net7.n1797 net7.n1796 0.047
R28669 net7.n1778 net7.n1776 0.047
R28670 net7.n1776 net7.n1775 0.047
R28671 net7.n1768 net7.n1766 0.047
R28672 net7.n1720 net7.n1719 0.047
R28673 net7.n1575 net7.n1574 0.047
R28674 net7.n1467 net7.n1465 0.047
R28675 net7.n1472 net7.n1471 0.047
R28676 net7.n1475 net7.n1473 0.047
R28677 net7.n1497 net7.n1496 0.047
R28678 net7.n1635 net7.n1634 0.047
R28679 net7.n1435 net7.n1434 0.047
R28680 net7.n1416 net7.n1414 0.047
R28681 net7.n1414 net7.n1413 0.047
R28682 net7.n1406 net7.n1404 0.047
R28683 net7.n1358 net7.n1357 0.047
R28684 net7.n1213 net7.n1212 0.047
R28685 net7.n1105 net7.n1103 0.047
R28686 net7.n1110 net7.n1109 0.047
R28687 net7.n1113 net7.n1111 0.047
R28688 net7.n1135 net7.n1134 0.047
R28689 net7.n1273 net7.n1272 0.047
R28690 net7.n1073 net7.n1072 0.047
R28691 net7.n1054 net7.n1052 0.047
R28692 net7.n1052 net7.n1051 0.047
R28693 net7.n1044 net7.n1042 0.047
R28694 net7.n996 net7.n995 0.047
R28695 net7.n851 net7.n850 0.047
R28696 net7.n743 net7.n741 0.047
R28697 net7.n748 net7.n747 0.047
R28698 net7.n751 net7.n749 0.047
R28699 net7.n773 net7.n772 0.047
R28700 net7.n911 net7.n910 0.047
R28701 net7.n711 net7.n710 0.047
R28702 net7.n692 net7.n690 0.047
R28703 net7.n690 net7.n689 0.047
R28704 net7.n682 net7.n680 0.047
R28705 net7.n634 net7.n633 0.047
R28706 net7.n489 net7.n488 0.047
R28707 net7.n381 net7.n379 0.047
R28708 net7.n386 net7.n385 0.047
R28709 net7.n389 net7.n387 0.047
R28710 net7.n411 net7.n410 0.047
R28711 net7.n549 net7.n548 0.047
R28712 net7.n350 net7.n349 0.047
R28713 net7.n331 net7.n329 0.047
R28714 net7.n329 net7.n328 0.047
R28715 net7.n321 net7.n319 0.047
R28716 net7.n273 net7.n272 0.047
R28717 net7.n128 net7.n127 0.047
R28718 net7.n20 net7.n18 0.047
R28719 net7.n25 net7.n24 0.047
R28720 net7.n28 net7.n26 0.047
R28721 net7.n50 net7.n49 0.047
R28722 net7.n188 net7.n187 0.047
R28723 net7.n3691 net7.n3690 0.047
R28724 net7.n3674 net7.n3672 0.047
R28725 net7.n3672 net7.n3671 0.047
R28726 net7.n3667 net7.n3665 0.047
R28727 net7.n3803 net7.n3802 0.047
R28728 net7.n3824 net7.n3823 0.047
R28729 net7.n3944 net7.n3942 0.047
R28730 net7.n3949 net7.n3948 0.047
R28731 net7.n3952 net7.n3950 0.047
R28732 net7.n3974 net7.n3973 0.047
R28733 net7.n3882 net7.n3880 0.047
R28734 net7.n4052 net7.n4051 0.047
R28735 net7.n4035 net7.n4033 0.047
R28736 net7.n4033 net7.n4032 0.047
R28737 net7.n4028 net7.n4026 0.047
R28738 net7.n4164 net7.n4163 0.047
R28739 net7.n4185 net7.n4184 0.047
R28740 net7.n4305 net7.n4303 0.047
R28741 net7.n4310 net7.n4309 0.047
R28742 net7.n4313 net7.n4311 0.047
R28743 net7.n4335 net7.n4334 0.047
R28744 net7.n4243 net7.n4241 0.047
R28745 net7.n4414 net7.n4413 0.047
R28746 net7.n4397 net7.n4395 0.047
R28747 net7.n4395 net7.n4394 0.047
R28748 net7.n4390 net7.n4388 0.047
R28749 net7.n4526 net7.n4525 0.047
R28750 net7.n4547 net7.n4546 0.047
R28751 net7.n4667 net7.n4665 0.047
R28752 net7.n4672 net7.n4671 0.047
R28753 net7.n4675 net7.n4673 0.047
R28754 net7.n4697 net7.n4696 0.047
R28755 net7.n4605 net7.n4603 0.047
R28756 net7.n4776 net7.n4775 0.047
R28757 net7.n4759 net7.n4757 0.047
R28758 net7.n4757 net7.n4756 0.047
R28759 net7.n4752 net7.n4750 0.047
R28760 net7.n4888 net7.n4887 0.047
R28761 net7.n4909 net7.n4908 0.047
R28762 net7.n5029 net7.n5027 0.047
R28763 net7.n5034 net7.n5033 0.047
R28764 net7.n5037 net7.n5035 0.047
R28765 net7.n5059 net7.n5058 0.047
R28766 net7.n4967 net7.n4965 0.047
R28767 net7.n5138 net7.n5137 0.047
R28768 net7.n5121 net7.n5119 0.047
R28769 net7.n5119 net7.n5118 0.047
R28770 net7.n5114 net7.n5112 0.047
R28771 net7.n5250 net7.n5249 0.047
R28772 net7.n5271 net7.n5270 0.047
R28773 net7.n5391 net7.n5389 0.047
R28774 net7.n5396 net7.n5395 0.047
R28775 net7.n5399 net7.n5397 0.047
R28776 net7.n5421 net7.n5420 0.047
R28777 net7.n5329 net7.n5327 0.047
R28778 net7.n5500 net7.n5499 0.047
R28779 net7.n5483 net7.n5481 0.047
R28780 net7.n5481 net7.n5480 0.047
R28781 net7.n5476 net7.n5474 0.047
R28782 net7.n5612 net7.n5611 0.047
R28783 net7.n5633 net7.n5632 0.047
R28784 net7.n5753 net7.n5751 0.047
R28785 net7.n5758 net7.n5757 0.047
R28786 net7.n5761 net7.n5759 0.047
R28787 net7.n5783 net7.n5782 0.047
R28788 net7.n5691 net7.n5689 0.047
R28789 net7.n5862 net7.n5861 0.047
R28790 net7.n5845 net7.n5843 0.047
R28791 net7.n5843 net7.n5842 0.047
R28792 net7.n5838 net7.n5836 0.047
R28793 net7.n5974 net7.n5973 0.047
R28794 net7.n5995 net7.n5994 0.047
R28795 net7.n6115 net7.n6113 0.047
R28796 net7.n6120 net7.n6119 0.047
R28797 net7.n6123 net7.n6121 0.047
R28798 net7.n6145 net7.n6144 0.047
R28799 net7.n6053 net7.n6051 0.047
R28800 net7.n6224 net7.n6223 0.047
R28801 net7.n6207 net7.n6205 0.047
R28802 net7.n6205 net7.n6204 0.047
R28803 net7.n6200 net7.n6198 0.047
R28804 net7.n6336 net7.n6335 0.047
R28805 net7.n6357 net7.n6356 0.047
R28806 net7.n6477 net7.n6475 0.047
R28807 net7.n6482 net7.n6481 0.047
R28808 net7.n6485 net7.n6483 0.047
R28809 net7.n6507 net7.n6506 0.047
R28810 net7.n6415 net7.n6413 0.047
R28811 net7.n6586 net7.n6585 0.047
R28812 net7.n6569 net7.n6567 0.047
R28813 net7.n6567 net7.n6566 0.047
R28814 net7.n6562 net7.n6560 0.047
R28815 net7.n6698 net7.n6697 0.047
R28816 net7.n6719 net7.n6718 0.047
R28817 net7.n6839 net7.n6837 0.047
R28818 net7.n6844 net7.n6843 0.047
R28819 net7.n6847 net7.n6845 0.047
R28820 net7.n6869 net7.n6868 0.047
R28821 net7.n6777 net7.n6775 0.047
R28822 net7.n6948 net7.n6947 0.047
R28823 net7.n6931 net7.n6929 0.047
R28824 net7.n6929 net7.n6928 0.047
R28825 net7.n6924 net7.n6922 0.047
R28826 net7.n7060 net7.n7059 0.047
R28827 net7.n7081 net7.n7080 0.047
R28828 net7.n7201 net7.n7199 0.047
R28829 net7.n7206 net7.n7205 0.047
R28830 net7.n7209 net7.n7207 0.047
R28831 net7.n7231 net7.n7230 0.047
R28832 net7.n7139 net7.n7137 0.047
R28833 net7.n3532 net7.n3531 0.045
R28834 net7.n3386 net7.n3385 0.045
R28835 net7.n3170 net7.n3169 0.045
R28836 net7.n3024 net7.n3023 0.045
R28837 net7.n2808 net7.n2807 0.045
R28838 net7.n2662 net7.n2661 0.045
R28839 net7.n2446 net7.n2445 0.045
R28840 net7.n2300 net7.n2299 0.045
R28841 net7.n2084 net7.n2083 0.045
R28842 net7.n1938 net7.n1937 0.045
R28843 net7.n1722 net7.n1721 0.045
R28844 net7.n1576 net7.n1575 0.045
R28845 net7.n1360 net7.n1359 0.045
R28846 net7.n1214 net7.n1213 0.045
R28847 net7.n998 net7.n997 0.045
R28848 net7.n852 net7.n851 0.045
R28849 net7.n636 net7.n635 0.045
R28850 net7.n490 net7.n489 0.045
R28851 net7.n275 net7.n274 0.045
R28852 net7.n129 net7.n128 0.045
R28853 net7.n3801 net7.n3800 0.045
R28854 net7.n3825 net7.n3824 0.045
R28855 net7.n4162 net7.n4161 0.045
R28856 net7.n4186 net7.n4185 0.045
R28857 net7.n4524 net7.n4523 0.045
R28858 net7.n4548 net7.n4547 0.045
R28859 net7.n4886 net7.n4885 0.045
R28860 net7.n4910 net7.n4909 0.045
R28861 net7.n5248 net7.n5247 0.045
R28862 net7.n5272 net7.n5271 0.045
R28863 net7.n5610 net7.n5609 0.045
R28864 net7.n5634 net7.n5633 0.045
R28865 net7.n5972 net7.n5971 0.045
R28866 net7.n5996 net7.n5995 0.045
R28867 net7.n6334 net7.n6333 0.045
R28868 net7.n6358 net7.n6357 0.045
R28869 net7.n6696 net7.n6695 0.045
R28870 net7.n6720 net7.n6719 0.045
R28871 net7.n7058 net7.n7057 0.045
R28872 net7.n7082 net7.n7081 0.045
R28873 net7.n3555 net7.n3554 0.043
R28874 net7.n3346 net7.n3340 0.043
R28875 net7.n3438 net7.n3437 0.043
R28876 net7.n3348 net7.n3347 0.043
R28877 net7.n3333 net7.n3332 0.043
R28878 net7.n3193 net7.n3192 0.043
R28879 net7.n2984 net7.n2978 0.043
R28880 net7.n3076 net7.n3075 0.043
R28881 net7.n2986 net7.n2985 0.043
R28882 net7.n2971 net7.n2970 0.043
R28883 net7.n2831 net7.n2830 0.043
R28884 net7.n2622 net7.n2616 0.043
R28885 net7.n2714 net7.n2713 0.043
R28886 net7.n2624 net7.n2623 0.043
R28887 net7.n2609 net7.n2608 0.043
R28888 net7.n2469 net7.n2468 0.043
R28889 net7.n2260 net7.n2254 0.043
R28890 net7.n2352 net7.n2351 0.043
R28891 net7.n2262 net7.n2261 0.043
R28892 net7.n2247 net7.n2246 0.043
R28893 net7.n2107 net7.n2106 0.043
R28894 net7.n1898 net7.n1892 0.043
R28895 net7.n1990 net7.n1989 0.043
R28896 net7.n1900 net7.n1899 0.043
R28897 net7.n1885 net7.n1884 0.043
R28898 net7.n1745 net7.n1744 0.043
R28899 net7.n1536 net7.n1530 0.043
R28900 net7.n1628 net7.n1627 0.043
R28901 net7.n1538 net7.n1537 0.043
R28902 net7.n1523 net7.n1522 0.043
R28903 net7.n1383 net7.n1382 0.043
R28904 net7.n1174 net7.n1168 0.043
R28905 net7.n1266 net7.n1265 0.043
R28906 net7.n1176 net7.n1175 0.043
R28907 net7.n1161 net7.n1160 0.043
R28908 net7.n1021 net7.n1020 0.043
R28909 net7.n812 net7.n806 0.043
R28910 net7.n904 net7.n903 0.043
R28911 net7.n814 net7.n813 0.043
R28912 net7.n799 net7.n798 0.043
R28913 net7.n659 net7.n658 0.043
R28914 net7.n450 net7.n444 0.043
R28915 net7.n542 net7.n541 0.043
R28916 net7.n452 net7.n451 0.043
R28917 net7.n437 net7.n436 0.043
R28918 net7.n298 net7.n297 0.043
R28919 net7.n89 net7.n83 0.043
R28920 net7.n181 net7.n180 0.043
R28921 net7.n91 net7.n90 0.043
R28922 net7.n76 net7.n75 0.043
R28923 net7.n3811 net7.n3810 0.043
R28924 net7.n3932 net7.n3928 0.043
R28925 net7.n3714 net7.n3713 0.043
R28926 net7.n3732 net7.n3731 0.043
R28927 net7.n4172 net7.n4171 0.043
R28928 net7.n4293 net7.n4289 0.043
R28929 net7.n4075 net7.n4074 0.043
R28930 net7.n4093 net7.n4092 0.043
R28931 net7.n4534 net7.n4533 0.043
R28932 net7.n4655 net7.n4651 0.043
R28933 net7.n4437 net7.n4436 0.043
R28934 net7.n4455 net7.n4454 0.043
R28935 net7.n4896 net7.n4895 0.043
R28936 net7.n5017 net7.n5013 0.043
R28937 net7.n4799 net7.n4798 0.043
R28938 net7.n4817 net7.n4816 0.043
R28939 net7.n5258 net7.n5257 0.043
R28940 net7.n5379 net7.n5375 0.043
R28941 net7.n5161 net7.n5160 0.043
R28942 net7.n5179 net7.n5178 0.043
R28943 net7.n5620 net7.n5619 0.043
R28944 net7.n5741 net7.n5737 0.043
R28945 net7.n5523 net7.n5522 0.043
R28946 net7.n5541 net7.n5540 0.043
R28947 net7.n5982 net7.n5981 0.043
R28948 net7.n6103 net7.n6099 0.043
R28949 net7.n5885 net7.n5884 0.043
R28950 net7.n5903 net7.n5902 0.043
R28951 net7.n6344 net7.n6343 0.043
R28952 net7.n6465 net7.n6461 0.043
R28953 net7.n6247 net7.n6246 0.043
R28954 net7.n6265 net7.n6264 0.043
R28955 net7.n6706 net7.n6705 0.043
R28956 net7.n6827 net7.n6823 0.043
R28957 net7.n6609 net7.n6608 0.043
R28958 net7.n6627 net7.n6626 0.043
R28959 net7.n7068 net7.n7067 0.043
R28960 net7.n7189 net7.n7185 0.043
R28961 net7.n6971 net7.n6970 0.043
R28962 net7.n6989 net7.n6988 0.043
R28963 net7.n3610 net7.n3607 0.043
R28964 net7.n3248 net7.n3245 0.043
R28965 net7.n2886 net7.n2883 0.043
R28966 net7.n2524 net7.n2521 0.043
R28967 net7.n2162 net7.n2159 0.043
R28968 net7.n1800 net7.n1797 0.043
R28969 net7.n1438 net7.n1435 0.043
R28970 net7.n1076 net7.n1073 0.043
R28971 net7.n714 net7.n711 0.043
R28972 net7.n353 net7.n350 0.043
R28973 net7.n3693 net7.n3691 0.043
R28974 net7.n4054 net7.n4052 0.043
R28975 net7.n4416 net7.n4414 0.043
R28976 net7.n4778 net7.n4776 0.043
R28977 net7.n5140 net7.n5138 0.043
R28978 net7.n5502 net7.n5500 0.043
R28979 net7.n5864 net7.n5862 0.043
R28980 net7.n6226 net7.n6224 0.043
R28981 net7.n6588 net7.n6586 0.043
R28982 net7.n6950 net7.n6948 0.043
R28983 net7.n3575 net7.n3574 0.041
R28984 net7.n3568 net7.n3564 0.041
R28985 net7.n3376 net7.n3375 0.041
R28986 net7.n3400 net7.n3399 0.041
R28987 net7.n3297 net7.n3296 0.041
R28988 net7.n3482 net7.n3481 0.041
R28989 net7.n3356 net7.n3355 0.041
R28990 net7.n3213 net7.n3212 0.041
R28991 net7.n3206 net7.n3202 0.041
R28992 net7.n3014 net7.n3013 0.041
R28993 net7.n3038 net7.n3037 0.041
R28994 net7.n2935 net7.n2934 0.041
R28995 net7.n3120 net7.n3119 0.041
R28996 net7.n2994 net7.n2993 0.041
R28997 net7.n2851 net7.n2850 0.041
R28998 net7.n2844 net7.n2840 0.041
R28999 net7.n2652 net7.n2651 0.041
R29000 net7.n2676 net7.n2675 0.041
R29001 net7.n2573 net7.n2572 0.041
R29002 net7.n2758 net7.n2757 0.041
R29003 net7.n2632 net7.n2631 0.041
R29004 net7.n2489 net7.n2488 0.041
R29005 net7.n2482 net7.n2478 0.041
R29006 net7.n2290 net7.n2289 0.041
R29007 net7.n2314 net7.n2313 0.041
R29008 net7.n2211 net7.n2210 0.041
R29009 net7.n2396 net7.n2395 0.041
R29010 net7.n2270 net7.n2269 0.041
R29011 net7.n2127 net7.n2126 0.041
R29012 net7.n2120 net7.n2116 0.041
R29013 net7.n1928 net7.n1927 0.041
R29014 net7.n1952 net7.n1951 0.041
R29015 net7.n1849 net7.n1848 0.041
R29016 net7.n2034 net7.n2033 0.041
R29017 net7.n1908 net7.n1907 0.041
R29018 net7.n1765 net7.n1764 0.041
R29019 net7.n1758 net7.n1754 0.041
R29020 net7.n1566 net7.n1565 0.041
R29021 net7.n1590 net7.n1589 0.041
R29022 net7.n1487 net7.n1486 0.041
R29023 net7.n1672 net7.n1671 0.041
R29024 net7.n1546 net7.n1545 0.041
R29025 net7.n1403 net7.n1402 0.041
R29026 net7.n1396 net7.n1392 0.041
R29027 net7.n1204 net7.n1203 0.041
R29028 net7.n1228 net7.n1227 0.041
R29029 net7.n1125 net7.n1124 0.041
R29030 net7.n1310 net7.n1309 0.041
R29031 net7.n1184 net7.n1183 0.041
R29032 net7.n1041 net7.n1040 0.041
R29033 net7.n1034 net7.n1030 0.041
R29034 net7.n842 net7.n841 0.041
R29035 net7.n866 net7.n865 0.041
R29036 net7.n763 net7.n762 0.041
R29037 net7.n948 net7.n947 0.041
R29038 net7.n822 net7.n821 0.041
R29039 net7.n679 net7.n678 0.041
R29040 net7.n672 net7.n668 0.041
R29041 net7.n480 net7.n479 0.041
R29042 net7.n504 net7.n503 0.041
R29043 net7.n401 net7.n400 0.041
R29044 net7.n586 net7.n585 0.041
R29045 net7.n460 net7.n459 0.041
R29046 net7.n318 net7.n317 0.041
R29047 net7.n311 net7.n307 0.041
R29048 net7.n119 net7.n118 0.041
R29049 net7.n143 net7.n142 0.041
R29050 net7.n40 net7.n39 0.041
R29051 net7.n225 net7.n224 0.041
R29052 net7.n99 net7.n98 0.041
R29053 net7.n3664 net7.n3663 0.041
R29054 net7.n3657 net7.n3656 0.041
R29055 net7.n3815 net7.n3814 0.041
R29056 net7.n3915 net7.n3914 0.041
R29057 net7.n3964 net7.n3963 0.041
R29058 net7.n3722 net7.n3721 0.041
R29059 net7.n3770 net7.n3766 0.041
R29060 net7.n4025 net7.n4024 0.041
R29061 net7.n4018 net7.n4017 0.041
R29062 net7.n4176 net7.n4175 0.041
R29063 net7.n4276 net7.n4275 0.041
R29064 net7.n4325 net7.n4324 0.041
R29065 net7.n4083 net7.n4082 0.041
R29066 net7.n4131 net7.n4127 0.041
R29067 net7.n4387 net7.n4386 0.041
R29068 net7.n4380 net7.n4379 0.041
R29069 net7.n4538 net7.n4537 0.041
R29070 net7.n4638 net7.n4637 0.041
R29071 net7.n4687 net7.n4686 0.041
R29072 net7.n4445 net7.n4444 0.041
R29073 net7.n4493 net7.n4489 0.041
R29074 net7.n4749 net7.n4748 0.041
R29075 net7.n4742 net7.n4741 0.041
R29076 net7.n4900 net7.n4899 0.041
R29077 net7.n5000 net7.n4999 0.041
R29078 net7.n5049 net7.n5048 0.041
R29079 net7.n4807 net7.n4806 0.041
R29080 net7.n4855 net7.n4851 0.041
R29081 net7.n5111 net7.n5110 0.041
R29082 net7.n5104 net7.n5103 0.041
R29083 net7.n5262 net7.n5261 0.041
R29084 net7.n5362 net7.n5361 0.041
R29085 net7.n5411 net7.n5410 0.041
R29086 net7.n5169 net7.n5168 0.041
R29087 net7.n5217 net7.n5213 0.041
R29088 net7.n5473 net7.n5472 0.041
R29089 net7.n5466 net7.n5465 0.041
R29090 net7.n5624 net7.n5623 0.041
R29091 net7.n5724 net7.n5723 0.041
R29092 net7.n5773 net7.n5772 0.041
R29093 net7.n5531 net7.n5530 0.041
R29094 net7.n5579 net7.n5575 0.041
R29095 net7.n5835 net7.n5834 0.041
R29096 net7.n5828 net7.n5827 0.041
R29097 net7.n5986 net7.n5985 0.041
R29098 net7.n6086 net7.n6085 0.041
R29099 net7.n6135 net7.n6134 0.041
R29100 net7.n5893 net7.n5892 0.041
R29101 net7.n5941 net7.n5937 0.041
R29102 net7.n6197 net7.n6196 0.041
R29103 net7.n6190 net7.n6189 0.041
R29104 net7.n6348 net7.n6347 0.041
R29105 net7.n6448 net7.n6447 0.041
R29106 net7.n6497 net7.n6496 0.041
R29107 net7.n6255 net7.n6254 0.041
R29108 net7.n6303 net7.n6299 0.041
R29109 net7.n6559 net7.n6558 0.041
R29110 net7.n6552 net7.n6551 0.041
R29111 net7.n6710 net7.n6709 0.041
R29112 net7.n6810 net7.n6809 0.041
R29113 net7.n6859 net7.n6858 0.041
R29114 net7.n6617 net7.n6616 0.041
R29115 net7.n6665 net7.n6661 0.041
R29116 net7.n6921 net7.n6920 0.041
R29117 net7.n6914 net7.n6913 0.041
R29118 net7.n7072 net7.n7071 0.041
R29119 net7.n7172 net7.n7171 0.041
R29120 net7.n7221 net7.n7220 0.041
R29121 net7.n6979 net7.n6978 0.041
R29122 net7.n7027 net7.n7023 0.041
R29123 net7.n3977 net7.n3974 0.041
R29124 net7.n4338 net7.n4335 0.041
R29125 net7.n4700 net7.n4697 0.041
R29126 net7.n5062 net7.n5059 0.041
R29127 net7.n5424 net7.n5421 0.041
R29128 net7.n5786 net7.n5783 0.041
R29129 net7.n6148 net7.n6145 0.041
R29130 net7.n6510 net7.n6507 0.041
R29131 net7.n6872 net7.n6869 0.041
R29132 net7.n7234 net7.n7231 0.041
R29133 net7.n3309 net7.n3307 0.041
R29134 net7.n2947 net7.n2945 0.041
R29135 net7.n2585 net7.n2583 0.041
R29136 net7.n2223 net7.n2221 0.041
R29137 net7.n1861 net7.n1859 0.041
R29138 net7.n1499 net7.n1497 0.041
R29139 net7.n1137 net7.n1135 0.041
R29140 net7.n775 net7.n773 0.041
R29141 net7.n413 net7.n411 0.041
R29142 net7.n52 net7.n50 0.041
R29143 net7.n3597 net7.n3596 0.039
R29144 net7.n3553 net7.n3552 0.039
R29145 net7.n3404 net7.n3401 0.039
R29146 net7.n3274 net7.n3273 0.039
R29147 net7.n3334 net7.n3329 0.039
R29148 net7.n3235 net7.n3234 0.039
R29149 net7.n3191 net7.n3190 0.039
R29150 net7.n3042 net7.n3039 0.039
R29151 net7.n2912 net7.n2911 0.039
R29152 net7.n2972 net7.n2967 0.039
R29153 net7.n2873 net7.n2872 0.039
R29154 net7.n2829 net7.n2828 0.039
R29155 net7.n2680 net7.n2677 0.039
R29156 net7.n2550 net7.n2549 0.039
R29157 net7.n2610 net7.n2605 0.039
R29158 net7.n2511 net7.n2510 0.039
R29159 net7.n2467 net7.n2466 0.039
R29160 net7.n2318 net7.n2315 0.039
R29161 net7.n2188 net7.n2187 0.039
R29162 net7.n2248 net7.n2243 0.039
R29163 net7.n2149 net7.n2148 0.039
R29164 net7.n2105 net7.n2104 0.039
R29165 net7.n1956 net7.n1953 0.039
R29166 net7.n1826 net7.n1825 0.039
R29167 net7.n1886 net7.n1881 0.039
R29168 net7.n1787 net7.n1786 0.039
R29169 net7.n1743 net7.n1742 0.039
R29170 net7.n1594 net7.n1591 0.039
R29171 net7.n1464 net7.n1463 0.039
R29172 net7.n1524 net7.n1519 0.039
R29173 net7.n1425 net7.n1424 0.039
R29174 net7.n1381 net7.n1380 0.039
R29175 net7.n1232 net7.n1229 0.039
R29176 net7.n1102 net7.n1101 0.039
R29177 net7.n1162 net7.n1157 0.039
R29178 net7.n1063 net7.n1062 0.039
R29179 net7.n1019 net7.n1018 0.039
R29180 net7.n870 net7.n867 0.039
R29181 net7.n740 net7.n739 0.039
R29182 net7.n800 net7.n795 0.039
R29183 net7.n701 net7.n700 0.039
R29184 net7.n657 net7.n656 0.039
R29185 net7.n508 net7.n505 0.039
R29186 net7.n378 net7.n377 0.039
R29187 net7.n438 net7.n433 0.039
R29188 net7.n340 net7.n339 0.039
R29189 net7.n296 net7.n295 0.039
R29190 net7.n147 net7.n144 0.039
R29191 net7.n17 net7.n16 0.039
R29192 net7.n77 net7.n72 0.039
R29193 net7.n3683 net7.n3682 0.039
R29194 net7.n3780 net7.n3777 0.039
R29195 net7.n3913 net7.n3912 0.039
R29196 net7.n3941 net7.n3940 0.039
R29197 net7.n3874 net7.n3872 0.039
R29198 net7.n4044 net7.n4043 0.039
R29199 net7.n4141 net7.n4138 0.039
R29200 net7.n4274 net7.n4273 0.039
R29201 net7.n4302 net7.n4301 0.039
R29202 net7.n4235 net7.n4233 0.039
R29203 net7.n4406 net7.n4405 0.039
R29204 net7.n4503 net7.n4500 0.039
R29205 net7.n4636 net7.n4635 0.039
R29206 net7.n4664 net7.n4663 0.039
R29207 net7.n4597 net7.n4595 0.039
R29208 net7.n4768 net7.n4767 0.039
R29209 net7.n4865 net7.n4862 0.039
R29210 net7.n4998 net7.n4997 0.039
R29211 net7.n5026 net7.n5025 0.039
R29212 net7.n4959 net7.n4957 0.039
R29213 net7.n5130 net7.n5129 0.039
R29214 net7.n5227 net7.n5224 0.039
R29215 net7.n5360 net7.n5359 0.039
R29216 net7.n5388 net7.n5387 0.039
R29217 net7.n5321 net7.n5319 0.039
R29218 net7.n5492 net7.n5491 0.039
R29219 net7.n5589 net7.n5586 0.039
R29220 net7.n5722 net7.n5721 0.039
R29221 net7.n5750 net7.n5749 0.039
R29222 net7.n5683 net7.n5681 0.039
R29223 net7.n5854 net7.n5853 0.039
R29224 net7.n5951 net7.n5948 0.039
R29225 net7.n6084 net7.n6083 0.039
R29226 net7.n6112 net7.n6111 0.039
R29227 net7.n6045 net7.n6043 0.039
R29228 net7.n6216 net7.n6215 0.039
R29229 net7.n6313 net7.n6310 0.039
R29230 net7.n6446 net7.n6445 0.039
R29231 net7.n6474 net7.n6473 0.039
R29232 net7.n6407 net7.n6405 0.039
R29233 net7.n6578 net7.n6577 0.039
R29234 net7.n6675 net7.n6672 0.039
R29235 net7.n6808 net7.n6807 0.039
R29236 net7.n6836 net7.n6835 0.039
R29237 net7.n6769 net7.n6767 0.039
R29238 net7.n6940 net7.n6939 0.039
R29239 net7.n7037 net7.n7034 0.039
R29240 net7.n7170 net7.n7169 0.039
R29241 net7.n7198 net7.n7197 0.039
R29242 net7.n7131 net7.n7129 0.039
R29243 net7.n3563 net7.n3562 0.037
R29244 net7.n3201 net7.n3200 0.037
R29245 net7.n2839 net7.n2838 0.037
R29246 net7.n2477 net7.n2476 0.037
R29247 net7.n2115 net7.n2114 0.037
R29248 net7.n1753 net7.n1752 0.037
R29249 net7.n1391 net7.n1390 0.037
R29250 net7.n1029 net7.n1028 0.037
R29251 net7.n667 net7.n666 0.037
R29252 net7.n306 net7.n305 0.037
R29253 net7.n3655 net7.n3654 0.037
R29254 net7.n4016 net7.n4015 0.037
R29255 net7.n4378 net7.n4377 0.037
R29256 net7.n4740 net7.n4739 0.037
R29257 net7.n5102 net7.n5101 0.037
R29258 net7.n5464 net7.n5463 0.037
R29259 net7.n5826 net7.n5825 0.037
R29260 net7.n6188 net7.n6187 0.037
R29261 net7.n6550 net7.n6549 0.037
R29262 net7.n6912 net7.n6911 0.037
R29263 net7.n3264 net7.n3263 0.035
R29264 net7.n2902 net7.n2901 0.035
R29265 net7.n2540 net7.n2539 0.035
R29266 net7.n2178 net7.n2177 0.035
R29267 net7.n1816 net7.n1815 0.035
R29268 net7.n1454 net7.n1453 0.035
R29269 net7.n1092 net7.n1091 0.035
R29270 net7.n730 net7.n729 0.035
R29271 net7.n368 net7.n367 0.035
R29272 net7.n7 net7.n6 0.035
R29273 net7.n3927 net7.n3926 0.035
R29274 net7.n3625 net7.n3624 0.035
R29275 net7.n4288 net7.n4287 0.035
R29276 net7.n3986 net7.n3985 0.035
R29277 net7.n4650 net7.n4649 0.035
R29278 net7.n4348 net7.n4347 0.035
R29279 net7.n5012 net7.n5011 0.035
R29280 net7.n4710 net7.n4709 0.035
R29281 net7.n5374 net7.n5373 0.035
R29282 net7.n5072 net7.n5071 0.035
R29283 net7.n5736 net7.n5735 0.035
R29284 net7.n5434 net7.n5433 0.035
R29285 net7.n6098 net7.n6097 0.035
R29286 net7.n5796 net7.n5795 0.035
R29287 net7.n6460 net7.n6459 0.035
R29288 net7.n6158 net7.n6157 0.035
R29289 net7.n6822 net7.n6821 0.035
R29290 net7.n6520 net7.n6519 0.035
R29291 net7.n7184 net7.n7183 0.035
R29292 net7.n6882 net7.n6881 0.035
R29293 net7.n3542 net7.n3541 0.034
R29294 net7.n3374 net7.n3373 0.034
R29295 net7.n3487 net7.n3486 0.034
R29296 net7.n3480 net7.n3479 0.034
R29297 net7.n3436 net7.n3435 0.034
R29298 net7.n3425 net7.n3424 0.034
R29299 net7.n3347 net7.n3338 0.034
R29300 net7.n3332 net7.n3331 0.034
R29301 net7.n3180 net7.n3179 0.034
R29302 net7.n3012 net7.n3011 0.034
R29303 net7.n3125 net7.n3124 0.034
R29304 net7.n3118 net7.n3117 0.034
R29305 net7.n3074 net7.n3073 0.034
R29306 net7.n3063 net7.n3062 0.034
R29307 net7.n2985 net7.n2976 0.034
R29308 net7.n2970 net7.n2969 0.034
R29309 net7.n2818 net7.n2817 0.034
R29310 net7.n2650 net7.n2649 0.034
R29311 net7.n2763 net7.n2762 0.034
R29312 net7.n2756 net7.n2755 0.034
R29313 net7.n2712 net7.n2711 0.034
R29314 net7.n2701 net7.n2700 0.034
R29315 net7.n2623 net7.n2614 0.034
R29316 net7.n2608 net7.n2607 0.034
R29317 net7.n2456 net7.n2455 0.034
R29318 net7.n2288 net7.n2287 0.034
R29319 net7.n2401 net7.n2400 0.034
R29320 net7.n2394 net7.n2393 0.034
R29321 net7.n2350 net7.n2349 0.034
R29322 net7.n2339 net7.n2338 0.034
R29323 net7.n2261 net7.n2252 0.034
R29324 net7.n2246 net7.n2245 0.034
R29325 net7.n2094 net7.n2093 0.034
R29326 net7.n1926 net7.n1925 0.034
R29327 net7.n2039 net7.n2038 0.034
R29328 net7.n2032 net7.n2031 0.034
R29329 net7.n1988 net7.n1987 0.034
R29330 net7.n1977 net7.n1976 0.034
R29331 net7.n1899 net7.n1890 0.034
R29332 net7.n1884 net7.n1883 0.034
R29333 net7.n1732 net7.n1731 0.034
R29334 net7.n1564 net7.n1563 0.034
R29335 net7.n1677 net7.n1676 0.034
R29336 net7.n1670 net7.n1669 0.034
R29337 net7.n1626 net7.n1625 0.034
R29338 net7.n1615 net7.n1614 0.034
R29339 net7.n1537 net7.n1528 0.034
R29340 net7.n1522 net7.n1521 0.034
R29341 net7.n1370 net7.n1369 0.034
R29342 net7.n1202 net7.n1201 0.034
R29343 net7.n1315 net7.n1314 0.034
R29344 net7.n1308 net7.n1307 0.034
R29345 net7.n1264 net7.n1263 0.034
R29346 net7.n1253 net7.n1252 0.034
R29347 net7.n1175 net7.n1166 0.034
R29348 net7.n1160 net7.n1159 0.034
R29349 net7.n1008 net7.n1007 0.034
R29350 net7.n840 net7.n839 0.034
R29351 net7.n953 net7.n952 0.034
R29352 net7.n946 net7.n945 0.034
R29353 net7.n902 net7.n901 0.034
R29354 net7.n891 net7.n890 0.034
R29355 net7.n813 net7.n804 0.034
R29356 net7.n798 net7.n797 0.034
R29357 net7.n646 net7.n645 0.034
R29358 net7.n478 net7.n477 0.034
R29359 net7.n591 net7.n590 0.034
R29360 net7.n584 net7.n583 0.034
R29361 net7.n540 net7.n539 0.034
R29362 net7.n529 net7.n528 0.034
R29363 net7.n451 net7.n442 0.034
R29364 net7.n436 net7.n435 0.034
R29365 net7.n285 net7.n284 0.034
R29366 net7.n117 net7.n116 0.034
R29367 net7.n230 net7.n229 0.034
R29368 net7.n223 net7.n222 0.034
R29369 net7.n179 net7.n178 0.034
R29370 net7.n168 net7.n167 0.034
R29371 net7.n90 net7.n81 0.034
R29372 net7.n75 net7.n74 0.034
R29373 net7.n3793 net7.n3790 0.034
R29374 net7.n3813 net7.n3812 0.034
R29375 net7.n3713 net7.n3712 0.034
R29376 net7.n3720 net7.n3719 0.034
R29377 net7.n3765 net7.n3764 0.034
R29378 net7.n3775 net7.n3774 0.034
R29379 net7.n3871 net7.n3870 0.034
R29380 net7.n3879 net7.n3878 0.034
R29381 net7.n4154 net7.n4151 0.034
R29382 net7.n4174 net7.n4173 0.034
R29383 net7.n4074 net7.n4073 0.034
R29384 net7.n4081 net7.n4080 0.034
R29385 net7.n4126 net7.n4125 0.034
R29386 net7.n4136 net7.n4135 0.034
R29387 net7.n4232 net7.n4231 0.034
R29388 net7.n4240 net7.n4239 0.034
R29389 net7.n4516 net7.n4513 0.034
R29390 net7.n4536 net7.n4535 0.034
R29391 net7.n4436 net7.n4435 0.034
R29392 net7.n4443 net7.n4442 0.034
R29393 net7.n4488 net7.n4487 0.034
R29394 net7.n4498 net7.n4497 0.034
R29395 net7.n4594 net7.n4593 0.034
R29396 net7.n4602 net7.n4601 0.034
R29397 net7.n4878 net7.n4875 0.034
R29398 net7.n4898 net7.n4897 0.034
R29399 net7.n4798 net7.n4797 0.034
R29400 net7.n4805 net7.n4804 0.034
R29401 net7.n4850 net7.n4849 0.034
R29402 net7.n4860 net7.n4859 0.034
R29403 net7.n4956 net7.n4955 0.034
R29404 net7.n4964 net7.n4963 0.034
R29405 net7.n5240 net7.n5237 0.034
R29406 net7.n5260 net7.n5259 0.034
R29407 net7.n5160 net7.n5159 0.034
R29408 net7.n5167 net7.n5166 0.034
R29409 net7.n5212 net7.n5211 0.034
R29410 net7.n5222 net7.n5221 0.034
R29411 net7.n5318 net7.n5317 0.034
R29412 net7.n5326 net7.n5325 0.034
R29413 net7.n5602 net7.n5599 0.034
R29414 net7.n5622 net7.n5621 0.034
R29415 net7.n5522 net7.n5521 0.034
R29416 net7.n5529 net7.n5528 0.034
R29417 net7.n5574 net7.n5573 0.034
R29418 net7.n5584 net7.n5583 0.034
R29419 net7.n5680 net7.n5679 0.034
R29420 net7.n5688 net7.n5687 0.034
R29421 net7.n5964 net7.n5961 0.034
R29422 net7.n5984 net7.n5983 0.034
R29423 net7.n5884 net7.n5883 0.034
R29424 net7.n5891 net7.n5890 0.034
R29425 net7.n5936 net7.n5935 0.034
R29426 net7.n5946 net7.n5945 0.034
R29427 net7.n6042 net7.n6041 0.034
R29428 net7.n6050 net7.n6049 0.034
R29429 net7.n6326 net7.n6323 0.034
R29430 net7.n6346 net7.n6345 0.034
R29431 net7.n6246 net7.n6245 0.034
R29432 net7.n6253 net7.n6252 0.034
R29433 net7.n6298 net7.n6297 0.034
R29434 net7.n6308 net7.n6307 0.034
R29435 net7.n6404 net7.n6403 0.034
R29436 net7.n6412 net7.n6411 0.034
R29437 net7.n6688 net7.n6685 0.034
R29438 net7.n6708 net7.n6707 0.034
R29439 net7.n6608 net7.n6607 0.034
R29440 net7.n6615 net7.n6614 0.034
R29441 net7.n6660 net7.n6659 0.034
R29442 net7.n6670 net7.n6669 0.034
R29443 net7.n6766 net7.n6765 0.034
R29444 net7.n6774 net7.n6773 0.034
R29445 net7.n7050 net7.n7047 0.034
R29446 net7.n7070 net7.n7069 0.034
R29447 net7.n6970 net7.n6969 0.034
R29448 net7.n6977 net7.n6976 0.034
R29449 net7.n7022 net7.n7021 0.034
R29450 net7.n7032 net7.n7031 0.034
R29451 net7.n7128 net7.n7127 0.034
R29452 net7.n7136 net7.n7135 0.034
R29453 net7.n3605 net7.n3604 0.032
R29454 net7.n3412 net7.n3409 0.032
R29455 net7.n3305 net7.n3304 0.032
R29456 net7.n3443 net7.n3442 0.032
R29457 net7.n3243 net7.n3242 0.032
R29458 net7.n3050 net7.n3047 0.032
R29459 net7.n2943 net7.n2942 0.032
R29460 net7.n3081 net7.n3080 0.032
R29461 net7.n2881 net7.n2880 0.032
R29462 net7.n2688 net7.n2685 0.032
R29463 net7.n2581 net7.n2580 0.032
R29464 net7.n2719 net7.n2718 0.032
R29465 net7.n2519 net7.n2518 0.032
R29466 net7.n2326 net7.n2323 0.032
R29467 net7.n2219 net7.n2218 0.032
R29468 net7.n2357 net7.n2356 0.032
R29469 net7.n2157 net7.n2156 0.032
R29470 net7.n1964 net7.n1961 0.032
R29471 net7.n1857 net7.n1856 0.032
R29472 net7.n1995 net7.n1994 0.032
R29473 net7.n1795 net7.n1794 0.032
R29474 net7.n1602 net7.n1599 0.032
R29475 net7.n1495 net7.n1494 0.032
R29476 net7.n1633 net7.n1632 0.032
R29477 net7.n1433 net7.n1432 0.032
R29478 net7.n1240 net7.n1237 0.032
R29479 net7.n1133 net7.n1132 0.032
R29480 net7.n1271 net7.n1270 0.032
R29481 net7.n1071 net7.n1070 0.032
R29482 net7.n878 net7.n875 0.032
R29483 net7.n771 net7.n770 0.032
R29484 net7.n909 net7.n908 0.032
R29485 net7.n709 net7.n708 0.032
R29486 net7.n516 net7.n513 0.032
R29487 net7.n409 net7.n408 0.032
R29488 net7.n547 net7.n546 0.032
R29489 net7.n348 net7.n347 0.032
R29490 net7.n155 net7.n152 0.032
R29491 net7.n48 net7.n47 0.032
R29492 net7.n186 net7.n185 0.032
R29493 net7.n3689 net7.n3688 0.032
R29494 net7.n3836 net7.n3833 0.032
R29495 net7.n3972 net7.n3971 0.032
R29496 net7.n3757 net7.n3756 0.032
R29497 net7.n4050 net7.n4049 0.032
R29498 net7.n4197 net7.n4194 0.032
R29499 net7.n4333 net7.n4332 0.032
R29500 net7.n4118 net7.n4117 0.032
R29501 net7.n4412 net7.n4411 0.032
R29502 net7.n4559 net7.n4556 0.032
R29503 net7.n4695 net7.n4694 0.032
R29504 net7.n4480 net7.n4479 0.032
R29505 net7.n4774 net7.n4773 0.032
R29506 net7.n4921 net7.n4918 0.032
R29507 net7.n5057 net7.n5056 0.032
R29508 net7.n4842 net7.n4841 0.032
R29509 net7.n5136 net7.n5135 0.032
R29510 net7.n5283 net7.n5280 0.032
R29511 net7.n5419 net7.n5418 0.032
R29512 net7.n5204 net7.n5203 0.032
R29513 net7.n5498 net7.n5497 0.032
R29514 net7.n5645 net7.n5642 0.032
R29515 net7.n5781 net7.n5780 0.032
R29516 net7.n5566 net7.n5565 0.032
R29517 net7.n5860 net7.n5859 0.032
R29518 net7.n6007 net7.n6004 0.032
R29519 net7.n6143 net7.n6142 0.032
R29520 net7.n5928 net7.n5927 0.032
R29521 net7.n6222 net7.n6221 0.032
R29522 net7.n6369 net7.n6366 0.032
R29523 net7.n6505 net7.n6504 0.032
R29524 net7.n6290 net7.n6289 0.032
R29525 net7.n6584 net7.n6583 0.032
R29526 net7.n6731 net7.n6728 0.032
R29527 net7.n6867 net7.n6866 0.032
R29528 net7.n6652 net7.n6651 0.032
R29529 net7.n6946 net7.n6945 0.032
R29530 net7.n7093 net7.n7090 0.032
R29531 net7.n7229 net7.n7228 0.032
R29532 net7.n7014 net7.n7013 0.032
R29533 net7.n3508 net7.n3507 0.031
R29534 net7.n3489 net7.n3485 0.031
R29535 net7.n3466 net7.n3465 0.031
R29536 net7.n3447 net7.n3441 0.031
R29537 net7.n3422 net7.n3421 0.031
R29538 net7.n3358 net7.n3352 0.031
R29539 net7.n3327 net7.n3326 0.031
R29540 net7.n3312 net7.n3311 0.031
R29541 net7.n3146 net7.n3145 0.031
R29542 net7.n3127 net7.n3123 0.031
R29543 net7.n3104 net7.n3103 0.031
R29544 net7.n3085 net7.n3079 0.031
R29545 net7.n3060 net7.n3059 0.031
R29546 net7.n2996 net7.n2990 0.031
R29547 net7.n2965 net7.n2964 0.031
R29548 net7.n2950 net7.n2949 0.031
R29549 net7.n2784 net7.n2783 0.031
R29550 net7.n2765 net7.n2761 0.031
R29551 net7.n2742 net7.n2741 0.031
R29552 net7.n2723 net7.n2717 0.031
R29553 net7.n2698 net7.n2697 0.031
R29554 net7.n2634 net7.n2628 0.031
R29555 net7.n2603 net7.n2602 0.031
R29556 net7.n2588 net7.n2587 0.031
R29557 net7.n2422 net7.n2421 0.031
R29558 net7.n2403 net7.n2399 0.031
R29559 net7.n2380 net7.n2379 0.031
R29560 net7.n2361 net7.n2355 0.031
R29561 net7.n2336 net7.n2335 0.031
R29562 net7.n2272 net7.n2266 0.031
R29563 net7.n2241 net7.n2240 0.031
R29564 net7.n2226 net7.n2225 0.031
R29565 net7.n2060 net7.n2059 0.031
R29566 net7.n2041 net7.n2037 0.031
R29567 net7.n2018 net7.n2017 0.031
R29568 net7.n1999 net7.n1993 0.031
R29569 net7.n1974 net7.n1973 0.031
R29570 net7.n1910 net7.n1904 0.031
R29571 net7.n1879 net7.n1878 0.031
R29572 net7.n1864 net7.n1863 0.031
R29573 net7.n1698 net7.n1697 0.031
R29574 net7.n1679 net7.n1675 0.031
R29575 net7.n1656 net7.n1655 0.031
R29576 net7.n1637 net7.n1631 0.031
R29577 net7.n1612 net7.n1611 0.031
R29578 net7.n1548 net7.n1542 0.031
R29579 net7.n1517 net7.n1516 0.031
R29580 net7.n1502 net7.n1501 0.031
R29581 net7.n1336 net7.n1335 0.031
R29582 net7.n1317 net7.n1313 0.031
R29583 net7.n1294 net7.n1293 0.031
R29584 net7.n1275 net7.n1269 0.031
R29585 net7.n1250 net7.n1249 0.031
R29586 net7.n1186 net7.n1180 0.031
R29587 net7.n1155 net7.n1154 0.031
R29588 net7.n1140 net7.n1139 0.031
R29589 net7.n974 net7.n973 0.031
R29590 net7.n955 net7.n951 0.031
R29591 net7.n932 net7.n931 0.031
R29592 net7.n913 net7.n907 0.031
R29593 net7.n888 net7.n887 0.031
R29594 net7.n824 net7.n818 0.031
R29595 net7.n793 net7.n792 0.031
R29596 net7.n778 net7.n777 0.031
R29597 net7.n612 net7.n611 0.031
R29598 net7.n593 net7.n589 0.031
R29599 net7.n570 net7.n569 0.031
R29600 net7.n551 net7.n545 0.031
R29601 net7.n526 net7.n525 0.031
R29602 net7.n462 net7.n456 0.031
R29603 net7.n431 net7.n430 0.031
R29604 net7.n416 net7.n415 0.031
R29605 net7.n251 net7.n250 0.031
R29606 net7.n232 net7.n228 0.031
R29607 net7.n209 net7.n208 0.031
R29608 net7.n190 net7.n184 0.031
R29609 net7.n165 net7.n164 0.031
R29610 net7.n101 net7.n95 0.031
R29611 net7.n70 net7.n69 0.031
R29612 net7.n55 net7.n54 0.031
R29613 net7.n3696 net7.n3695 0.031
R29614 net7.n3710 net7.n3709 0.031
R29615 net7.n3734 net7.n3728 0.031
R29616 net7.n3753 net7.n3752 0.031
R29617 net7.n3841 net7.n3773 0.031
R29618 net7.n3860 net7.n3859 0.031
R29619 net7.n3883 net7.n3877 0.031
R29620 net7.n3903 net7.n3902 0.031
R29621 net7.n4057 net7.n4056 0.031
R29622 net7.n4071 net7.n4070 0.031
R29623 net7.n4095 net7.n4089 0.031
R29624 net7.n4114 net7.n4113 0.031
R29625 net7.n4202 net7.n4134 0.031
R29626 net7.n4221 net7.n4220 0.031
R29627 net7.n4244 net7.n4238 0.031
R29628 net7.n4264 net7.n4263 0.031
R29629 net7.n4419 net7.n4418 0.031
R29630 net7.n4433 net7.n4432 0.031
R29631 net7.n4457 net7.n4451 0.031
R29632 net7.n4476 net7.n4475 0.031
R29633 net7.n4564 net7.n4496 0.031
R29634 net7.n4583 net7.n4582 0.031
R29635 net7.n4606 net7.n4600 0.031
R29636 net7.n4626 net7.n4625 0.031
R29637 net7.n4781 net7.n4780 0.031
R29638 net7.n4795 net7.n4794 0.031
R29639 net7.n4819 net7.n4813 0.031
R29640 net7.n4838 net7.n4837 0.031
R29641 net7.n4926 net7.n4858 0.031
R29642 net7.n4945 net7.n4944 0.031
R29643 net7.n4968 net7.n4962 0.031
R29644 net7.n4988 net7.n4987 0.031
R29645 net7.n5143 net7.n5142 0.031
R29646 net7.n5157 net7.n5156 0.031
R29647 net7.n5181 net7.n5175 0.031
R29648 net7.n5200 net7.n5199 0.031
R29649 net7.n5288 net7.n5220 0.031
R29650 net7.n5307 net7.n5306 0.031
R29651 net7.n5330 net7.n5324 0.031
R29652 net7.n5350 net7.n5349 0.031
R29653 net7.n5505 net7.n5504 0.031
R29654 net7.n5519 net7.n5518 0.031
R29655 net7.n5543 net7.n5537 0.031
R29656 net7.n5562 net7.n5561 0.031
R29657 net7.n5650 net7.n5582 0.031
R29658 net7.n5669 net7.n5668 0.031
R29659 net7.n5692 net7.n5686 0.031
R29660 net7.n5712 net7.n5711 0.031
R29661 net7.n5867 net7.n5866 0.031
R29662 net7.n5881 net7.n5880 0.031
R29663 net7.n5905 net7.n5899 0.031
R29664 net7.n5924 net7.n5923 0.031
R29665 net7.n6012 net7.n5944 0.031
R29666 net7.n6031 net7.n6030 0.031
R29667 net7.n6054 net7.n6048 0.031
R29668 net7.n6074 net7.n6073 0.031
R29669 net7.n6229 net7.n6228 0.031
R29670 net7.n6243 net7.n6242 0.031
R29671 net7.n6267 net7.n6261 0.031
R29672 net7.n6286 net7.n6285 0.031
R29673 net7.n6374 net7.n6306 0.031
R29674 net7.n6393 net7.n6392 0.031
R29675 net7.n6416 net7.n6410 0.031
R29676 net7.n6436 net7.n6435 0.031
R29677 net7.n6591 net7.n6590 0.031
R29678 net7.n6605 net7.n6604 0.031
R29679 net7.n6629 net7.n6623 0.031
R29680 net7.n6648 net7.n6647 0.031
R29681 net7.n6736 net7.n6668 0.031
R29682 net7.n6755 net7.n6754 0.031
R29683 net7.n6778 net7.n6772 0.031
R29684 net7.n6798 net7.n6797 0.031
R29685 net7.n6953 net7.n6952 0.031
R29686 net7.n6967 net7.n6966 0.031
R29687 net7.n6991 net7.n6985 0.031
R29688 net7.n7010 net7.n7009 0.031
R29689 net7.n7098 net7.n7030 0.031
R29690 net7.n7117 net7.n7116 0.031
R29691 net7.n7140 net7.n7134 0.031
R29692 net7.n7160 net7.n7159 0.031
R29693 net7.n3584 net7.n3580 0.03
R29694 net7.n3528 net7.n3525 0.03
R29695 net7.n3383 net7.n3380 0.03
R29696 net7.n3278 net7.n3277 0.03
R29697 net7.n3295 net7.n3294 0.03
R29698 net7.n3427 net7.n3426 0.03
R29699 net7.n3222 net7.n3218 0.03
R29700 net7.n3166 net7.n3163 0.03
R29701 net7.n3021 net7.n3018 0.03
R29702 net7.n2916 net7.n2915 0.03
R29703 net7.n2933 net7.n2932 0.03
R29704 net7.n3065 net7.n3064 0.03
R29705 net7.n2860 net7.n2856 0.03
R29706 net7.n2804 net7.n2801 0.03
R29707 net7.n2659 net7.n2656 0.03
R29708 net7.n2554 net7.n2553 0.03
R29709 net7.n2571 net7.n2570 0.03
R29710 net7.n2703 net7.n2702 0.03
R29711 net7.n2498 net7.n2494 0.03
R29712 net7.n2442 net7.n2439 0.03
R29713 net7.n2297 net7.n2294 0.03
R29714 net7.n2192 net7.n2191 0.03
R29715 net7.n2209 net7.n2208 0.03
R29716 net7.n2341 net7.n2340 0.03
R29717 net7.n2136 net7.n2132 0.03
R29718 net7.n2080 net7.n2077 0.03
R29719 net7.n1935 net7.n1932 0.03
R29720 net7.n1830 net7.n1829 0.03
R29721 net7.n1847 net7.n1846 0.03
R29722 net7.n1979 net7.n1978 0.03
R29723 net7.n1774 net7.n1770 0.03
R29724 net7.n1718 net7.n1715 0.03
R29725 net7.n1573 net7.n1570 0.03
R29726 net7.n1468 net7.n1467 0.03
R29727 net7.n1485 net7.n1484 0.03
R29728 net7.n1617 net7.n1616 0.03
R29729 net7.n1412 net7.n1408 0.03
R29730 net7.n1356 net7.n1353 0.03
R29731 net7.n1211 net7.n1208 0.03
R29732 net7.n1106 net7.n1105 0.03
R29733 net7.n1123 net7.n1122 0.03
R29734 net7.n1255 net7.n1254 0.03
R29735 net7.n1050 net7.n1046 0.03
R29736 net7.n994 net7.n991 0.03
R29737 net7.n849 net7.n846 0.03
R29738 net7.n744 net7.n743 0.03
R29739 net7.n761 net7.n760 0.03
R29740 net7.n893 net7.n892 0.03
R29741 net7.n688 net7.n684 0.03
R29742 net7.n632 net7.n629 0.03
R29743 net7.n487 net7.n484 0.03
R29744 net7.n382 net7.n381 0.03
R29745 net7.n399 net7.n398 0.03
R29746 net7.n531 net7.n530 0.03
R29747 net7.n327 net7.n323 0.03
R29748 net7.n271 net7.n268 0.03
R29749 net7.n126 net7.n123 0.03
R29750 net7.n21 net7.n20 0.03
R29751 net7.n38 net7.n37 0.03
R29752 net7.n170 net7.n169 0.03
R29753 net7.n3670 net7.n3669 0.03
R29754 net7.n3809 net7.n3806 0.03
R29755 net7.n3822 net7.n3819 0.03
R29756 net7.n3945 net7.n3944 0.03
R29757 net7.n3962 net7.n3961 0.03
R29758 net7.n3768 net7.n3767 0.03
R29759 net7.n3892 net7.n3891 0.03
R29760 net7.n4031 net7.n4030 0.03
R29761 net7.n4170 net7.n4167 0.03
R29762 net7.n4183 net7.n4180 0.03
R29763 net7.n4306 net7.n4305 0.03
R29764 net7.n4323 net7.n4322 0.03
R29765 net7.n4129 net7.n4128 0.03
R29766 net7.n4253 net7.n4252 0.03
R29767 net7.n4393 net7.n4392 0.03
R29768 net7.n4532 net7.n4529 0.03
R29769 net7.n4545 net7.n4542 0.03
R29770 net7.n4668 net7.n4667 0.03
R29771 net7.n4685 net7.n4684 0.03
R29772 net7.n4491 net7.n4490 0.03
R29773 net7.n4615 net7.n4614 0.03
R29774 net7.n4755 net7.n4754 0.03
R29775 net7.n4894 net7.n4891 0.03
R29776 net7.n4907 net7.n4904 0.03
R29777 net7.n5030 net7.n5029 0.03
R29778 net7.n5047 net7.n5046 0.03
R29779 net7.n4853 net7.n4852 0.03
R29780 net7.n4977 net7.n4976 0.03
R29781 net7.n5117 net7.n5116 0.03
R29782 net7.n5256 net7.n5253 0.03
R29783 net7.n5269 net7.n5266 0.03
R29784 net7.n5392 net7.n5391 0.03
R29785 net7.n5409 net7.n5408 0.03
R29786 net7.n5215 net7.n5214 0.03
R29787 net7.n5339 net7.n5338 0.03
R29788 net7.n5479 net7.n5478 0.03
R29789 net7.n5618 net7.n5615 0.03
R29790 net7.n5631 net7.n5628 0.03
R29791 net7.n5754 net7.n5753 0.03
R29792 net7.n5771 net7.n5770 0.03
R29793 net7.n5577 net7.n5576 0.03
R29794 net7.n5701 net7.n5700 0.03
R29795 net7.n5841 net7.n5840 0.03
R29796 net7.n5980 net7.n5977 0.03
R29797 net7.n5993 net7.n5990 0.03
R29798 net7.n6116 net7.n6115 0.03
R29799 net7.n6133 net7.n6132 0.03
R29800 net7.n5939 net7.n5938 0.03
R29801 net7.n6063 net7.n6062 0.03
R29802 net7.n6203 net7.n6202 0.03
R29803 net7.n6342 net7.n6339 0.03
R29804 net7.n6355 net7.n6352 0.03
R29805 net7.n6478 net7.n6477 0.03
R29806 net7.n6495 net7.n6494 0.03
R29807 net7.n6301 net7.n6300 0.03
R29808 net7.n6425 net7.n6424 0.03
R29809 net7.n6565 net7.n6564 0.03
R29810 net7.n6704 net7.n6701 0.03
R29811 net7.n6717 net7.n6714 0.03
R29812 net7.n6840 net7.n6839 0.03
R29813 net7.n6857 net7.n6856 0.03
R29814 net7.n6663 net7.n6662 0.03
R29815 net7.n6787 net7.n6786 0.03
R29816 net7.n6927 net7.n6926 0.03
R29817 net7.n7066 net7.n7063 0.03
R29818 net7.n7079 net7.n7076 0.03
R29819 net7.n7202 net7.n7201 0.03
R29820 net7.n7219 net7.n7218 0.03
R29821 net7.n7025 net7.n7024 0.03
R29822 net7.n7149 net7.n7148 0.03
R29823 net7.n3694 net7.n3628 0.029
R29824 net7.n4055 net7.n3989 0.029
R29825 net7.n4417 net7.n4351 0.029
R29826 net7.n4779 net7.n4713 0.029
R29827 net7.n5141 net7.n5075 0.029
R29828 net7.n5503 net7.n5437 0.029
R29829 net7.n5865 net7.n5799 0.029
R29830 net7.n6227 net7.n6161 0.029
R29831 net7.n6589 net7.n6523 0.029
R29832 net7.n6951 net7.n6885 0.029
R29833 net7.n3595 net7.n3594 0.028
R29834 net7.n3538 net7.n3536 0.028
R29835 net7.n3417 net7.n3414 0.028
R29836 net7.n3407 net7.n3406 0.028
R29837 net7.n3498 net7.n3497 0.028
R29838 net7.n3473 net7.n3472 0.028
R29839 net7.n3471 net7.n3470 0.028
R29840 net7.n3432 net7.n3431 0.028
R29841 net7.n3233 net7.n3232 0.028
R29842 net7.n3176 net7.n3174 0.028
R29843 net7.n3055 net7.n3052 0.028
R29844 net7.n3045 net7.n3044 0.028
R29845 net7.n3136 net7.n3135 0.028
R29846 net7.n3111 net7.n3110 0.028
R29847 net7.n3109 net7.n3108 0.028
R29848 net7.n3070 net7.n3069 0.028
R29849 net7.n2871 net7.n2870 0.028
R29850 net7.n2814 net7.n2812 0.028
R29851 net7.n2693 net7.n2690 0.028
R29852 net7.n2683 net7.n2682 0.028
R29853 net7.n2774 net7.n2773 0.028
R29854 net7.n2749 net7.n2748 0.028
R29855 net7.n2747 net7.n2746 0.028
R29856 net7.n2708 net7.n2707 0.028
R29857 net7.n2509 net7.n2508 0.028
R29858 net7.n2452 net7.n2450 0.028
R29859 net7.n2331 net7.n2328 0.028
R29860 net7.n2321 net7.n2320 0.028
R29861 net7.n2412 net7.n2411 0.028
R29862 net7.n2387 net7.n2386 0.028
R29863 net7.n2385 net7.n2384 0.028
R29864 net7.n2346 net7.n2345 0.028
R29865 net7.n2147 net7.n2146 0.028
R29866 net7.n2090 net7.n2088 0.028
R29867 net7.n1969 net7.n1966 0.028
R29868 net7.n1959 net7.n1958 0.028
R29869 net7.n2050 net7.n2049 0.028
R29870 net7.n2025 net7.n2024 0.028
R29871 net7.n2023 net7.n2022 0.028
R29872 net7.n1984 net7.n1983 0.028
R29873 net7.n1785 net7.n1784 0.028
R29874 net7.n1728 net7.n1726 0.028
R29875 net7.n1607 net7.n1604 0.028
R29876 net7.n1597 net7.n1596 0.028
R29877 net7.n1688 net7.n1687 0.028
R29878 net7.n1663 net7.n1662 0.028
R29879 net7.n1661 net7.n1660 0.028
R29880 net7.n1622 net7.n1621 0.028
R29881 net7.n1423 net7.n1422 0.028
R29882 net7.n1366 net7.n1364 0.028
R29883 net7.n1245 net7.n1242 0.028
R29884 net7.n1235 net7.n1234 0.028
R29885 net7.n1326 net7.n1325 0.028
R29886 net7.n1301 net7.n1300 0.028
R29887 net7.n1299 net7.n1298 0.028
R29888 net7.n1260 net7.n1259 0.028
R29889 net7.n1061 net7.n1060 0.028
R29890 net7.n1004 net7.n1002 0.028
R29891 net7.n883 net7.n880 0.028
R29892 net7.n873 net7.n872 0.028
R29893 net7.n964 net7.n963 0.028
R29894 net7.n939 net7.n938 0.028
R29895 net7.n937 net7.n936 0.028
R29896 net7.n898 net7.n897 0.028
R29897 net7.n699 net7.n698 0.028
R29898 net7.n642 net7.n640 0.028
R29899 net7.n521 net7.n518 0.028
R29900 net7.n511 net7.n510 0.028
R29901 net7.n602 net7.n601 0.028
R29902 net7.n577 net7.n576 0.028
R29903 net7.n575 net7.n574 0.028
R29904 net7.n536 net7.n535 0.028
R29905 net7.n338 net7.n337 0.028
R29906 net7.n281 net7.n279 0.028
R29907 net7.n160 net7.n157 0.028
R29908 net7.n150 net7.n149 0.028
R29909 net7.n241 net7.n240 0.028
R29910 net7.n216 net7.n215 0.028
R29911 net7.n214 net7.n213 0.028
R29912 net7.n175 net7.n174 0.028
R29913 net7.n3681 net7.n3680 0.028
R29914 net7.n3796 net7.n3795 0.028
R29915 net7.n3839 net7.n3838 0.028
R29916 net7.n3831 net7.n3830 0.028
R29917 net7.n3724 net7.n3723 0.028
R29918 net7.n3730 net7.n3729 0.028
R29919 net7.n3759 net7.n3758 0.028
R29920 net7.n3850 net7.n3849 0.028
R29921 net7.n4042 net7.n4041 0.028
R29922 net7.n4157 net7.n4156 0.028
R29923 net7.n4200 net7.n4199 0.028
R29924 net7.n4192 net7.n4191 0.028
R29925 net7.n4085 net7.n4084 0.028
R29926 net7.n4091 net7.n4090 0.028
R29927 net7.n4120 net7.n4119 0.028
R29928 net7.n4211 net7.n4210 0.028
R29929 net7.n4404 net7.n4403 0.028
R29930 net7.n4519 net7.n4518 0.028
R29931 net7.n4562 net7.n4561 0.028
R29932 net7.n4554 net7.n4553 0.028
R29933 net7.n4447 net7.n4446 0.028
R29934 net7.n4453 net7.n4452 0.028
R29935 net7.n4482 net7.n4481 0.028
R29936 net7.n4573 net7.n4572 0.028
R29937 net7.n4766 net7.n4765 0.028
R29938 net7.n4881 net7.n4880 0.028
R29939 net7.n4924 net7.n4923 0.028
R29940 net7.n4916 net7.n4915 0.028
R29941 net7.n4809 net7.n4808 0.028
R29942 net7.n4815 net7.n4814 0.028
R29943 net7.n4844 net7.n4843 0.028
R29944 net7.n4935 net7.n4934 0.028
R29945 net7.n5128 net7.n5127 0.028
R29946 net7.n5243 net7.n5242 0.028
R29947 net7.n5286 net7.n5285 0.028
R29948 net7.n5278 net7.n5277 0.028
R29949 net7.n5171 net7.n5170 0.028
R29950 net7.n5177 net7.n5176 0.028
R29951 net7.n5206 net7.n5205 0.028
R29952 net7.n5297 net7.n5296 0.028
R29953 net7.n5490 net7.n5489 0.028
R29954 net7.n5605 net7.n5604 0.028
R29955 net7.n5648 net7.n5647 0.028
R29956 net7.n5640 net7.n5639 0.028
R29957 net7.n5533 net7.n5532 0.028
R29958 net7.n5539 net7.n5538 0.028
R29959 net7.n5568 net7.n5567 0.028
R29960 net7.n5659 net7.n5658 0.028
R29961 net7.n5852 net7.n5851 0.028
R29962 net7.n5967 net7.n5966 0.028
R29963 net7.n6010 net7.n6009 0.028
R29964 net7.n6002 net7.n6001 0.028
R29965 net7.n5895 net7.n5894 0.028
R29966 net7.n5901 net7.n5900 0.028
R29967 net7.n5930 net7.n5929 0.028
R29968 net7.n6021 net7.n6020 0.028
R29969 net7.n6214 net7.n6213 0.028
R29970 net7.n6329 net7.n6328 0.028
R29971 net7.n6372 net7.n6371 0.028
R29972 net7.n6364 net7.n6363 0.028
R29973 net7.n6257 net7.n6256 0.028
R29974 net7.n6263 net7.n6262 0.028
R29975 net7.n6292 net7.n6291 0.028
R29976 net7.n6383 net7.n6382 0.028
R29977 net7.n6576 net7.n6575 0.028
R29978 net7.n6691 net7.n6690 0.028
R29979 net7.n6734 net7.n6733 0.028
R29980 net7.n6726 net7.n6725 0.028
R29981 net7.n6619 net7.n6618 0.028
R29982 net7.n6625 net7.n6624 0.028
R29983 net7.n6654 net7.n6653 0.028
R29984 net7.n6745 net7.n6744 0.028
R29985 net7.n6938 net7.n6937 0.028
R29986 net7.n7053 net7.n7052 0.028
R29987 net7.n7096 net7.n7095 0.028
R29988 net7.n7088 net7.n7087 0.028
R29989 net7.n6981 net7.n6980 0.028
R29990 net7.n6987 net7.n6986 0.028
R29991 net7.n7016 net7.n7015 0.028
R29992 net7.n7107 net7.n7106 0.028
R29993 net7.n3310 net7.n3267 0.027
R29994 net7.n2948 net7.n2905 0.027
R29995 net7.n2586 net7.n2543 0.027
R29996 net7.n2224 net7.n2181 0.027
R29997 net7.n1862 net7.n1819 0.027
R29998 net7.n1500 net7.n1457 0.027
R29999 net7.n1138 net7.n1095 0.027
R30000 net7.n776 net7.n733 0.027
R30001 net7.n414 net7.n371 0.027
R30002 net7.n53 net7.n10 0.027
R30003 net7.n3500 net7.n3496 0.027
R30004 net7.n3458 net7.n3454 0.027
R30005 net7.n3369 net7.n3365 0.027
R30006 net7.n3319 net7.n3315 0.027
R30007 net7.n3138 net7.n3134 0.027
R30008 net7.n3096 net7.n3092 0.027
R30009 net7.n3007 net7.n3003 0.027
R30010 net7.n2957 net7.n2953 0.027
R30011 net7.n2776 net7.n2772 0.027
R30012 net7.n2734 net7.n2730 0.027
R30013 net7.n2645 net7.n2641 0.027
R30014 net7.n2595 net7.n2591 0.027
R30015 net7.n2414 net7.n2410 0.027
R30016 net7.n2372 net7.n2368 0.027
R30017 net7.n2283 net7.n2279 0.027
R30018 net7.n2233 net7.n2229 0.027
R30019 net7.n2052 net7.n2048 0.027
R30020 net7.n2010 net7.n2006 0.027
R30021 net7.n1921 net7.n1917 0.027
R30022 net7.n1871 net7.n1867 0.027
R30023 net7.n1690 net7.n1686 0.027
R30024 net7.n1648 net7.n1644 0.027
R30025 net7.n1559 net7.n1555 0.027
R30026 net7.n1509 net7.n1505 0.027
R30027 net7.n1328 net7.n1324 0.027
R30028 net7.n1286 net7.n1282 0.027
R30029 net7.n1197 net7.n1193 0.027
R30030 net7.n1147 net7.n1143 0.027
R30031 net7.n966 net7.n962 0.027
R30032 net7.n924 net7.n920 0.027
R30033 net7.n835 net7.n831 0.027
R30034 net7.n785 net7.n781 0.027
R30035 net7.n604 net7.n600 0.027
R30036 net7.n562 net7.n558 0.027
R30037 net7.n473 net7.n469 0.027
R30038 net7.n423 net7.n419 0.027
R30039 net7.n243 net7.n239 0.027
R30040 net7.n201 net7.n197 0.027
R30041 net7.n112 net7.n108 0.027
R30042 net7.n62 net7.n58 0.027
R30043 net7.n3703 net7.n3699 0.027
R30044 net7.n3745 net7.n3741 0.027
R30045 net7.n3852 net7.n3848 0.027
R30046 net7.n3894 net7.n3890 0.027
R30047 net7.n4064 net7.n4060 0.027
R30048 net7.n4106 net7.n4102 0.027
R30049 net7.n4213 net7.n4209 0.027
R30050 net7.n4255 net7.n4251 0.027
R30051 net7.n4426 net7.n4422 0.027
R30052 net7.n4468 net7.n4464 0.027
R30053 net7.n4575 net7.n4571 0.027
R30054 net7.n4617 net7.n4613 0.027
R30055 net7.n4788 net7.n4784 0.027
R30056 net7.n4830 net7.n4826 0.027
R30057 net7.n4937 net7.n4933 0.027
R30058 net7.n4979 net7.n4975 0.027
R30059 net7.n5150 net7.n5146 0.027
R30060 net7.n5192 net7.n5188 0.027
R30061 net7.n5299 net7.n5295 0.027
R30062 net7.n5341 net7.n5337 0.027
R30063 net7.n5512 net7.n5508 0.027
R30064 net7.n5554 net7.n5550 0.027
R30065 net7.n5661 net7.n5657 0.027
R30066 net7.n5703 net7.n5699 0.027
R30067 net7.n5874 net7.n5870 0.027
R30068 net7.n5916 net7.n5912 0.027
R30069 net7.n6023 net7.n6019 0.027
R30070 net7.n6065 net7.n6061 0.027
R30071 net7.n6236 net7.n6232 0.027
R30072 net7.n6278 net7.n6274 0.027
R30073 net7.n6385 net7.n6381 0.027
R30074 net7.n6427 net7.n6423 0.027
R30075 net7.n6598 net7.n6594 0.027
R30076 net7.n6640 net7.n6636 0.027
R30077 net7.n6747 net7.n6743 0.027
R30078 net7.n6789 net7.n6785 0.027
R30079 net7.n6960 net7.n6956 0.027
R30080 net7.n7002 net7.n6998 0.027
R30081 net7.n7109 net7.n7105 0.027
R30082 net7.n7151 net7.n7147 0.027
R30083 net7.n3545 net7.n3544 0.026
R30084 net7.n3613 net7.n3612 0.026
R30085 net7.n3456 net7.n3455 0.026
R30086 net7.n3354 net7.n3353 0.026
R30087 net7.n3337 net7.n3336 0.026
R30088 net7.n3183 net7.n3182 0.026
R30089 net7.n3251 net7.n3250 0.026
R30090 net7.n3094 net7.n3093 0.026
R30091 net7.n2992 net7.n2991 0.026
R30092 net7.n2975 net7.n2974 0.026
R30093 net7.n2821 net7.n2820 0.026
R30094 net7.n2889 net7.n2888 0.026
R30095 net7.n2732 net7.n2731 0.026
R30096 net7.n2630 net7.n2629 0.026
R30097 net7.n2613 net7.n2612 0.026
R30098 net7.n2459 net7.n2458 0.026
R30099 net7.n2527 net7.n2526 0.026
R30100 net7.n2370 net7.n2369 0.026
R30101 net7.n2268 net7.n2267 0.026
R30102 net7.n2251 net7.n2250 0.026
R30103 net7.n2097 net7.n2096 0.026
R30104 net7.n2165 net7.n2164 0.026
R30105 net7.n2008 net7.n2007 0.026
R30106 net7.n1906 net7.n1905 0.026
R30107 net7.n1889 net7.n1888 0.026
R30108 net7.n1735 net7.n1734 0.026
R30109 net7.n1803 net7.n1802 0.026
R30110 net7.n1646 net7.n1645 0.026
R30111 net7.n1544 net7.n1543 0.026
R30112 net7.n1527 net7.n1526 0.026
R30113 net7.n1373 net7.n1372 0.026
R30114 net7.n1441 net7.n1440 0.026
R30115 net7.n1284 net7.n1283 0.026
R30116 net7.n1182 net7.n1181 0.026
R30117 net7.n1165 net7.n1164 0.026
R30118 net7.n1011 net7.n1010 0.026
R30119 net7.n1079 net7.n1078 0.026
R30120 net7.n922 net7.n921 0.026
R30121 net7.n820 net7.n819 0.026
R30122 net7.n803 net7.n802 0.026
R30123 net7.n649 net7.n648 0.026
R30124 net7.n717 net7.n716 0.026
R30125 net7.n560 net7.n559 0.026
R30126 net7.n458 net7.n457 0.026
R30127 net7.n441 net7.n440 0.026
R30128 net7.n288 net7.n287 0.026
R30129 net7.n356 net7.n355 0.026
R30130 net7.n199 net7.n198 0.026
R30131 net7.n97 net7.n96 0.026
R30132 net7.n80 net7.n79 0.026
R30133 net7.n3788 net7.n3787 0.026
R30134 net7.n3627 net7.n3626 0.026
R30135 net7.n3864 net7.n3863 0.026
R30136 net7.n3866 net7.n3865 0.026
R30137 net7.n4149 net7.n4148 0.026
R30138 net7.n3988 net7.n3987 0.026
R30139 net7.n4225 net7.n4224 0.026
R30140 net7.n4227 net7.n4226 0.026
R30141 net7.n4511 net7.n4510 0.026
R30142 net7.n4350 net7.n4349 0.026
R30143 net7.n4587 net7.n4586 0.026
R30144 net7.n4589 net7.n4588 0.026
R30145 net7.n4873 net7.n4872 0.026
R30146 net7.n4712 net7.n4711 0.026
R30147 net7.n4949 net7.n4948 0.026
R30148 net7.n4951 net7.n4950 0.026
R30149 net7.n5235 net7.n5234 0.026
R30150 net7.n5074 net7.n5073 0.026
R30151 net7.n5311 net7.n5310 0.026
R30152 net7.n5313 net7.n5312 0.026
R30153 net7.n5597 net7.n5596 0.026
R30154 net7.n5436 net7.n5435 0.026
R30155 net7.n5673 net7.n5672 0.026
R30156 net7.n5675 net7.n5674 0.026
R30157 net7.n5959 net7.n5958 0.026
R30158 net7.n5798 net7.n5797 0.026
R30159 net7.n6035 net7.n6034 0.026
R30160 net7.n6037 net7.n6036 0.026
R30161 net7.n6321 net7.n6320 0.026
R30162 net7.n6160 net7.n6159 0.026
R30163 net7.n6397 net7.n6396 0.026
R30164 net7.n6399 net7.n6398 0.026
R30165 net7.n6683 net7.n6682 0.026
R30166 net7.n6522 net7.n6521 0.026
R30167 net7.n6759 net7.n6758 0.026
R30168 net7.n6761 net7.n6760 0.026
R30169 net7.n7045 net7.n7044 0.026
R30170 net7.n6884 net7.n6883 0.026
R30171 net7.n7121 net7.n7120 0.026
R30172 net7.n7123 net7.n7122 0.026
R30173 net7.n3405 net7.n3404 0.024
R30174 net7.n3506 net7.n3505 0.024
R30175 net7.n3495 net7.n3494 0.024
R30176 net7.n3464 net7.n3463 0.024
R30177 net7.n3453 net7.n3452 0.024
R30178 net7.n3420 net7.n3419 0.024
R30179 net7.n3364 net7.n3363 0.024
R30180 net7.n3259 net7.n3258 0.024
R30181 net7.n3266 net7.n3265 0.024
R30182 net7.n3043 net7.n3042 0.024
R30183 net7.n3144 net7.n3143 0.024
R30184 net7.n3133 net7.n3132 0.024
R30185 net7.n3102 net7.n3101 0.024
R30186 net7.n3091 net7.n3090 0.024
R30187 net7.n3058 net7.n3057 0.024
R30188 net7.n3002 net7.n3001 0.024
R30189 net7.n2897 net7.n2896 0.024
R30190 net7.n2904 net7.n2903 0.024
R30191 net7.n2681 net7.n2680 0.024
R30192 net7.n2782 net7.n2781 0.024
R30193 net7.n2771 net7.n2770 0.024
R30194 net7.n2740 net7.n2739 0.024
R30195 net7.n2729 net7.n2728 0.024
R30196 net7.n2696 net7.n2695 0.024
R30197 net7.n2640 net7.n2639 0.024
R30198 net7.n2535 net7.n2534 0.024
R30199 net7.n2542 net7.n2541 0.024
R30200 net7.n2319 net7.n2318 0.024
R30201 net7.n2420 net7.n2419 0.024
R30202 net7.n2409 net7.n2408 0.024
R30203 net7.n2378 net7.n2377 0.024
R30204 net7.n2367 net7.n2366 0.024
R30205 net7.n2334 net7.n2333 0.024
R30206 net7.n2278 net7.n2277 0.024
R30207 net7.n2173 net7.n2172 0.024
R30208 net7.n2180 net7.n2179 0.024
R30209 net7.n1957 net7.n1956 0.024
R30210 net7.n2058 net7.n2057 0.024
R30211 net7.n2047 net7.n2046 0.024
R30212 net7.n2016 net7.n2015 0.024
R30213 net7.n2005 net7.n2004 0.024
R30214 net7.n1972 net7.n1971 0.024
R30215 net7.n1916 net7.n1915 0.024
R30216 net7.n1811 net7.n1810 0.024
R30217 net7.n1818 net7.n1817 0.024
R30218 net7.n1595 net7.n1594 0.024
R30219 net7.n1696 net7.n1695 0.024
R30220 net7.n1685 net7.n1684 0.024
R30221 net7.n1654 net7.n1653 0.024
R30222 net7.n1643 net7.n1642 0.024
R30223 net7.n1610 net7.n1609 0.024
R30224 net7.n1554 net7.n1553 0.024
R30225 net7.n1449 net7.n1448 0.024
R30226 net7.n1456 net7.n1455 0.024
R30227 net7.n1233 net7.n1232 0.024
R30228 net7.n1334 net7.n1333 0.024
R30229 net7.n1323 net7.n1322 0.024
R30230 net7.n1292 net7.n1291 0.024
R30231 net7.n1281 net7.n1280 0.024
R30232 net7.n1248 net7.n1247 0.024
R30233 net7.n1192 net7.n1191 0.024
R30234 net7.n1087 net7.n1086 0.024
R30235 net7.n1094 net7.n1093 0.024
R30236 net7.n871 net7.n870 0.024
R30237 net7.n972 net7.n971 0.024
R30238 net7.n961 net7.n960 0.024
R30239 net7.n930 net7.n929 0.024
R30240 net7.n919 net7.n918 0.024
R30241 net7.n886 net7.n885 0.024
R30242 net7.n830 net7.n829 0.024
R30243 net7.n725 net7.n724 0.024
R30244 net7.n732 net7.n731 0.024
R30245 net7.n509 net7.n508 0.024
R30246 net7.n610 net7.n609 0.024
R30247 net7.n599 net7.n598 0.024
R30248 net7.n568 net7.n567 0.024
R30249 net7.n557 net7.n556 0.024
R30250 net7.n524 net7.n523 0.024
R30251 net7.n468 net7.n467 0.024
R30252 net7.n363 net7.n362 0.024
R30253 net7.n370 net7.n369 0.024
R30254 net7.n148 net7.n147 0.024
R30255 net7.n249 net7.n248 0.024
R30256 net7.n238 net7.n237 0.024
R30257 net7.n207 net7.n206 0.024
R30258 net7.n196 net7.n195 0.024
R30259 net7.n163 net7.n162 0.024
R30260 net7.n107 net7.n106 0.024
R30261 net7.n2 net7.n1 0.024
R30262 net7.n9 net7.n8 0.024
R30263 net7.n3623 net7.n3622 0.024
R30264 net7.n3621 net7.n3620 0.024
R30265 net7.n3708 net7.n3707 0.024
R30266 net7.n3740 net7.n3738 0.024
R30267 net7.n3751 net7.n3749 0.024
R30268 net7.n3847 net7.n3845 0.024
R30269 net7.n3858 net7.n3856 0.024
R30270 net7.n3889 net7.n3887 0.024
R30271 net7.n3907 net7.n3906 0.024
R30272 net7.n3984 net7.n3983 0.024
R30273 net7.n3982 net7.n3981 0.024
R30274 net7.n4069 net7.n4068 0.024
R30275 net7.n4101 net7.n4099 0.024
R30276 net7.n4112 net7.n4110 0.024
R30277 net7.n4208 net7.n4206 0.024
R30278 net7.n4219 net7.n4217 0.024
R30279 net7.n4250 net7.n4248 0.024
R30280 net7.n4268 net7.n4267 0.024
R30281 net7.n4346 net7.n4345 0.024
R30282 net7.n4344 net7.n4343 0.024
R30283 net7.n4431 net7.n4430 0.024
R30284 net7.n4463 net7.n4461 0.024
R30285 net7.n4474 net7.n4472 0.024
R30286 net7.n4570 net7.n4568 0.024
R30287 net7.n4581 net7.n4579 0.024
R30288 net7.n4612 net7.n4610 0.024
R30289 net7.n4630 net7.n4629 0.024
R30290 net7.n4708 net7.n4707 0.024
R30291 net7.n4706 net7.n4705 0.024
R30292 net7.n4793 net7.n4792 0.024
R30293 net7.n4825 net7.n4823 0.024
R30294 net7.n4836 net7.n4834 0.024
R30295 net7.n4932 net7.n4930 0.024
R30296 net7.n4943 net7.n4941 0.024
R30297 net7.n4974 net7.n4972 0.024
R30298 net7.n4992 net7.n4991 0.024
R30299 net7.n5070 net7.n5069 0.024
R30300 net7.n5068 net7.n5067 0.024
R30301 net7.n5155 net7.n5154 0.024
R30302 net7.n5187 net7.n5185 0.024
R30303 net7.n5198 net7.n5196 0.024
R30304 net7.n5294 net7.n5292 0.024
R30305 net7.n5305 net7.n5303 0.024
R30306 net7.n5336 net7.n5334 0.024
R30307 net7.n5354 net7.n5353 0.024
R30308 net7.n5432 net7.n5431 0.024
R30309 net7.n5430 net7.n5429 0.024
R30310 net7.n5517 net7.n5516 0.024
R30311 net7.n5549 net7.n5547 0.024
R30312 net7.n5560 net7.n5558 0.024
R30313 net7.n5656 net7.n5654 0.024
R30314 net7.n5667 net7.n5665 0.024
R30315 net7.n5698 net7.n5696 0.024
R30316 net7.n5716 net7.n5715 0.024
R30317 net7.n5794 net7.n5793 0.024
R30318 net7.n5792 net7.n5791 0.024
R30319 net7.n5879 net7.n5878 0.024
R30320 net7.n5911 net7.n5909 0.024
R30321 net7.n5922 net7.n5920 0.024
R30322 net7.n6018 net7.n6016 0.024
R30323 net7.n6029 net7.n6027 0.024
R30324 net7.n6060 net7.n6058 0.024
R30325 net7.n6078 net7.n6077 0.024
R30326 net7.n6156 net7.n6155 0.024
R30327 net7.n6154 net7.n6153 0.024
R30328 net7.n6241 net7.n6240 0.024
R30329 net7.n6273 net7.n6271 0.024
R30330 net7.n6284 net7.n6282 0.024
R30331 net7.n6380 net7.n6378 0.024
R30332 net7.n6391 net7.n6389 0.024
R30333 net7.n6422 net7.n6420 0.024
R30334 net7.n6440 net7.n6439 0.024
R30335 net7.n6518 net7.n6517 0.024
R30336 net7.n6516 net7.n6515 0.024
R30337 net7.n6603 net7.n6602 0.024
R30338 net7.n6635 net7.n6633 0.024
R30339 net7.n6646 net7.n6644 0.024
R30340 net7.n6742 net7.n6740 0.024
R30341 net7.n6753 net7.n6751 0.024
R30342 net7.n6784 net7.n6782 0.024
R30343 net7.n6802 net7.n6801 0.024
R30344 net7.n6880 net7.n6879 0.024
R30345 net7.n6878 net7.n6877 0.024
R30346 net7.n6965 net7.n6964 0.024
R30347 net7.n6997 net7.n6995 0.024
R30348 net7.n7008 net7.n7006 0.024
R30349 net7.n7104 net7.n7102 0.024
R30350 net7.n7115 net7.n7113 0.024
R30351 net7.n7146 net7.n7144 0.024
R30352 net7.n7164 net7.n7163 0.024
R30353 net7.n3549 net7.n3547 0.022
R30354 net7.n3544 net7.n3543 0.022
R30355 net7.n3615 net7.n3614 0.022
R30356 net7.n3324 net7.n3323 0.022
R30357 net7.n3262 net7.n3261 0.022
R30358 net7.n3267 net7.n3266 0.022
R30359 net7.n3187 net7.n3185 0.022
R30360 net7.n3182 net7.n3181 0.022
R30361 net7.n3253 net7.n3252 0.022
R30362 net7.n2962 net7.n2961 0.022
R30363 net7.n2900 net7.n2899 0.022
R30364 net7.n2905 net7.n2904 0.022
R30365 net7.n2825 net7.n2823 0.022
R30366 net7.n2820 net7.n2819 0.022
R30367 net7.n2891 net7.n2890 0.022
R30368 net7.n2600 net7.n2599 0.022
R30369 net7.n2538 net7.n2537 0.022
R30370 net7.n2543 net7.n2542 0.022
R30371 net7.n2463 net7.n2461 0.022
R30372 net7.n2458 net7.n2457 0.022
R30373 net7.n2529 net7.n2528 0.022
R30374 net7.n2238 net7.n2237 0.022
R30375 net7.n2176 net7.n2175 0.022
R30376 net7.n2181 net7.n2180 0.022
R30377 net7.n2101 net7.n2099 0.022
R30378 net7.n2096 net7.n2095 0.022
R30379 net7.n2167 net7.n2166 0.022
R30380 net7.n1876 net7.n1875 0.022
R30381 net7.n1814 net7.n1813 0.022
R30382 net7.n1819 net7.n1818 0.022
R30383 net7.n1739 net7.n1737 0.022
R30384 net7.n1734 net7.n1733 0.022
R30385 net7.n1805 net7.n1804 0.022
R30386 net7.n1514 net7.n1513 0.022
R30387 net7.n1452 net7.n1451 0.022
R30388 net7.n1457 net7.n1456 0.022
R30389 net7.n1377 net7.n1375 0.022
R30390 net7.n1372 net7.n1371 0.022
R30391 net7.n1443 net7.n1442 0.022
R30392 net7.n1152 net7.n1151 0.022
R30393 net7.n1090 net7.n1089 0.022
R30394 net7.n1095 net7.n1094 0.022
R30395 net7.n1015 net7.n1013 0.022
R30396 net7.n1010 net7.n1009 0.022
R30397 net7.n1081 net7.n1080 0.022
R30398 net7.n790 net7.n789 0.022
R30399 net7.n728 net7.n727 0.022
R30400 net7.n733 net7.n732 0.022
R30401 net7.n653 net7.n651 0.022
R30402 net7.n648 net7.n647 0.022
R30403 net7.n719 net7.n718 0.022
R30404 net7.n428 net7.n427 0.022
R30405 net7.n366 net7.n365 0.022
R30406 net7.n371 net7.n370 0.022
R30407 net7.n292 net7.n290 0.022
R30408 net7.n287 net7.n286 0.022
R30409 net7.n358 net7.n357 0.022
R30410 net7.n67 net7.n66 0.022
R30411 net7.n5 net7.n4 0.022
R30412 net7.n10 net7.n9 0.022
R30413 net7.n3783 net7.n3782 0.022
R30414 net7.n3789 net7.n3788 0.022
R30415 net7.n3743 net7.n3742 0.022
R30416 net7.n3901 net7.n3899 0.022
R30417 net7.n3908 net7.n3907 0.022
R30418 net7.n4144 net7.n4143 0.022
R30419 net7.n4150 net7.n4149 0.022
R30420 net7.n4104 net7.n4103 0.022
R30421 net7.n4262 net7.n4260 0.022
R30422 net7.n4269 net7.n4268 0.022
R30423 net7.n4506 net7.n4505 0.022
R30424 net7.n4512 net7.n4511 0.022
R30425 net7.n4466 net7.n4465 0.022
R30426 net7.n4624 net7.n4622 0.022
R30427 net7.n4631 net7.n4630 0.022
R30428 net7.n4868 net7.n4867 0.022
R30429 net7.n4874 net7.n4873 0.022
R30430 net7.n4828 net7.n4827 0.022
R30431 net7.n4986 net7.n4984 0.022
R30432 net7.n4993 net7.n4992 0.022
R30433 net7.n5230 net7.n5229 0.022
R30434 net7.n5236 net7.n5235 0.022
R30435 net7.n5190 net7.n5189 0.022
R30436 net7.n5348 net7.n5346 0.022
R30437 net7.n5355 net7.n5354 0.022
R30438 net7.n5592 net7.n5591 0.022
R30439 net7.n5598 net7.n5597 0.022
R30440 net7.n5552 net7.n5551 0.022
R30441 net7.n5710 net7.n5708 0.022
R30442 net7.n5717 net7.n5716 0.022
R30443 net7.n5954 net7.n5953 0.022
R30444 net7.n5960 net7.n5959 0.022
R30445 net7.n5914 net7.n5913 0.022
R30446 net7.n6072 net7.n6070 0.022
R30447 net7.n6079 net7.n6078 0.022
R30448 net7.n6316 net7.n6315 0.022
R30449 net7.n6322 net7.n6321 0.022
R30450 net7.n6276 net7.n6275 0.022
R30451 net7.n6434 net7.n6432 0.022
R30452 net7.n6441 net7.n6440 0.022
R30453 net7.n6678 net7.n6677 0.022
R30454 net7.n6684 net7.n6683 0.022
R30455 net7.n6638 net7.n6637 0.022
R30456 net7.n6796 net7.n6794 0.022
R30457 net7.n6803 net7.n6802 0.022
R30458 net7.n7040 net7.n7039 0.022
R30459 net7.n7046 net7.n7045 0.022
R30460 net7.n7000 net7.n6999 0.022
R30461 net7.n7158 net7.n7156 0.022
R30462 net7.n7165 net7.n7164 0.022
R30463 net7.n3560 net7.n3559 0.02
R30464 net7.n3408 net7.n3407 0.02
R30465 net7.n3397 net7.n3396 0.02
R30466 net7.n3614 net7.n3613 0.02
R30467 net7.n3367 net7.n3366 0.02
R30468 net7.n3198 net7.n3197 0.02
R30469 net7.n3046 net7.n3045 0.02
R30470 net7.n3035 net7.n3034 0.02
R30471 net7.n3252 net7.n3251 0.02
R30472 net7.n3005 net7.n3004 0.02
R30473 net7.n2836 net7.n2835 0.02
R30474 net7.n2684 net7.n2683 0.02
R30475 net7.n2673 net7.n2672 0.02
R30476 net7.n2890 net7.n2889 0.02
R30477 net7.n2643 net7.n2642 0.02
R30478 net7.n2474 net7.n2473 0.02
R30479 net7.n2322 net7.n2321 0.02
R30480 net7.n2311 net7.n2310 0.02
R30481 net7.n2528 net7.n2527 0.02
R30482 net7.n2281 net7.n2280 0.02
R30483 net7.n2112 net7.n2111 0.02
R30484 net7.n1960 net7.n1959 0.02
R30485 net7.n1949 net7.n1948 0.02
R30486 net7.n2166 net7.n2165 0.02
R30487 net7.n1919 net7.n1918 0.02
R30488 net7.n1750 net7.n1749 0.02
R30489 net7.n1598 net7.n1597 0.02
R30490 net7.n1587 net7.n1586 0.02
R30491 net7.n1804 net7.n1803 0.02
R30492 net7.n1557 net7.n1556 0.02
R30493 net7.n1388 net7.n1387 0.02
R30494 net7.n1236 net7.n1235 0.02
R30495 net7.n1225 net7.n1224 0.02
R30496 net7.n1442 net7.n1441 0.02
R30497 net7.n1195 net7.n1194 0.02
R30498 net7.n1026 net7.n1025 0.02
R30499 net7.n874 net7.n873 0.02
R30500 net7.n863 net7.n862 0.02
R30501 net7.n1080 net7.n1079 0.02
R30502 net7.n833 net7.n832 0.02
R30503 net7.n664 net7.n663 0.02
R30504 net7.n512 net7.n511 0.02
R30505 net7.n501 net7.n500 0.02
R30506 net7.n718 net7.n717 0.02
R30507 net7.n471 net7.n470 0.02
R30508 net7.n303 net7.n302 0.02
R30509 net7.n151 net7.n150 0.02
R30510 net7.n140 net7.n139 0.02
R30511 net7.n357 net7.n356 0.02
R30512 net7.n110 net7.n109 0.02
R30513 net7.n3652 net7.n3651 0.02
R30514 net7.n3832 net7.n3831 0.02
R30515 net7.n3920 net7.n3919 0.02
R30516 net7.n3628 net7.n3627 0.02
R30517 net7.n3701 net7.n3700 0.02
R30518 net7.n3909 net7.n3908 0.02
R30519 net7.n4013 net7.n4012 0.02
R30520 net7.n4193 net7.n4192 0.02
R30521 net7.n4281 net7.n4280 0.02
R30522 net7.n3989 net7.n3988 0.02
R30523 net7.n4062 net7.n4061 0.02
R30524 net7.n4270 net7.n4269 0.02
R30525 net7.n4375 net7.n4374 0.02
R30526 net7.n4555 net7.n4554 0.02
R30527 net7.n4643 net7.n4642 0.02
R30528 net7.n4351 net7.n4350 0.02
R30529 net7.n4424 net7.n4423 0.02
R30530 net7.n4632 net7.n4631 0.02
R30531 net7.n4737 net7.n4736 0.02
R30532 net7.n4917 net7.n4916 0.02
R30533 net7.n5005 net7.n5004 0.02
R30534 net7.n4713 net7.n4712 0.02
R30535 net7.n4786 net7.n4785 0.02
R30536 net7.n4994 net7.n4993 0.02
R30537 net7.n5099 net7.n5098 0.02
R30538 net7.n5279 net7.n5278 0.02
R30539 net7.n5367 net7.n5366 0.02
R30540 net7.n5075 net7.n5074 0.02
R30541 net7.n5148 net7.n5147 0.02
R30542 net7.n5356 net7.n5355 0.02
R30543 net7.n5461 net7.n5460 0.02
R30544 net7.n5641 net7.n5640 0.02
R30545 net7.n5729 net7.n5728 0.02
R30546 net7.n5437 net7.n5436 0.02
R30547 net7.n5510 net7.n5509 0.02
R30548 net7.n5718 net7.n5717 0.02
R30549 net7.n5823 net7.n5822 0.02
R30550 net7.n6003 net7.n6002 0.02
R30551 net7.n6091 net7.n6090 0.02
R30552 net7.n5799 net7.n5798 0.02
R30553 net7.n5872 net7.n5871 0.02
R30554 net7.n6080 net7.n6079 0.02
R30555 net7.n6185 net7.n6184 0.02
R30556 net7.n6365 net7.n6364 0.02
R30557 net7.n6453 net7.n6452 0.02
R30558 net7.n6161 net7.n6160 0.02
R30559 net7.n6234 net7.n6233 0.02
R30560 net7.n6442 net7.n6441 0.02
R30561 net7.n6547 net7.n6546 0.02
R30562 net7.n6727 net7.n6726 0.02
R30563 net7.n6815 net7.n6814 0.02
R30564 net7.n6523 net7.n6522 0.02
R30565 net7.n6596 net7.n6595 0.02
R30566 net7.n6804 net7.n6803 0.02
R30567 net7.n6909 net7.n6908 0.02
R30568 net7.n7089 net7.n7088 0.02
R30569 net7.n7177 net7.n7176 0.02
R30570 net7.n6885 net7.n6884 0.02
R30571 net7.n6958 net7.n6957 0.02
R30572 net7.n7166 net7.n7165 0.02
R30573 net7.n3317 net7.n3316 0.018
R30574 net7.n2955 net7.n2954 0.018
R30575 net7.n2593 net7.n2592 0.018
R30576 net7.n2231 net7.n2230 0.018
R30577 net7.n1869 net7.n1868 0.018
R30578 net7.n1507 net7.n1506 0.018
R30579 net7.n1145 net7.n1144 0.018
R30580 net7.n783 net7.n782 0.018
R30581 net7.n421 net7.n420 0.018
R30582 net7.n60 net7.n59 0.018
R30583 net7.n3572 net7.n3571 0.017
R30584 net7.n3292 net7.n3288 0.017
R30585 net7.n3318 net7.n3317 0.017
R30586 net7.n3210 net7.n3209 0.017
R30587 net7.n2930 net7.n2926 0.017
R30588 net7.n2956 net7.n2955 0.017
R30589 net7.n2848 net7.n2847 0.017
R30590 net7.n2568 net7.n2564 0.017
R30591 net7.n2594 net7.n2593 0.017
R30592 net7.n2486 net7.n2485 0.017
R30593 net7.n2206 net7.n2202 0.017
R30594 net7.n2232 net7.n2231 0.017
R30595 net7.n2124 net7.n2123 0.017
R30596 net7.n1844 net7.n1840 0.017
R30597 net7.n1870 net7.n1869 0.017
R30598 net7.n1762 net7.n1761 0.017
R30599 net7.n1482 net7.n1478 0.017
R30600 net7.n1508 net7.n1507 0.017
R30601 net7.n1400 net7.n1399 0.017
R30602 net7.n1120 net7.n1116 0.017
R30603 net7.n1146 net7.n1145 0.017
R30604 net7.n1038 net7.n1037 0.017
R30605 net7.n758 net7.n754 0.017
R30606 net7.n784 net7.n783 0.017
R30607 net7.n676 net7.n675 0.017
R30608 net7.n396 net7.n392 0.017
R30609 net7.n422 net7.n421 0.017
R30610 net7.n315 net7.n314 0.017
R30611 net7.n35 net7.n31 0.017
R30612 net7.n61 net7.n60 0.017
R30613 net7.n3661 net7.n3660 0.017
R30614 net7.n3935 net7.n3934 0.017
R30615 net7.n3959 net7.n3955 0.017
R30616 net7.n3865 net7.n3864 0.017
R30617 net7.n3889 net7.n3888 0.017
R30618 net7.n4022 net7.n4021 0.017
R30619 net7.n4296 net7.n4295 0.017
R30620 net7.n4320 net7.n4316 0.017
R30621 net7.n4226 net7.n4225 0.017
R30622 net7.n4250 net7.n4249 0.017
R30623 net7.n4384 net7.n4383 0.017
R30624 net7.n4658 net7.n4657 0.017
R30625 net7.n4682 net7.n4678 0.017
R30626 net7.n4588 net7.n4587 0.017
R30627 net7.n4612 net7.n4611 0.017
R30628 net7.n4746 net7.n4745 0.017
R30629 net7.n5020 net7.n5019 0.017
R30630 net7.n5044 net7.n5040 0.017
R30631 net7.n4950 net7.n4949 0.017
R30632 net7.n4974 net7.n4973 0.017
R30633 net7.n5108 net7.n5107 0.017
R30634 net7.n5382 net7.n5381 0.017
R30635 net7.n5406 net7.n5402 0.017
R30636 net7.n5312 net7.n5311 0.017
R30637 net7.n5336 net7.n5335 0.017
R30638 net7.n5470 net7.n5469 0.017
R30639 net7.n5744 net7.n5743 0.017
R30640 net7.n5768 net7.n5764 0.017
R30641 net7.n5674 net7.n5673 0.017
R30642 net7.n5698 net7.n5697 0.017
R30643 net7.n5832 net7.n5831 0.017
R30644 net7.n6106 net7.n6105 0.017
R30645 net7.n6130 net7.n6126 0.017
R30646 net7.n6036 net7.n6035 0.017
R30647 net7.n6060 net7.n6059 0.017
R30648 net7.n6194 net7.n6193 0.017
R30649 net7.n6468 net7.n6467 0.017
R30650 net7.n6492 net7.n6488 0.017
R30651 net7.n6398 net7.n6397 0.017
R30652 net7.n6422 net7.n6421 0.017
R30653 net7.n6556 net7.n6555 0.017
R30654 net7.n6830 net7.n6829 0.017
R30655 net7.n6854 net7.n6850 0.017
R30656 net7.n6760 net7.n6759 0.017
R30657 net7.n6784 net7.n6783 0.017
R30658 net7.n6918 net7.n6917 0.017
R30659 net7.n7192 net7.n7191 0.017
R30660 net7.n7216 net7.n7212 0.017
R30661 net7.n7122 net7.n7121 0.017
R30662 net7.n7146 net7.n7145 0.017
R30663 net7.n3509 net7.n3508 0.016
R30664 net7.n3485 net7.n3484 0.016
R30665 net7.n3467 net7.n3466 0.016
R30666 net7.n3441 net7.n3440 0.016
R30667 net7.n3423 net7.n3422 0.016
R30668 net7.n3352 net7.n3351 0.016
R30669 net7.n3328 net7.n3327 0.016
R30670 net7.n3147 net7.n3146 0.016
R30671 net7.n3123 net7.n3122 0.016
R30672 net7.n3105 net7.n3104 0.016
R30673 net7.n3079 net7.n3078 0.016
R30674 net7.n3061 net7.n3060 0.016
R30675 net7.n2990 net7.n2989 0.016
R30676 net7.n2966 net7.n2965 0.016
R30677 net7.n2785 net7.n2784 0.016
R30678 net7.n2761 net7.n2760 0.016
R30679 net7.n2743 net7.n2742 0.016
R30680 net7.n2717 net7.n2716 0.016
R30681 net7.n2699 net7.n2698 0.016
R30682 net7.n2628 net7.n2627 0.016
R30683 net7.n2604 net7.n2603 0.016
R30684 net7.n2423 net7.n2422 0.016
R30685 net7.n2399 net7.n2398 0.016
R30686 net7.n2381 net7.n2380 0.016
R30687 net7.n2355 net7.n2354 0.016
R30688 net7.n2337 net7.n2336 0.016
R30689 net7.n2266 net7.n2265 0.016
R30690 net7.n2242 net7.n2241 0.016
R30691 net7.n2061 net7.n2060 0.016
R30692 net7.n2037 net7.n2036 0.016
R30693 net7.n2019 net7.n2018 0.016
R30694 net7.n1993 net7.n1992 0.016
R30695 net7.n1975 net7.n1974 0.016
R30696 net7.n1904 net7.n1903 0.016
R30697 net7.n1880 net7.n1879 0.016
R30698 net7.n1699 net7.n1698 0.016
R30699 net7.n1675 net7.n1674 0.016
R30700 net7.n1657 net7.n1656 0.016
R30701 net7.n1631 net7.n1630 0.016
R30702 net7.n1613 net7.n1612 0.016
R30703 net7.n1542 net7.n1541 0.016
R30704 net7.n1518 net7.n1517 0.016
R30705 net7.n1337 net7.n1336 0.016
R30706 net7.n1313 net7.n1312 0.016
R30707 net7.n1295 net7.n1294 0.016
R30708 net7.n1269 net7.n1268 0.016
R30709 net7.n1251 net7.n1250 0.016
R30710 net7.n1180 net7.n1179 0.016
R30711 net7.n1156 net7.n1155 0.016
R30712 net7.n975 net7.n974 0.016
R30713 net7.n951 net7.n950 0.016
R30714 net7.n933 net7.n932 0.016
R30715 net7.n907 net7.n906 0.016
R30716 net7.n889 net7.n888 0.016
R30717 net7.n818 net7.n817 0.016
R30718 net7.n794 net7.n793 0.016
R30719 net7.n613 net7.n612 0.016
R30720 net7.n589 net7.n588 0.016
R30721 net7.n571 net7.n570 0.016
R30722 net7.n545 net7.n544 0.016
R30723 net7.n527 net7.n526 0.016
R30724 net7.n456 net7.n455 0.016
R30725 net7.n432 net7.n431 0.016
R30726 net7.n252 net7.n251 0.016
R30727 net7.n228 net7.n227 0.016
R30728 net7.n210 net7.n209 0.016
R30729 net7.n184 net7.n183 0.016
R30730 net7.n166 net7.n165 0.016
R30731 net7.n95 net7.n94 0.016
R30732 net7.n71 net7.n70 0.016
R30733 net7.n3711 net7.n3710 0.016
R30734 net7.n3728 net7.n3727 0.016
R30735 net7.n3754 net7.n3753 0.016
R30736 net7.n3773 net7.n3772 0.016
R30737 net7.n3861 net7.n3860 0.016
R30738 net7.n3877 net7.n3876 0.016
R30739 net7.n3904 net7.n3903 0.016
R30740 net7.n4072 net7.n4071 0.016
R30741 net7.n4089 net7.n4088 0.016
R30742 net7.n4115 net7.n4114 0.016
R30743 net7.n4134 net7.n4133 0.016
R30744 net7.n4222 net7.n4221 0.016
R30745 net7.n4238 net7.n4237 0.016
R30746 net7.n4265 net7.n4264 0.016
R30747 net7.n4434 net7.n4433 0.016
R30748 net7.n4451 net7.n4450 0.016
R30749 net7.n4477 net7.n4476 0.016
R30750 net7.n4496 net7.n4495 0.016
R30751 net7.n4584 net7.n4583 0.016
R30752 net7.n4600 net7.n4599 0.016
R30753 net7.n4627 net7.n4626 0.016
R30754 net7.n4796 net7.n4795 0.016
R30755 net7.n4813 net7.n4812 0.016
R30756 net7.n4839 net7.n4838 0.016
R30757 net7.n4858 net7.n4857 0.016
R30758 net7.n4946 net7.n4945 0.016
R30759 net7.n4962 net7.n4961 0.016
R30760 net7.n4989 net7.n4988 0.016
R30761 net7.n5158 net7.n5157 0.016
R30762 net7.n5175 net7.n5174 0.016
R30763 net7.n5201 net7.n5200 0.016
R30764 net7.n5220 net7.n5219 0.016
R30765 net7.n5308 net7.n5307 0.016
R30766 net7.n5324 net7.n5323 0.016
R30767 net7.n5351 net7.n5350 0.016
R30768 net7.n5520 net7.n5519 0.016
R30769 net7.n5537 net7.n5536 0.016
R30770 net7.n5563 net7.n5562 0.016
R30771 net7.n5582 net7.n5581 0.016
R30772 net7.n5670 net7.n5669 0.016
R30773 net7.n5686 net7.n5685 0.016
R30774 net7.n5713 net7.n5712 0.016
R30775 net7.n5882 net7.n5881 0.016
R30776 net7.n5899 net7.n5898 0.016
R30777 net7.n5925 net7.n5924 0.016
R30778 net7.n5944 net7.n5943 0.016
R30779 net7.n6032 net7.n6031 0.016
R30780 net7.n6048 net7.n6047 0.016
R30781 net7.n6075 net7.n6074 0.016
R30782 net7.n6244 net7.n6243 0.016
R30783 net7.n6261 net7.n6260 0.016
R30784 net7.n6287 net7.n6286 0.016
R30785 net7.n6306 net7.n6305 0.016
R30786 net7.n6394 net7.n6393 0.016
R30787 net7.n6410 net7.n6409 0.016
R30788 net7.n6437 net7.n6436 0.016
R30789 net7.n6606 net7.n6605 0.016
R30790 net7.n6623 net7.n6622 0.016
R30791 net7.n6649 net7.n6648 0.016
R30792 net7.n6668 net7.n6667 0.016
R30793 net7.n6756 net7.n6755 0.016
R30794 net7.n6772 net7.n6771 0.016
R30795 net7.n6799 net7.n6798 0.016
R30796 net7.n6968 net7.n6967 0.016
R30797 net7.n6985 net7.n6984 0.016
R30798 net7.n7011 net7.n7010 0.016
R30799 net7.n7030 net7.n7029 0.016
R30800 net7.n7118 net7.n7117 0.016
R30801 net7.n7134 net7.n7133 0.016
R30802 net7.n7161 net7.n7160 0.016
R30803 net7.n3600 net7.n3599 0.015
R30804 net7.n3594 net7.n3593 0.015
R30805 net7.n3592 net7.n3591 0.015
R30806 net7.n3409 net7.n3408 0.015
R30807 net7.n3294 net7.n3293 0.015
R30808 net7.n3300 net7.n3299 0.015
R30809 net7.n3505 net7.n3504 0.015
R30810 net7.n3495 net7.n3492 0.015
R30811 net7.n3494 net7.n3493 0.015
R30812 net7.n3472 net7.n3471 0.015
R30813 net7.n3463 net7.n3462 0.015
R30814 net7.n3452 net7.n3451 0.015
R30815 net7.n3419 net7.n3418 0.015
R30816 net7.n3368 net7.n3367 0.015
R30817 net7.n3363 net7.n3362 0.015
R30818 net7.n3323 net7.n3322 0.015
R30819 net7.n3260 net7.n3259 0.015
R30820 net7.n3238 net7.n3237 0.015
R30821 net7.n3232 net7.n3231 0.015
R30822 net7.n3230 net7.n3229 0.015
R30823 net7.n3047 net7.n3046 0.015
R30824 net7.n2932 net7.n2931 0.015
R30825 net7.n2938 net7.n2937 0.015
R30826 net7.n3143 net7.n3142 0.015
R30827 net7.n3133 net7.n3130 0.015
R30828 net7.n3132 net7.n3131 0.015
R30829 net7.n3110 net7.n3109 0.015
R30830 net7.n3101 net7.n3100 0.015
R30831 net7.n3090 net7.n3089 0.015
R30832 net7.n3057 net7.n3056 0.015
R30833 net7.n3006 net7.n3005 0.015
R30834 net7.n3001 net7.n3000 0.015
R30835 net7.n2961 net7.n2960 0.015
R30836 net7.n2898 net7.n2897 0.015
R30837 net7.n2876 net7.n2875 0.015
R30838 net7.n2870 net7.n2869 0.015
R30839 net7.n2868 net7.n2867 0.015
R30840 net7.n2685 net7.n2684 0.015
R30841 net7.n2570 net7.n2569 0.015
R30842 net7.n2576 net7.n2575 0.015
R30843 net7.n2781 net7.n2780 0.015
R30844 net7.n2771 net7.n2768 0.015
R30845 net7.n2770 net7.n2769 0.015
R30846 net7.n2748 net7.n2747 0.015
R30847 net7.n2739 net7.n2738 0.015
R30848 net7.n2728 net7.n2727 0.015
R30849 net7.n2695 net7.n2694 0.015
R30850 net7.n2644 net7.n2643 0.015
R30851 net7.n2639 net7.n2638 0.015
R30852 net7.n2599 net7.n2598 0.015
R30853 net7.n2536 net7.n2535 0.015
R30854 net7.n2514 net7.n2513 0.015
R30855 net7.n2508 net7.n2507 0.015
R30856 net7.n2506 net7.n2505 0.015
R30857 net7.n2323 net7.n2322 0.015
R30858 net7.n2208 net7.n2207 0.015
R30859 net7.n2214 net7.n2213 0.015
R30860 net7.n2419 net7.n2418 0.015
R30861 net7.n2409 net7.n2406 0.015
R30862 net7.n2408 net7.n2407 0.015
R30863 net7.n2386 net7.n2385 0.015
R30864 net7.n2377 net7.n2376 0.015
R30865 net7.n2366 net7.n2365 0.015
R30866 net7.n2333 net7.n2332 0.015
R30867 net7.n2282 net7.n2281 0.015
R30868 net7.n2277 net7.n2276 0.015
R30869 net7.n2237 net7.n2236 0.015
R30870 net7.n2174 net7.n2173 0.015
R30871 net7.n2152 net7.n2151 0.015
R30872 net7.n2146 net7.n2145 0.015
R30873 net7.n2144 net7.n2143 0.015
R30874 net7.n1961 net7.n1960 0.015
R30875 net7.n1846 net7.n1845 0.015
R30876 net7.n1852 net7.n1851 0.015
R30877 net7.n2057 net7.n2056 0.015
R30878 net7.n2047 net7.n2044 0.015
R30879 net7.n2046 net7.n2045 0.015
R30880 net7.n2024 net7.n2023 0.015
R30881 net7.n2015 net7.n2014 0.015
R30882 net7.n2004 net7.n2003 0.015
R30883 net7.n1971 net7.n1970 0.015
R30884 net7.n1920 net7.n1919 0.015
R30885 net7.n1915 net7.n1914 0.015
R30886 net7.n1875 net7.n1874 0.015
R30887 net7.n1812 net7.n1811 0.015
R30888 net7.n1790 net7.n1789 0.015
R30889 net7.n1784 net7.n1783 0.015
R30890 net7.n1782 net7.n1781 0.015
R30891 net7.n1599 net7.n1598 0.015
R30892 net7.n1484 net7.n1483 0.015
R30893 net7.n1490 net7.n1489 0.015
R30894 net7.n1695 net7.n1694 0.015
R30895 net7.n1685 net7.n1682 0.015
R30896 net7.n1684 net7.n1683 0.015
R30897 net7.n1662 net7.n1661 0.015
R30898 net7.n1653 net7.n1652 0.015
R30899 net7.n1642 net7.n1641 0.015
R30900 net7.n1609 net7.n1608 0.015
R30901 net7.n1558 net7.n1557 0.015
R30902 net7.n1553 net7.n1552 0.015
R30903 net7.n1513 net7.n1512 0.015
R30904 net7.n1450 net7.n1449 0.015
R30905 net7.n1428 net7.n1427 0.015
R30906 net7.n1422 net7.n1421 0.015
R30907 net7.n1420 net7.n1419 0.015
R30908 net7.n1237 net7.n1236 0.015
R30909 net7.n1122 net7.n1121 0.015
R30910 net7.n1128 net7.n1127 0.015
R30911 net7.n1333 net7.n1332 0.015
R30912 net7.n1323 net7.n1320 0.015
R30913 net7.n1322 net7.n1321 0.015
R30914 net7.n1300 net7.n1299 0.015
R30915 net7.n1291 net7.n1290 0.015
R30916 net7.n1280 net7.n1279 0.015
R30917 net7.n1247 net7.n1246 0.015
R30918 net7.n1196 net7.n1195 0.015
R30919 net7.n1191 net7.n1190 0.015
R30920 net7.n1151 net7.n1150 0.015
R30921 net7.n1088 net7.n1087 0.015
R30922 net7.n1066 net7.n1065 0.015
R30923 net7.n1060 net7.n1059 0.015
R30924 net7.n1058 net7.n1057 0.015
R30925 net7.n875 net7.n874 0.015
R30926 net7.n760 net7.n759 0.015
R30927 net7.n766 net7.n765 0.015
R30928 net7.n971 net7.n970 0.015
R30929 net7.n961 net7.n958 0.015
R30930 net7.n960 net7.n959 0.015
R30931 net7.n938 net7.n937 0.015
R30932 net7.n929 net7.n928 0.015
R30933 net7.n918 net7.n917 0.015
R30934 net7.n885 net7.n884 0.015
R30935 net7.n834 net7.n833 0.015
R30936 net7.n829 net7.n828 0.015
R30937 net7.n789 net7.n788 0.015
R30938 net7.n726 net7.n725 0.015
R30939 net7.n704 net7.n703 0.015
R30940 net7.n698 net7.n697 0.015
R30941 net7.n696 net7.n695 0.015
R30942 net7.n513 net7.n512 0.015
R30943 net7.n398 net7.n397 0.015
R30944 net7.n404 net7.n403 0.015
R30945 net7.n609 net7.n608 0.015
R30946 net7.n599 net7.n596 0.015
R30947 net7.n598 net7.n597 0.015
R30948 net7.n576 net7.n575 0.015
R30949 net7.n567 net7.n566 0.015
R30950 net7.n556 net7.n555 0.015
R30951 net7.n523 net7.n522 0.015
R30952 net7.n472 net7.n471 0.015
R30953 net7.n467 net7.n466 0.015
R30954 net7.n427 net7.n426 0.015
R30955 net7.n364 net7.n363 0.015
R30956 net7.n343 net7.n342 0.015
R30957 net7.n337 net7.n336 0.015
R30958 net7.n335 net7.n334 0.015
R30959 net7.n152 net7.n151 0.015
R30960 net7.n37 net7.n36 0.015
R30961 net7.n43 net7.n42 0.015
R30962 net7.n248 net7.n247 0.015
R30963 net7.n238 net7.n235 0.015
R30964 net7.n237 net7.n236 0.015
R30965 net7.n215 net7.n214 0.015
R30966 net7.n206 net7.n205 0.015
R30967 net7.n195 net7.n194 0.015
R30968 net7.n162 net7.n161 0.015
R30969 net7.n111 net7.n110 0.015
R30970 net7.n106 net7.n105 0.015
R30971 net7.n66 net7.n65 0.015
R30972 net7.n3 net7.n2 0.015
R30973 net7.n3686 net7.n3685 0.015
R30974 net7.n3680 net7.n3679 0.015
R30975 net7.n3678 net7.n3677 0.015
R30976 net7.n3833 net7.n3832 0.015
R30977 net7.n3961 net7.n3960 0.015
R30978 net7.n3967 net7.n3966 0.015
R30979 net7.n3622 net7.n3621 0.015
R30980 net7.n3702 net7.n3701 0.015
R30981 net7.n3707 net7.n3706 0.015
R30982 net7.n3738 net7.n3737 0.015
R30983 net7.n3749 net7.n3748 0.015
R30984 net7.n3758 net7.n3757 0.015
R30985 net7.n3845 net7.n3844 0.015
R30986 net7.n3847 net7.n3846 0.015
R30987 net7.n3856 net7.n3855 0.015
R30988 net7.n3887 net7.n3886 0.015
R30989 net7.n3898 net7.n3897 0.015
R30990 net7.n4047 net7.n4046 0.015
R30991 net7.n4041 net7.n4040 0.015
R30992 net7.n4039 net7.n4038 0.015
R30993 net7.n4194 net7.n4193 0.015
R30994 net7.n4322 net7.n4321 0.015
R30995 net7.n4328 net7.n4327 0.015
R30996 net7.n3983 net7.n3982 0.015
R30997 net7.n4063 net7.n4062 0.015
R30998 net7.n4068 net7.n4067 0.015
R30999 net7.n4099 net7.n4098 0.015
R31000 net7.n4110 net7.n4109 0.015
R31001 net7.n4119 net7.n4118 0.015
R31002 net7.n4206 net7.n4205 0.015
R31003 net7.n4208 net7.n4207 0.015
R31004 net7.n4217 net7.n4216 0.015
R31005 net7.n4248 net7.n4247 0.015
R31006 net7.n4259 net7.n4258 0.015
R31007 net7.n4409 net7.n4408 0.015
R31008 net7.n4403 net7.n4402 0.015
R31009 net7.n4401 net7.n4400 0.015
R31010 net7.n4556 net7.n4555 0.015
R31011 net7.n4684 net7.n4683 0.015
R31012 net7.n4690 net7.n4689 0.015
R31013 net7.n4345 net7.n4344 0.015
R31014 net7.n4425 net7.n4424 0.015
R31015 net7.n4430 net7.n4429 0.015
R31016 net7.n4461 net7.n4460 0.015
R31017 net7.n4472 net7.n4471 0.015
R31018 net7.n4481 net7.n4480 0.015
R31019 net7.n4568 net7.n4567 0.015
R31020 net7.n4570 net7.n4569 0.015
R31021 net7.n4579 net7.n4578 0.015
R31022 net7.n4610 net7.n4609 0.015
R31023 net7.n4621 net7.n4620 0.015
R31024 net7.n4771 net7.n4770 0.015
R31025 net7.n4765 net7.n4764 0.015
R31026 net7.n4763 net7.n4762 0.015
R31027 net7.n4918 net7.n4917 0.015
R31028 net7.n5046 net7.n5045 0.015
R31029 net7.n5052 net7.n5051 0.015
R31030 net7.n4707 net7.n4706 0.015
R31031 net7.n4787 net7.n4786 0.015
R31032 net7.n4792 net7.n4791 0.015
R31033 net7.n4823 net7.n4822 0.015
R31034 net7.n4834 net7.n4833 0.015
R31035 net7.n4843 net7.n4842 0.015
R31036 net7.n4930 net7.n4929 0.015
R31037 net7.n4932 net7.n4931 0.015
R31038 net7.n4941 net7.n4940 0.015
R31039 net7.n4972 net7.n4971 0.015
R31040 net7.n4983 net7.n4982 0.015
R31041 net7.n5133 net7.n5132 0.015
R31042 net7.n5127 net7.n5126 0.015
R31043 net7.n5125 net7.n5124 0.015
R31044 net7.n5280 net7.n5279 0.015
R31045 net7.n5408 net7.n5407 0.015
R31046 net7.n5414 net7.n5413 0.015
R31047 net7.n5069 net7.n5068 0.015
R31048 net7.n5149 net7.n5148 0.015
R31049 net7.n5154 net7.n5153 0.015
R31050 net7.n5185 net7.n5184 0.015
R31051 net7.n5196 net7.n5195 0.015
R31052 net7.n5205 net7.n5204 0.015
R31053 net7.n5292 net7.n5291 0.015
R31054 net7.n5294 net7.n5293 0.015
R31055 net7.n5303 net7.n5302 0.015
R31056 net7.n5334 net7.n5333 0.015
R31057 net7.n5345 net7.n5344 0.015
R31058 net7.n5495 net7.n5494 0.015
R31059 net7.n5489 net7.n5488 0.015
R31060 net7.n5487 net7.n5486 0.015
R31061 net7.n5642 net7.n5641 0.015
R31062 net7.n5770 net7.n5769 0.015
R31063 net7.n5776 net7.n5775 0.015
R31064 net7.n5431 net7.n5430 0.015
R31065 net7.n5511 net7.n5510 0.015
R31066 net7.n5516 net7.n5515 0.015
R31067 net7.n5547 net7.n5546 0.015
R31068 net7.n5558 net7.n5557 0.015
R31069 net7.n5567 net7.n5566 0.015
R31070 net7.n5654 net7.n5653 0.015
R31071 net7.n5656 net7.n5655 0.015
R31072 net7.n5665 net7.n5664 0.015
R31073 net7.n5696 net7.n5695 0.015
R31074 net7.n5707 net7.n5706 0.015
R31075 net7.n5857 net7.n5856 0.015
R31076 net7.n5851 net7.n5850 0.015
R31077 net7.n5849 net7.n5848 0.015
R31078 net7.n6004 net7.n6003 0.015
R31079 net7.n6132 net7.n6131 0.015
R31080 net7.n6138 net7.n6137 0.015
R31081 net7.n5793 net7.n5792 0.015
R31082 net7.n5873 net7.n5872 0.015
R31083 net7.n5878 net7.n5877 0.015
R31084 net7.n5909 net7.n5908 0.015
R31085 net7.n5920 net7.n5919 0.015
R31086 net7.n5929 net7.n5928 0.015
R31087 net7.n6016 net7.n6015 0.015
R31088 net7.n6018 net7.n6017 0.015
R31089 net7.n6027 net7.n6026 0.015
R31090 net7.n6058 net7.n6057 0.015
R31091 net7.n6069 net7.n6068 0.015
R31092 net7.n6219 net7.n6218 0.015
R31093 net7.n6213 net7.n6212 0.015
R31094 net7.n6211 net7.n6210 0.015
R31095 net7.n6366 net7.n6365 0.015
R31096 net7.n6494 net7.n6493 0.015
R31097 net7.n6500 net7.n6499 0.015
R31098 net7.n6155 net7.n6154 0.015
R31099 net7.n6235 net7.n6234 0.015
R31100 net7.n6240 net7.n6239 0.015
R31101 net7.n6271 net7.n6270 0.015
R31102 net7.n6282 net7.n6281 0.015
R31103 net7.n6291 net7.n6290 0.015
R31104 net7.n6378 net7.n6377 0.015
R31105 net7.n6380 net7.n6379 0.015
R31106 net7.n6389 net7.n6388 0.015
R31107 net7.n6420 net7.n6419 0.015
R31108 net7.n6431 net7.n6430 0.015
R31109 net7.n6581 net7.n6580 0.015
R31110 net7.n6575 net7.n6574 0.015
R31111 net7.n6573 net7.n6572 0.015
R31112 net7.n6728 net7.n6727 0.015
R31113 net7.n6856 net7.n6855 0.015
R31114 net7.n6862 net7.n6861 0.015
R31115 net7.n6517 net7.n6516 0.015
R31116 net7.n6597 net7.n6596 0.015
R31117 net7.n6602 net7.n6601 0.015
R31118 net7.n6633 net7.n6632 0.015
R31119 net7.n6644 net7.n6643 0.015
R31120 net7.n6653 net7.n6652 0.015
R31121 net7.n6740 net7.n6739 0.015
R31122 net7.n6742 net7.n6741 0.015
R31123 net7.n6751 net7.n6750 0.015
R31124 net7.n6782 net7.n6781 0.015
R31125 net7.n6793 net7.n6792 0.015
R31126 net7.n6943 net7.n6942 0.015
R31127 net7.n6937 net7.n6936 0.015
R31128 net7.n6935 net7.n6934 0.015
R31129 net7.n7090 net7.n7089 0.015
R31130 net7.n7218 net7.n7217 0.015
R31131 net7.n7224 net7.n7223 0.015
R31132 net7.n6879 net7.n6878 0.015
R31133 net7.n6959 net7.n6958 0.015
R31134 net7.n6964 net7.n6963 0.015
R31135 net7.n6995 net7.n6994 0.015
R31136 net7.n7006 net7.n7005 0.015
R31137 net7.n7015 net7.n7014 0.015
R31138 net7.n7102 net7.n7101 0.015
R31139 net7.n7104 net7.n7103 0.015
R31140 net7.n7113 net7.n7112 0.015
R31141 net7.n7144 net7.n7143 0.015
R31142 net7.n7155 net7.n7154 0.015
R31143 net7.n3603 net7.n3600 0.013
R31144 net7.n3543 net7.n3542 0.013
R31145 net7.n3303 net7.n3300 0.013
R31146 net7.n3506 net7.n3503 0.013
R31147 net7.n3453 net7.n3450 0.013
R31148 net7.n3426 net7.n3425 0.013
R31149 net7.n3263 net7.n3262 0.013
R31150 net7.n3241 net7.n3238 0.013
R31151 net7.n3181 net7.n3180 0.013
R31152 net7.n2941 net7.n2938 0.013
R31153 net7.n3144 net7.n3141 0.013
R31154 net7.n3091 net7.n3088 0.013
R31155 net7.n3064 net7.n3063 0.013
R31156 net7.n2901 net7.n2900 0.013
R31157 net7.n2879 net7.n2876 0.013
R31158 net7.n2819 net7.n2818 0.013
R31159 net7.n2579 net7.n2576 0.013
R31160 net7.n2782 net7.n2779 0.013
R31161 net7.n2729 net7.n2726 0.013
R31162 net7.n2702 net7.n2701 0.013
R31163 net7.n2539 net7.n2538 0.013
R31164 net7.n2517 net7.n2514 0.013
R31165 net7.n2457 net7.n2456 0.013
R31166 net7.n2217 net7.n2214 0.013
R31167 net7.n2420 net7.n2417 0.013
R31168 net7.n2367 net7.n2364 0.013
R31169 net7.n2340 net7.n2339 0.013
R31170 net7.n2177 net7.n2176 0.013
R31171 net7.n2155 net7.n2152 0.013
R31172 net7.n2095 net7.n2094 0.013
R31173 net7.n1855 net7.n1852 0.013
R31174 net7.n2058 net7.n2055 0.013
R31175 net7.n2005 net7.n2002 0.013
R31176 net7.n1978 net7.n1977 0.013
R31177 net7.n1815 net7.n1814 0.013
R31178 net7.n1793 net7.n1790 0.013
R31179 net7.n1733 net7.n1732 0.013
R31180 net7.n1493 net7.n1490 0.013
R31181 net7.n1696 net7.n1693 0.013
R31182 net7.n1643 net7.n1640 0.013
R31183 net7.n1616 net7.n1615 0.013
R31184 net7.n1453 net7.n1452 0.013
R31185 net7.n1431 net7.n1428 0.013
R31186 net7.n1371 net7.n1370 0.013
R31187 net7.n1131 net7.n1128 0.013
R31188 net7.n1334 net7.n1331 0.013
R31189 net7.n1281 net7.n1278 0.013
R31190 net7.n1254 net7.n1253 0.013
R31191 net7.n1091 net7.n1090 0.013
R31192 net7.n1069 net7.n1066 0.013
R31193 net7.n1009 net7.n1008 0.013
R31194 net7.n769 net7.n766 0.013
R31195 net7.n972 net7.n969 0.013
R31196 net7.n919 net7.n916 0.013
R31197 net7.n892 net7.n891 0.013
R31198 net7.n729 net7.n728 0.013
R31199 net7.n707 net7.n704 0.013
R31200 net7.n647 net7.n646 0.013
R31201 net7.n407 net7.n404 0.013
R31202 net7.n610 net7.n607 0.013
R31203 net7.n557 net7.n554 0.013
R31204 net7.n530 net7.n529 0.013
R31205 net7.n367 net7.n366 0.013
R31206 net7.n346 net7.n343 0.013
R31207 net7.n286 net7.n285 0.013
R31208 net7.n46 net7.n43 0.013
R31209 net7.n249 net7.n246 0.013
R31210 net7.n196 net7.n193 0.013
R31211 net7.n169 net7.n168 0.013
R31212 net7.n6 net7.n5 0.013
R31213 net7.n3687 net7.n3686 0.013
R31214 net7.n3790 net7.n3789 0.013
R31215 net7.n3970 net7.n3967 0.013
R31216 net7.n3624 net7.n3623 0.013
R31217 net7.n3744 net7.n3743 0.013
R31218 net7.n3901 net7.n3900 0.013
R31219 net7.n4048 net7.n4047 0.013
R31220 net7.n4151 net7.n4150 0.013
R31221 net7.n4331 net7.n4328 0.013
R31222 net7.n3985 net7.n3984 0.013
R31223 net7.n4105 net7.n4104 0.013
R31224 net7.n4262 net7.n4261 0.013
R31225 net7.n4410 net7.n4409 0.013
R31226 net7.n4513 net7.n4512 0.013
R31227 net7.n4693 net7.n4690 0.013
R31228 net7.n4347 net7.n4346 0.013
R31229 net7.n4467 net7.n4466 0.013
R31230 net7.n4624 net7.n4623 0.013
R31231 net7.n4772 net7.n4771 0.013
R31232 net7.n4875 net7.n4874 0.013
R31233 net7.n5055 net7.n5052 0.013
R31234 net7.n4709 net7.n4708 0.013
R31235 net7.n4829 net7.n4828 0.013
R31236 net7.n4986 net7.n4985 0.013
R31237 net7.n5134 net7.n5133 0.013
R31238 net7.n5237 net7.n5236 0.013
R31239 net7.n5417 net7.n5414 0.013
R31240 net7.n5071 net7.n5070 0.013
R31241 net7.n5191 net7.n5190 0.013
R31242 net7.n5348 net7.n5347 0.013
R31243 net7.n5496 net7.n5495 0.013
R31244 net7.n5599 net7.n5598 0.013
R31245 net7.n5779 net7.n5776 0.013
R31246 net7.n5433 net7.n5432 0.013
R31247 net7.n5553 net7.n5552 0.013
R31248 net7.n5710 net7.n5709 0.013
R31249 net7.n5858 net7.n5857 0.013
R31250 net7.n5961 net7.n5960 0.013
R31251 net7.n6141 net7.n6138 0.013
R31252 net7.n5795 net7.n5794 0.013
R31253 net7.n5915 net7.n5914 0.013
R31254 net7.n6072 net7.n6071 0.013
R31255 net7.n6220 net7.n6219 0.013
R31256 net7.n6323 net7.n6322 0.013
R31257 net7.n6503 net7.n6500 0.013
R31258 net7.n6157 net7.n6156 0.013
R31259 net7.n6277 net7.n6276 0.013
R31260 net7.n6434 net7.n6433 0.013
R31261 net7.n6582 net7.n6581 0.013
R31262 net7.n6685 net7.n6684 0.013
R31263 net7.n6865 net7.n6862 0.013
R31264 net7.n6519 net7.n6518 0.013
R31265 net7.n6639 net7.n6638 0.013
R31266 net7.n6796 net7.n6795 0.013
R31267 net7.n6944 net7.n6943 0.013
R31268 net7.n7047 net7.n7046 0.013
R31269 net7.n7227 net7.n7224 0.013
R31270 net7.n6881 net7.n6880 0.013
R31271 net7.n7001 net7.n7000 0.013
R31272 net7.n7158 net7.n7157 0.013
R31273 net7.n3591 net7.n3590 0.011
R31274 net7.n3561 net7.n3560 0.011
R31275 net7.n3396 net7.n3395 0.011
R31276 net7.n3288 net7.n3287 0.011
R31277 net7.n3229 net7.n3228 0.011
R31278 net7.n3199 net7.n3198 0.011
R31279 net7.n3034 net7.n3033 0.011
R31280 net7.n2926 net7.n2925 0.011
R31281 net7.n2867 net7.n2866 0.011
R31282 net7.n2837 net7.n2836 0.011
R31283 net7.n2672 net7.n2671 0.011
R31284 net7.n2564 net7.n2563 0.011
R31285 net7.n2505 net7.n2504 0.011
R31286 net7.n2475 net7.n2474 0.011
R31287 net7.n2310 net7.n2309 0.011
R31288 net7.n2202 net7.n2201 0.011
R31289 net7.n2143 net7.n2142 0.011
R31290 net7.n2113 net7.n2112 0.011
R31291 net7.n1948 net7.n1947 0.011
R31292 net7.n1840 net7.n1839 0.011
R31293 net7.n1781 net7.n1780 0.011
R31294 net7.n1751 net7.n1750 0.011
R31295 net7.n1586 net7.n1585 0.011
R31296 net7.n1478 net7.n1477 0.011
R31297 net7.n1419 net7.n1418 0.011
R31298 net7.n1389 net7.n1388 0.011
R31299 net7.n1224 net7.n1223 0.011
R31300 net7.n1116 net7.n1115 0.011
R31301 net7.n1057 net7.n1056 0.011
R31302 net7.n1027 net7.n1026 0.011
R31303 net7.n862 net7.n861 0.011
R31304 net7.n754 net7.n753 0.011
R31305 net7.n695 net7.n694 0.011
R31306 net7.n665 net7.n664 0.011
R31307 net7.n500 net7.n499 0.011
R31308 net7.n392 net7.n391 0.011
R31309 net7.n334 net7.n333 0.011
R31310 net7.n304 net7.n303 0.011
R31311 net7.n139 net7.n138 0.011
R31312 net7.n31 net7.n30 0.011
R31313 net7.n3677 net7.n3676 0.011
R31314 net7.n3653 net7.n3652 0.011
R31315 net7.n3921 net7.n3920 0.011
R31316 net7.n3955 net7.n3954 0.011
R31317 net7.n4038 net7.n4037 0.011
R31318 net7.n4014 net7.n4013 0.011
R31319 net7.n4282 net7.n4281 0.011
R31320 net7.n4316 net7.n4315 0.011
R31321 net7.n4400 net7.n4399 0.011
R31322 net7.n4376 net7.n4375 0.011
R31323 net7.n4644 net7.n4643 0.011
R31324 net7.n4678 net7.n4677 0.011
R31325 net7.n4762 net7.n4761 0.011
R31326 net7.n4738 net7.n4737 0.011
R31327 net7.n5006 net7.n5005 0.011
R31328 net7.n5040 net7.n5039 0.011
R31329 net7.n5124 net7.n5123 0.011
R31330 net7.n5100 net7.n5099 0.011
R31331 net7.n5368 net7.n5367 0.011
R31332 net7.n5402 net7.n5401 0.011
R31333 net7.n5486 net7.n5485 0.011
R31334 net7.n5462 net7.n5461 0.011
R31335 net7.n5730 net7.n5729 0.011
R31336 net7.n5764 net7.n5763 0.011
R31337 net7.n5848 net7.n5847 0.011
R31338 net7.n5824 net7.n5823 0.011
R31339 net7.n6092 net7.n6091 0.011
R31340 net7.n6126 net7.n6125 0.011
R31341 net7.n6210 net7.n6209 0.011
R31342 net7.n6186 net7.n6185 0.011
R31343 net7.n6454 net7.n6453 0.011
R31344 net7.n6488 net7.n6487 0.011
R31345 net7.n6572 net7.n6571 0.011
R31346 net7.n6548 net7.n6547 0.011
R31347 net7.n6816 net7.n6815 0.011
R31348 net7.n6850 net7.n6849 0.011
R31349 net7.n6934 net7.n6933 0.011
R31350 net7.n6910 net7.n6909 0.011
R31351 net7.n7178 net7.n7177 0.011
R31352 net7.n7212 net7.n7211 0.011
R31353 net7.n3599 net7.n3597 0.009
R31354 net7.n3571 net7.n3570 0.009
R31355 net7.n3345 net7.n3344 0.009
R31356 net7.n3275 net7.n3274 0.009
R31357 net7.n3306 net7.n3305 0.009
R31358 net7.n3616 net7.n3615 0.009
R31359 net7.n3474 net7.n3473 0.009
R31360 net7.n3457 net7.n3456 0.009
R31361 net7.n3349 net7.n3337 0.009
R31362 net7.n3334 net7.n3333 0.009
R31363 net7.n3265 net7.n3264 0.009
R31364 net7.n3507 net7.n3502 0.009
R31365 net7.n3501 net7.n3500 0.009
R31366 net7.n3496 net7.n3491 0.009
R31367 net7.n3490 net7.n3489 0.009
R31368 net7.n3465 net7.n3460 0.009
R31369 net7.n3459 net7.n3458 0.009
R31370 net7.n3454 net7.n3449 0.009
R31371 net7.n3448 net7.n3447 0.009
R31372 net7.n3421 net7.n3371 0.009
R31373 net7.n3370 net7.n3369 0.009
R31374 net7.n3365 net7.n3360 0.009
R31375 net7.n3359 net7.n3358 0.009
R31376 net7.n3326 net7.n3321 0.009
R31377 net7.n3320 net7.n3319 0.009
R31378 net7.n3315 net7.n3314 0.009
R31379 net7.n3313 net7.n3312 0.009
R31380 net7.n3237 net7.n3235 0.009
R31381 net7.n3209 net7.n3208 0.009
R31382 net7.n2983 net7.n2982 0.009
R31383 net7.n2913 net7.n2912 0.009
R31384 net7.n2944 net7.n2943 0.009
R31385 net7.n3254 net7.n3253 0.009
R31386 net7.n3112 net7.n3111 0.009
R31387 net7.n3095 net7.n3094 0.009
R31388 net7.n2987 net7.n2975 0.009
R31389 net7.n2972 net7.n2971 0.009
R31390 net7.n2903 net7.n2902 0.009
R31391 net7.n3145 net7.n3140 0.009
R31392 net7.n3139 net7.n3138 0.009
R31393 net7.n3134 net7.n3129 0.009
R31394 net7.n3128 net7.n3127 0.009
R31395 net7.n3103 net7.n3098 0.009
R31396 net7.n3097 net7.n3096 0.009
R31397 net7.n3092 net7.n3087 0.009
R31398 net7.n3086 net7.n3085 0.009
R31399 net7.n3059 net7.n3009 0.009
R31400 net7.n3008 net7.n3007 0.009
R31401 net7.n3003 net7.n2998 0.009
R31402 net7.n2997 net7.n2996 0.009
R31403 net7.n2964 net7.n2959 0.009
R31404 net7.n2958 net7.n2957 0.009
R31405 net7.n2953 net7.n2952 0.009
R31406 net7.n2951 net7.n2950 0.009
R31407 net7.n2875 net7.n2873 0.009
R31408 net7.n2847 net7.n2846 0.009
R31409 net7.n2621 net7.n2620 0.009
R31410 net7.n2551 net7.n2550 0.009
R31411 net7.n2582 net7.n2581 0.009
R31412 net7.n2892 net7.n2891 0.009
R31413 net7.n2750 net7.n2749 0.009
R31414 net7.n2733 net7.n2732 0.009
R31415 net7.n2625 net7.n2613 0.009
R31416 net7.n2610 net7.n2609 0.009
R31417 net7.n2541 net7.n2540 0.009
R31418 net7.n2783 net7.n2778 0.009
R31419 net7.n2777 net7.n2776 0.009
R31420 net7.n2772 net7.n2767 0.009
R31421 net7.n2766 net7.n2765 0.009
R31422 net7.n2741 net7.n2736 0.009
R31423 net7.n2735 net7.n2734 0.009
R31424 net7.n2730 net7.n2725 0.009
R31425 net7.n2724 net7.n2723 0.009
R31426 net7.n2697 net7.n2647 0.009
R31427 net7.n2646 net7.n2645 0.009
R31428 net7.n2641 net7.n2636 0.009
R31429 net7.n2635 net7.n2634 0.009
R31430 net7.n2602 net7.n2597 0.009
R31431 net7.n2596 net7.n2595 0.009
R31432 net7.n2591 net7.n2590 0.009
R31433 net7.n2589 net7.n2588 0.009
R31434 net7.n2513 net7.n2511 0.009
R31435 net7.n2485 net7.n2484 0.009
R31436 net7.n2259 net7.n2258 0.009
R31437 net7.n2189 net7.n2188 0.009
R31438 net7.n2220 net7.n2219 0.009
R31439 net7.n2530 net7.n2529 0.009
R31440 net7.n2388 net7.n2387 0.009
R31441 net7.n2371 net7.n2370 0.009
R31442 net7.n2263 net7.n2251 0.009
R31443 net7.n2248 net7.n2247 0.009
R31444 net7.n2179 net7.n2178 0.009
R31445 net7.n2421 net7.n2416 0.009
R31446 net7.n2415 net7.n2414 0.009
R31447 net7.n2410 net7.n2405 0.009
R31448 net7.n2404 net7.n2403 0.009
R31449 net7.n2379 net7.n2374 0.009
R31450 net7.n2373 net7.n2372 0.009
R31451 net7.n2368 net7.n2363 0.009
R31452 net7.n2362 net7.n2361 0.009
R31453 net7.n2335 net7.n2285 0.009
R31454 net7.n2284 net7.n2283 0.009
R31455 net7.n2279 net7.n2274 0.009
R31456 net7.n2273 net7.n2272 0.009
R31457 net7.n2240 net7.n2235 0.009
R31458 net7.n2234 net7.n2233 0.009
R31459 net7.n2229 net7.n2228 0.009
R31460 net7.n2227 net7.n2226 0.009
R31461 net7.n2151 net7.n2149 0.009
R31462 net7.n2123 net7.n2122 0.009
R31463 net7.n1897 net7.n1896 0.009
R31464 net7.n1827 net7.n1826 0.009
R31465 net7.n1858 net7.n1857 0.009
R31466 net7.n2168 net7.n2167 0.009
R31467 net7.n2026 net7.n2025 0.009
R31468 net7.n2009 net7.n2008 0.009
R31469 net7.n1901 net7.n1889 0.009
R31470 net7.n1886 net7.n1885 0.009
R31471 net7.n1817 net7.n1816 0.009
R31472 net7.n2059 net7.n2054 0.009
R31473 net7.n2053 net7.n2052 0.009
R31474 net7.n2048 net7.n2043 0.009
R31475 net7.n2042 net7.n2041 0.009
R31476 net7.n2017 net7.n2012 0.009
R31477 net7.n2011 net7.n2010 0.009
R31478 net7.n2006 net7.n2001 0.009
R31479 net7.n2000 net7.n1999 0.009
R31480 net7.n1973 net7.n1923 0.009
R31481 net7.n1922 net7.n1921 0.009
R31482 net7.n1917 net7.n1912 0.009
R31483 net7.n1911 net7.n1910 0.009
R31484 net7.n1878 net7.n1873 0.009
R31485 net7.n1872 net7.n1871 0.009
R31486 net7.n1867 net7.n1866 0.009
R31487 net7.n1865 net7.n1864 0.009
R31488 net7.n1789 net7.n1787 0.009
R31489 net7.n1761 net7.n1760 0.009
R31490 net7.n1535 net7.n1534 0.009
R31491 net7.n1465 net7.n1464 0.009
R31492 net7.n1496 net7.n1495 0.009
R31493 net7.n1806 net7.n1805 0.009
R31494 net7.n1664 net7.n1663 0.009
R31495 net7.n1647 net7.n1646 0.009
R31496 net7.n1539 net7.n1527 0.009
R31497 net7.n1524 net7.n1523 0.009
R31498 net7.n1455 net7.n1454 0.009
R31499 net7.n1697 net7.n1692 0.009
R31500 net7.n1691 net7.n1690 0.009
R31501 net7.n1686 net7.n1681 0.009
R31502 net7.n1680 net7.n1679 0.009
R31503 net7.n1655 net7.n1650 0.009
R31504 net7.n1649 net7.n1648 0.009
R31505 net7.n1644 net7.n1639 0.009
R31506 net7.n1638 net7.n1637 0.009
R31507 net7.n1611 net7.n1561 0.009
R31508 net7.n1560 net7.n1559 0.009
R31509 net7.n1555 net7.n1550 0.009
R31510 net7.n1549 net7.n1548 0.009
R31511 net7.n1516 net7.n1511 0.009
R31512 net7.n1510 net7.n1509 0.009
R31513 net7.n1505 net7.n1504 0.009
R31514 net7.n1503 net7.n1502 0.009
R31515 net7.n1427 net7.n1425 0.009
R31516 net7.n1399 net7.n1398 0.009
R31517 net7.n1173 net7.n1172 0.009
R31518 net7.n1103 net7.n1102 0.009
R31519 net7.n1134 net7.n1133 0.009
R31520 net7.n1444 net7.n1443 0.009
R31521 net7.n1302 net7.n1301 0.009
R31522 net7.n1285 net7.n1284 0.009
R31523 net7.n1177 net7.n1165 0.009
R31524 net7.n1162 net7.n1161 0.009
R31525 net7.n1093 net7.n1092 0.009
R31526 net7.n1335 net7.n1330 0.009
R31527 net7.n1329 net7.n1328 0.009
R31528 net7.n1324 net7.n1319 0.009
R31529 net7.n1318 net7.n1317 0.009
R31530 net7.n1293 net7.n1288 0.009
R31531 net7.n1287 net7.n1286 0.009
R31532 net7.n1282 net7.n1277 0.009
R31533 net7.n1276 net7.n1275 0.009
R31534 net7.n1249 net7.n1199 0.009
R31535 net7.n1198 net7.n1197 0.009
R31536 net7.n1193 net7.n1188 0.009
R31537 net7.n1187 net7.n1186 0.009
R31538 net7.n1154 net7.n1149 0.009
R31539 net7.n1148 net7.n1147 0.009
R31540 net7.n1143 net7.n1142 0.009
R31541 net7.n1141 net7.n1140 0.009
R31542 net7.n1065 net7.n1063 0.009
R31543 net7.n1037 net7.n1036 0.009
R31544 net7.n811 net7.n810 0.009
R31545 net7.n741 net7.n740 0.009
R31546 net7.n772 net7.n771 0.009
R31547 net7.n1082 net7.n1081 0.009
R31548 net7.n940 net7.n939 0.009
R31549 net7.n923 net7.n922 0.009
R31550 net7.n815 net7.n803 0.009
R31551 net7.n800 net7.n799 0.009
R31552 net7.n731 net7.n730 0.009
R31553 net7.n973 net7.n968 0.009
R31554 net7.n967 net7.n966 0.009
R31555 net7.n962 net7.n957 0.009
R31556 net7.n956 net7.n955 0.009
R31557 net7.n931 net7.n926 0.009
R31558 net7.n925 net7.n924 0.009
R31559 net7.n920 net7.n915 0.009
R31560 net7.n914 net7.n913 0.009
R31561 net7.n887 net7.n837 0.009
R31562 net7.n836 net7.n835 0.009
R31563 net7.n831 net7.n826 0.009
R31564 net7.n825 net7.n824 0.009
R31565 net7.n792 net7.n787 0.009
R31566 net7.n786 net7.n785 0.009
R31567 net7.n781 net7.n780 0.009
R31568 net7.n779 net7.n778 0.009
R31569 net7.n703 net7.n701 0.009
R31570 net7.n675 net7.n674 0.009
R31571 net7.n449 net7.n448 0.009
R31572 net7.n379 net7.n378 0.009
R31573 net7.n410 net7.n409 0.009
R31574 net7.n720 net7.n719 0.009
R31575 net7.n578 net7.n577 0.009
R31576 net7.n561 net7.n560 0.009
R31577 net7.n453 net7.n441 0.009
R31578 net7.n438 net7.n437 0.009
R31579 net7.n369 net7.n368 0.009
R31580 net7.n611 net7.n606 0.009
R31581 net7.n605 net7.n604 0.009
R31582 net7.n600 net7.n595 0.009
R31583 net7.n594 net7.n593 0.009
R31584 net7.n569 net7.n564 0.009
R31585 net7.n563 net7.n562 0.009
R31586 net7.n558 net7.n553 0.009
R31587 net7.n552 net7.n551 0.009
R31588 net7.n525 net7.n475 0.009
R31589 net7.n474 net7.n473 0.009
R31590 net7.n469 net7.n464 0.009
R31591 net7.n463 net7.n462 0.009
R31592 net7.n430 net7.n425 0.009
R31593 net7.n424 net7.n423 0.009
R31594 net7.n419 net7.n418 0.009
R31595 net7.n417 net7.n416 0.009
R31596 net7.n342 net7.n340 0.009
R31597 net7.n314 net7.n313 0.009
R31598 net7.n88 net7.n87 0.009
R31599 net7.n18 net7.n17 0.009
R31600 net7.n49 net7.n48 0.009
R31601 net7.n359 net7.n358 0.009
R31602 net7.n217 net7.n216 0.009
R31603 net7.n200 net7.n199 0.009
R31604 net7.n92 net7.n80 0.009
R31605 net7.n77 net7.n76 0.009
R31606 net7.n8 net7.n7 0.009
R31607 net7.n250 net7.n245 0.009
R31608 net7.n244 net7.n243 0.009
R31609 net7.n239 net7.n234 0.009
R31610 net7.n233 net7.n232 0.009
R31611 net7.n208 net7.n203 0.009
R31612 net7.n202 net7.n201 0.009
R31613 net7.n197 net7.n192 0.009
R31614 net7.n191 net7.n190 0.009
R31615 net7.n164 net7.n114 0.009
R31616 net7.n113 net7.n112 0.009
R31617 net7.n108 net7.n103 0.009
R31618 net7.n102 net7.n101 0.009
R31619 net7.n69 net7.n64 0.009
R31620 net7.n63 net7.n62 0.009
R31621 net7.n58 net7.n57 0.009
R31622 net7.n56 net7.n55 0.009
R31623 net7.n3685 net7.n3683 0.009
R31624 net7.n3660 net7.n3659 0.009
R31625 net7.n3934 net7.n3933 0.009
R31626 net7.n3942 net7.n3941 0.009
R31627 net7.n3973 net7.n3972 0.009
R31628 net7.n3725 net7.n3724 0.009
R31629 net7.n3740 net7.n3739 0.009
R31630 net7.n3868 net7.n3866 0.009
R31631 net7.n3872 net7.n3871 0.009
R31632 net7.n3874 net7.n3873 0.009
R31633 net7.n3906 net7.n3905 0.009
R31634 net7.n3978 net7.n3909 0.009
R31635 net7.n3697 net7.n3696 0.009
R31636 net7.n3699 net7.n3698 0.009
R31637 net7.n3704 net7.n3703 0.009
R31638 net7.n3709 net7.n3705 0.009
R31639 net7.n3735 net7.n3734 0.009
R31640 net7.n3741 net7.n3736 0.009
R31641 net7.n3746 net7.n3745 0.009
R31642 net7.n3752 net7.n3747 0.009
R31643 net7.n3842 net7.n3841 0.009
R31644 net7.n3848 net7.n3843 0.009
R31645 net7.n3853 net7.n3852 0.009
R31646 net7.n3859 net7.n3854 0.009
R31647 net7.n3884 net7.n3883 0.009
R31648 net7.n3890 net7.n3885 0.009
R31649 net7.n3895 net7.n3894 0.009
R31650 net7.n3902 net7.n3896 0.009
R31651 net7.n4046 net7.n4044 0.009
R31652 net7.n4021 net7.n4020 0.009
R31653 net7.n4295 net7.n4294 0.009
R31654 net7.n4303 net7.n4302 0.009
R31655 net7.n4334 net7.n4333 0.009
R31656 net7.n4086 net7.n4085 0.009
R31657 net7.n4101 net7.n4100 0.009
R31658 net7.n4229 net7.n4227 0.009
R31659 net7.n4233 net7.n4232 0.009
R31660 net7.n4235 net7.n4234 0.009
R31661 net7.n4267 net7.n4266 0.009
R31662 net7.n4339 net7.n4270 0.009
R31663 net7.n4058 net7.n4057 0.009
R31664 net7.n4060 net7.n4059 0.009
R31665 net7.n4065 net7.n4064 0.009
R31666 net7.n4070 net7.n4066 0.009
R31667 net7.n4096 net7.n4095 0.009
R31668 net7.n4102 net7.n4097 0.009
R31669 net7.n4107 net7.n4106 0.009
R31670 net7.n4113 net7.n4108 0.009
R31671 net7.n4203 net7.n4202 0.009
R31672 net7.n4209 net7.n4204 0.009
R31673 net7.n4214 net7.n4213 0.009
R31674 net7.n4220 net7.n4215 0.009
R31675 net7.n4245 net7.n4244 0.009
R31676 net7.n4251 net7.n4246 0.009
R31677 net7.n4256 net7.n4255 0.009
R31678 net7.n4263 net7.n4257 0.009
R31679 net7.n4408 net7.n4406 0.009
R31680 net7.n4383 net7.n4382 0.009
R31681 net7.n4657 net7.n4656 0.009
R31682 net7.n4665 net7.n4664 0.009
R31683 net7.n4696 net7.n4695 0.009
R31684 net7.n4448 net7.n4447 0.009
R31685 net7.n4463 net7.n4462 0.009
R31686 net7.n4591 net7.n4589 0.009
R31687 net7.n4595 net7.n4594 0.009
R31688 net7.n4597 net7.n4596 0.009
R31689 net7.n4629 net7.n4628 0.009
R31690 net7.n4701 net7.n4632 0.009
R31691 net7.n4420 net7.n4419 0.009
R31692 net7.n4422 net7.n4421 0.009
R31693 net7.n4427 net7.n4426 0.009
R31694 net7.n4432 net7.n4428 0.009
R31695 net7.n4458 net7.n4457 0.009
R31696 net7.n4464 net7.n4459 0.009
R31697 net7.n4469 net7.n4468 0.009
R31698 net7.n4475 net7.n4470 0.009
R31699 net7.n4565 net7.n4564 0.009
R31700 net7.n4571 net7.n4566 0.009
R31701 net7.n4576 net7.n4575 0.009
R31702 net7.n4582 net7.n4577 0.009
R31703 net7.n4607 net7.n4606 0.009
R31704 net7.n4613 net7.n4608 0.009
R31705 net7.n4618 net7.n4617 0.009
R31706 net7.n4625 net7.n4619 0.009
R31707 net7.n4770 net7.n4768 0.009
R31708 net7.n4745 net7.n4744 0.009
R31709 net7.n5019 net7.n5018 0.009
R31710 net7.n5027 net7.n5026 0.009
R31711 net7.n5058 net7.n5057 0.009
R31712 net7.n4810 net7.n4809 0.009
R31713 net7.n4825 net7.n4824 0.009
R31714 net7.n4953 net7.n4951 0.009
R31715 net7.n4957 net7.n4956 0.009
R31716 net7.n4959 net7.n4958 0.009
R31717 net7.n4991 net7.n4990 0.009
R31718 net7.n5063 net7.n4994 0.009
R31719 net7.n4782 net7.n4781 0.009
R31720 net7.n4784 net7.n4783 0.009
R31721 net7.n4789 net7.n4788 0.009
R31722 net7.n4794 net7.n4790 0.009
R31723 net7.n4820 net7.n4819 0.009
R31724 net7.n4826 net7.n4821 0.009
R31725 net7.n4831 net7.n4830 0.009
R31726 net7.n4837 net7.n4832 0.009
R31727 net7.n4927 net7.n4926 0.009
R31728 net7.n4933 net7.n4928 0.009
R31729 net7.n4938 net7.n4937 0.009
R31730 net7.n4944 net7.n4939 0.009
R31731 net7.n4969 net7.n4968 0.009
R31732 net7.n4975 net7.n4970 0.009
R31733 net7.n4980 net7.n4979 0.009
R31734 net7.n4987 net7.n4981 0.009
R31735 net7.n5132 net7.n5130 0.009
R31736 net7.n5107 net7.n5106 0.009
R31737 net7.n5381 net7.n5380 0.009
R31738 net7.n5389 net7.n5388 0.009
R31739 net7.n5420 net7.n5419 0.009
R31740 net7.n5172 net7.n5171 0.009
R31741 net7.n5187 net7.n5186 0.009
R31742 net7.n5315 net7.n5313 0.009
R31743 net7.n5319 net7.n5318 0.009
R31744 net7.n5321 net7.n5320 0.009
R31745 net7.n5353 net7.n5352 0.009
R31746 net7.n5425 net7.n5356 0.009
R31747 net7.n5144 net7.n5143 0.009
R31748 net7.n5146 net7.n5145 0.009
R31749 net7.n5151 net7.n5150 0.009
R31750 net7.n5156 net7.n5152 0.009
R31751 net7.n5182 net7.n5181 0.009
R31752 net7.n5188 net7.n5183 0.009
R31753 net7.n5193 net7.n5192 0.009
R31754 net7.n5199 net7.n5194 0.009
R31755 net7.n5289 net7.n5288 0.009
R31756 net7.n5295 net7.n5290 0.009
R31757 net7.n5300 net7.n5299 0.009
R31758 net7.n5306 net7.n5301 0.009
R31759 net7.n5331 net7.n5330 0.009
R31760 net7.n5337 net7.n5332 0.009
R31761 net7.n5342 net7.n5341 0.009
R31762 net7.n5349 net7.n5343 0.009
R31763 net7.n5494 net7.n5492 0.009
R31764 net7.n5469 net7.n5468 0.009
R31765 net7.n5743 net7.n5742 0.009
R31766 net7.n5751 net7.n5750 0.009
R31767 net7.n5782 net7.n5781 0.009
R31768 net7.n5534 net7.n5533 0.009
R31769 net7.n5549 net7.n5548 0.009
R31770 net7.n5677 net7.n5675 0.009
R31771 net7.n5681 net7.n5680 0.009
R31772 net7.n5683 net7.n5682 0.009
R31773 net7.n5715 net7.n5714 0.009
R31774 net7.n5787 net7.n5718 0.009
R31775 net7.n5506 net7.n5505 0.009
R31776 net7.n5508 net7.n5507 0.009
R31777 net7.n5513 net7.n5512 0.009
R31778 net7.n5518 net7.n5514 0.009
R31779 net7.n5544 net7.n5543 0.009
R31780 net7.n5550 net7.n5545 0.009
R31781 net7.n5555 net7.n5554 0.009
R31782 net7.n5561 net7.n5556 0.009
R31783 net7.n5651 net7.n5650 0.009
R31784 net7.n5657 net7.n5652 0.009
R31785 net7.n5662 net7.n5661 0.009
R31786 net7.n5668 net7.n5663 0.009
R31787 net7.n5693 net7.n5692 0.009
R31788 net7.n5699 net7.n5694 0.009
R31789 net7.n5704 net7.n5703 0.009
R31790 net7.n5711 net7.n5705 0.009
R31791 net7.n5856 net7.n5854 0.009
R31792 net7.n5831 net7.n5830 0.009
R31793 net7.n6105 net7.n6104 0.009
R31794 net7.n6113 net7.n6112 0.009
R31795 net7.n6144 net7.n6143 0.009
R31796 net7.n5896 net7.n5895 0.009
R31797 net7.n5911 net7.n5910 0.009
R31798 net7.n6039 net7.n6037 0.009
R31799 net7.n6043 net7.n6042 0.009
R31800 net7.n6045 net7.n6044 0.009
R31801 net7.n6077 net7.n6076 0.009
R31802 net7.n6149 net7.n6080 0.009
R31803 net7.n5868 net7.n5867 0.009
R31804 net7.n5870 net7.n5869 0.009
R31805 net7.n5875 net7.n5874 0.009
R31806 net7.n5880 net7.n5876 0.009
R31807 net7.n5906 net7.n5905 0.009
R31808 net7.n5912 net7.n5907 0.009
R31809 net7.n5917 net7.n5916 0.009
R31810 net7.n5923 net7.n5918 0.009
R31811 net7.n6013 net7.n6012 0.009
R31812 net7.n6019 net7.n6014 0.009
R31813 net7.n6024 net7.n6023 0.009
R31814 net7.n6030 net7.n6025 0.009
R31815 net7.n6055 net7.n6054 0.009
R31816 net7.n6061 net7.n6056 0.009
R31817 net7.n6066 net7.n6065 0.009
R31818 net7.n6073 net7.n6067 0.009
R31819 net7.n6218 net7.n6216 0.009
R31820 net7.n6193 net7.n6192 0.009
R31821 net7.n6467 net7.n6466 0.009
R31822 net7.n6475 net7.n6474 0.009
R31823 net7.n6506 net7.n6505 0.009
R31824 net7.n6258 net7.n6257 0.009
R31825 net7.n6273 net7.n6272 0.009
R31826 net7.n6401 net7.n6399 0.009
R31827 net7.n6405 net7.n6404 0.009
R31828 net7.n6407 net7.n6406 0.009
R31829 net7.n6439 net7.n6438 0.009
R31830 net7.n6511 net7.n6442 0.009
R31831 net7.n6230 net7.n6229 0.009
R31832 net7.n6232 net7.n6231 0.009
R31833 net7.n6237 net7.n6236 0.009
R31834 net7.n6242 net7.n6238 0.009
R31835 net7.n6268 net7.n6267 0.009
R31836 net7.n6274 net7.n6269 0.009
R31837 net7.n6279 net7.n6278 0.009
R31838 net7.n6285 net7.n6280 0.009
R31839 net7.n6375 net7.n6374 0.009
R31840 net7.n6381 net7.n6376 0.009
R31841 net7.n6386 net7.n6385 0.009
R31842 net7.n6392 net7.n6387 0.009
R31843 net7.n6417 net7.n6416 0.009
R31844 net7.n6423 net7.n6418 0.009
R31845 net7.n6428 net7.n6427 0.009
R31846 net7.n6435 net7.n6429 0.009
R31847 net7.n6580 net7.n6578 0.009
R31848 net7.n6555 net7.n6554 0.009
R31849 net7.n6829 net7.n6828 0.009
R31850 net7.n6837 net7.n6836 0.009
R31851 net7.n6868 net7.n6867 0.009
R31852 net7.n6620 net7.n6619 0.009
R31853 net7.n6635 net7.n6634 0.009
R31854 net7.n6763 net7.n6761 0.009
R31855 net7.n6767 net7.n6766 0.009
R31856 net7.n6769 net7.n6768 0.009
R31857 net7.n6801 net7.n6800 0.009
R31858 net7.n6873 net7.n6804 0.009
R31859 net7.n6592 net7.n6591 0.009
R31860 net7.n6594 net7.n6593 0.009
R31861 net7.n6599 net7.n6598 0.009
R31862 net7.n6604 net7.n6600 0.009
R31863 net7.n6630 net7.n6629 0.009
R31864 net7.n6636 net7.n6631 0.009
R31865 net7.n6641 net7.n6640 0.009
R31866 net7.n6647 net7.n6642 0.009
R31867 net7.n6737 net7.n6736 0.009
R31868 net7.n6743 net7.n6738 0.009
R31869 net7.n6748 net7.n6747 0.009
R31870 net7.n6754 net7.n6749 0.009
R31871 net7.n6779 net7.n6778 0.009
R31872 net7.n6785 net7.n6780 0.009
R31873 net7.n6790 net7.n6789 0.009
R31874 net7.n6797 net7.n6791 0.009
R31875 net7.n6942 net7.n6940 0.009
R31876 net7.n6917 net7.n6916 0.009
R31877 net7.n7191 net7.n7190 0.009
R31878 net7.n7199 net7.n7198 0.009
R31879 net7.n7230 net7.n7229 0.009
R31880 net7.n6982 net7.n6981 0.009
R31881 net7.n6997 net7.n6996 0.009
R31882 net7.n7125 net7.n7123 0.009
R31883 net7.n7129 net7.n7128 0.009
R31884 net7.n7131 net7.n7130 0.009
R31885 net7.n7163 net7.n7162 0.009
R31886 net7.n7235 net7.n7166 0.009
R31887 net7.n6954 net7.n6953 0.009
R31888 net7.n6956 net7.n6955 0.009
R31889 net7.n6961 net7.n6960 0.009
R31890 net7.n6966 net7.n6962 0.009
R31891 net7.n6992 net7.n6991 0.009
R31892 net7.n6998 net7.n6993 0.009
R31893 net7.n7003 net7.n7002 0.009
R31894 net7.n7009 net7.n7004 0.009
R31895 net7.n7099 net7.n7098 0.009
R31896 net7.n7105 net7.n7100 0.009
R31897 net7.n7110 net7.n7109 0.009
R31898 net7.n7116 net7.n7111 0.009
R31899 net7.n7141 net7.n7140 0.009
R31900 net7.n7147 net7.n7142 0.009
R31901 net7.n7152 net7.n7151 0.009
R31902 net7.n7159 net7.n7153 0.009
R31903 net7.n3606 net7.n3605 0.007
R31904 net7.n3596 net7.n3595 0.007
R31905 net7.n3576 net7.n3575 0.007
R31906 net7.n3570 net7.n3569 0.007
R31907 net7.n3547 net7.n3546 0.007
R31908 net7.n3375 net7.n3374 0.007
R31909 net7.n3384 net7.n3383 0.007
R31910 net7.n3406 net7.n3405 0.007
R31911 net7.n3401 net7.n3400 0.007
R31912 net7.n3399 net7.n3398 0.007
R31913 net7.n3395 net7.n3394 0.007
R31914 net7.n3346 net7.n3345 0.007
R31915 net7.n3299 net7.n3297 0.007
R31916 net7.n3612 net7.n3611 0.007
R31917 net7.n3499 net7.n3498 0.007
R31918 net7.n3482 net7.n3477 0.007
R31919 net7.n3481 net7.n3480 0.007
R31920 net7.n3433 net7.n3432 0.007
R31921 net7.n3435 net7.n3434 0.007
R31922 net7.n3428 net7.n3427 0.007
R31923 net7.n3364 net7.n3361 0.007
R31924 net7.n3357 net7.n3356 0.007
R31925 net7.n3355 net7.n3354 0.007
R31926 net7.n3244 net7.n3243 0.007
R31927 net7.n3234 net7.n3233 0.007
R31928 net7.n3214 net7.n3213 0.007
R31929 net7.n3208 net7.n3207 0.007
R31930 net7.n3185 net7.n3184 0.007
R31931 net7.n3013 net7.n3012 0.007
R31932 net7.n3022 net7.n3021 0.007
R31933 net7.n3044 net7.n3043 0.007
R31934 net7.n3039 net7.n3038 0.007
R31935 net7.n3037 net7.n3036 0.007
R31936 net7.n3033 net7.n3032 0.007
R31937 net7.n2984 net7.n2983 0.007
R31938 net7.n2937 net7.n2935 0.007
R31939 net7.n3250 net7.n3249 0.007
R31940 net7.n3137 net7.n3136 0.007
R31941 net7.n3120 net7.n3115 0.007
R31942 net7.n3119 net7.n3118 0.007
R31943 net7.n3071 net7.n3070 0.007
R31944 net7.n3073 net7.n3072 0.007
R31945 net7.n3066 net7.n3065 0.007
R31946 net7.n3002 net7.n2999 0.007
R31947 net7.n2995 net7.n2994 0.007
R31948 net7.n2993 net7.n2992 0.007
R31949 net7.n2882 net7.n2881 0.007
R31950 net7.n2872 net7.n2871 0.007
R31951 net7.n2852 net7.n2851 0.007
R31952 net7.n2846 net7.n2845 0.007
R31953 net7.n2823 net7.n2822 0.007
R31954 net7.n2651 net7.n2650 0.007
R31955 net7.n2660 net7.n2659 0.007
R31956 net7.n2682 net7.n2681 0.007
R31957 net7.n2677 net7.n2676 0.007
R31958 net7.n2675 net7.n2674 0.007
R31959 net7.n2671 net7.n2670 0.007
R31960 net7.n2622 net7.n2621 0.007
R31961 net7.n2575 net7.n2573 0.007
R31962 net7.n2888 net7.n2887 0.007
R31963 net7.n2775 net7.n2774 0.007
R31964 net7.n2758 net7.n2753 0.007
R31965 net7.n2757 net7.n2756 0.007
R31966 net7.n2709 net7.n2708 0.007
R31967 net7.n2711 net7.n2710 0.007
R31968 net7.n2704 net7.n2703 0.007
R31969 net7.n2640 net7.n2637 0.007
R31970 net7.n2633 net7.n2632 0.007
R31971 net7.n2631 net7.n2630 0.007
R31972 net7.n2520 net7.n2519 0.007
R31973 net7.n2510 net7.n2509 0.007
R31974 net7.n2490 net7.n2489 0.007
R31975 net7.n2484 net7.n2483 0.007
R31976 net7.n2461 net7.n2460 0.007
R31977 net7.n2289 net7.n2288 0.007
R31978 net7.n2298 net7.n2297 0.007
R31979 net7.n2320 net7.n2319 0.007
R31980 net7.n2315 net7.n2314 0.007
R31981 net7.n2313 net7.n2312 0.007
R31982 net7.n2309 net7.n2308 0.007
R31983 net7.n2260 net7.n2259 0.007
R31984 net7.n2213 net7.n2211 0.007
R31985 net7.n2526 net7.n2525 0.007
R31986 net7.n2413 net7.n2412 0.007
R31987 net7.n2396 net7.n2391 0.007
R31988 net7.n2395 net7.n2394 0.007
R31989 net7.n2347 net7.n2346 0.007
R31990 net7.n2349 net7.n2348 0.007
R31991 net7.n2342 net7.n2341 0.007
R31992 net7.n2278 net7.n2275 0.007
R31993 net7.n2271 net7.n2270 0.007
R31994 net7.n2269 net7.n2268 0.007
R31995 net7.n2158 net7.n2157 0.007
R31996 net7.n2148 net7.n2147 0.007
R31997 net7.n2128 net7.n2127 0.007
R31998 net7.n2122 net7.n2121 0.007
R31999 net7.n2099 net7.n2098 0.007
R32000 net7.n1927 net7.n1926 0.007
R32001 net7.n1936 net7.n1935 0.007
R32002 net7.n1958 net7.n1957 0.007
R32003 net7.n1953 net7.n1952 0.007
R32004 net7.n1951 net7.n1950 0.007
R32005 net7.n1947 net7.n1946 0.007
R32006 net7.n1898 net7.n1897 0.007
R32007 net7.n1851 net7.n1849 0.007
R32008 net7.n2164 net7.n2163 0.007
R32009 net7.n2051 net7.n2050 0.007
R32010 net7.n2034 net7.n2029 0.007
R32011 net7.n2033 net7.n2032 0.007
R32012 net7.n1985 net7.n1984 0.007
R32013 net7.n1987 net7.n1986 0.007
R32014 net7.n1980 net7.n1979 0.007
R32015 net7.n1916 net7.n1913 0.007
R32016 net7.n1909 net7.n1908 0.007
R32017 net7.n1907 net7.n1906 0.007
R32018 net7.n1796 net7.n1795 0.007
R32019 net7.n1786 net7.n1785 0.007
R32020 net7.n1766 net7.n1765 0.007
R32021 net7.n1760 net7.n1759 0.007
R32022 net7.n1737 net7.n1736 0.007
R32023 net7.n1565 net7.n1564 0.007
R32024 net7.n1574 net7.n1573 0.007
R32025 net7.n1596 net7.n1595 0.007
R32026 net7.n1591 net7.n1590 0.007
R32027 net7.n1589 net7.n1588 0.007
R32028 net7.n1585 net7.n1584 0.007
R32029 net7.n1536 net7.n1535 0.007
R32030 net7.n1489 net7.n1487 0.007
R32031 net7.n1802 net7.n1801 0.007
R32032 net7.n1689 net7.n1688 0.007
R32033 net7.n1672 net7.n1667 0.007
R32034 net7.n1671 net7.n1670 0.007
R32035 net7.n1623 net7.n1622 0.007
R32036 net7.n1625 net7.n1624 0.007
R32037 net7.n1618 net7.n1617 0.007
R32038 net7.n1554 net7.n1551 0.007
R32039 net7.n1547 net7.n1546 0.007
R32040 net7.n1545 net7.n1544 0.007
R32041 net7.n1434 net7.n1433 0.007
R32042 net7.n1424 net7.n1423 0.007
R32043 net7.n1404 net7.n1403 0.007
R32044 net7.n1398 net7.n1397 0.007
R32045 net7.n1375 net7.n1374 0.007
R32046 net7.n1203 net7.n1202 0.007
R32047 net7.n1212 net7.n1211 0.007
R32048 net7.n1234 net7.n1233 0.007
R32049 net7.n1229 net7.n1228 0.007
R32050 net7.n1227 net7.n1226 0.007
R32051 net7.n1223 net7.n1222 0.007
R32052 net7.n1174 net7.n1173 0.007
R32053 net7.n1127 net7.n1125 0.007
R32054 net7.n1440 net7.n1439 0.007
R32055 net7.n1327 net7.n1326 0.007
R32056 net7.n1310 net7.n1305 0.007
R32057 net7.n1309 net7.n1308 0.007
R32058 net7.n1261 net7.n1260 0.007
R32059 net7.n1263 net7.n1262 0.007
R32060 net7.n1256 net7.n1255 0.007
R32061 net7.n1192 net7.n1189 0.007
R32062 net7.n1185 net7.n1184 0.007
R32063 net7.n1183 net7.n1182 0.007
R32064 net7.n1072 net7.n1071 0.007
R32065 net7.n1062 net7.n1061 0.007
R32066 net7.n1042 net7.n1041 0.007
R32067 net7.n1036 net7.n1035 0.007
R32068 net7.n1013 net7.n1012 0.007
R32069 net7.n841 net7.n840 0.007
R32070 net7.n850 net7.n849 0.007
R32071 net7.n872 net7.n871 0.007
R32072 net7.n867 net7.n866 0.007
R32073 net7.n865 net7.n864 0.007
R32074 net7.n861 net7.n860 0.007
R32075 net7.n812 net7.n811 0.007
R32076 net7.n765 net7.n763 0.007
R32077 net7.n1078 net7.n1077 0.007
R32078 net7.n965 net7.n964 0.007
R32079 net7.n948 net7.n943 0.007
R32080 net7.n947 net7.n946 0.007
R32081 net7.n899 net7.n898 0.007
R32082 net7.n901 net7.n900 0.007
R32083 net7.n894 net7.n893 0.007
R32084 net7.n830 net7.n827 0.007
R32085 net7.n823 net7.n822 0.007
R32086 net7.n821 net7.n820 0.007
R32087 net7.n710 net7.n709 0.007
R32088 net7.n700 net7.n699 0.007
R32089 net7.n680 net7.n679 0.007
R32090 net7.n674 net7.n673 0.007
R32091 net7.n651 net7.n650 0.007
R32092 net7.n479 net7.n478 0.007
R32093 net7.n488 net7.n487 0.007
R32094 net7.n510 net7.n509 0.007
R32095 net7.n505 net7.n504 0.007
R32096 net7.n503 net7.n502 0.007
R32097 net7.n499 net7.n498 0.007
R32098 net7.n450 net7.n449 0.007
R32099 net7.n403 net7.n401 0.007
R32100 net7.n716 net7.n715 0.007
R32101 net7.n603 net7.n602 0.007
R32102 net7.n586 net7.n581 0.007
R32103 net7.n585 net7.n584 0.007
R32104 net7.n537 net7.n536 0.007
R32105 net7.n539 net7.n538 0.007
R32106 net7.n532 net7.n531 0.007
R32107 net7.n468 net7.n465 0.007
R32108 net7.n461 net7.n460 0.007
R32109 net7.n459 net7.n458 0.007
R32110 net7.n349 net7.n348 0.007
R32111 net7.n339 net7.n338 0.007
R32112 net7.n319 net7.n318 0.007
R32113 net7.n313 net7.n312 0.007
R32114 net7.n290 net7.n289 0.007
R32115 net7.n118 net7.n117 0.007
R32116 net7.n127 net7.n126 0.007
R32117 net7.n149 net7.n148 0.007
R32118 net7.n144 net7.n143 0.007
R32119 net7.n142 net7.n141 0.007
R32120 net7.n138 net7.n137 0.007
R32121 net7.n89 net7.n88 0.007
R32122 net7.n42 net7.n40 0.007
R32123 net7.n355 net7.n354 0.007
R32124 net7.n242 net7.n241 0.007
R32125 net7.n225 net7.n220 0.007
R32126 net7.n224 net7.n223 0.007
R32127 net7.n176 net7.n175 0.007
R32128 net7.n178 net7.n177 0.007
R32129 net7.n171 net7.n170 0.007
R32130 net7.n107 net7.n104 0.007
R32131 net7.n100 net7.n99 0.007
R32132 net7.n98 net7.n97 0.007
R32133 net7.n3690 net7.n3689 0.007
R32134 net7.n3682 net7.n3681 0.007
R32135 net7.n3665 net7.n3664 0.007
R32136 net7.n3659 net7.n3658 0.007
R32137 net7.n3784 net7.n3783 0.007
R32138 net7.n3814 net7.n3813 0.007
R32139 net7.n3823 net7.n3822 0.007
R32140 net7.n3830 net7.n3829 0.007
R32141 net7.n3914 net7.n3913 0.007
R32142 net7.n3918 net7.n3915 0.007
R32143 net7.n3926 net7.n3921 0.007
R32144 net7.n3933 net7.n3932 0.007
R32145 net7.n3966 net7.n3964 0.007
R32146 net7.n3626 net7.n3625 0.007
R32147 net7.n3620 net7.n3619 0.007
R32148 net7.n3716 net7.n3715 0.007
R32149 net7.n3719 net7.n3718 0.007
R32150 net7.n3760 net7.n3759 0.007
R32151 net7.n3766 net7.n3765 0.007
R32152 net7.n3769 net7.n3768 0.007
R32153 net7.n3851 net7.n3850 0.007
R32154 net7.n3858 net7.n3857 0.007
R32155 net7.n3863 net7.n3862 0.007
R32156 net7.n4051 net7.n4050 0.007
R32157 net7.n4043 net7.n4042 0.007
R32158 net7.n4026 net7.n4025 0.007
R32159 net7.n4020 net7.n4019 0.007
R32160 net7.n4145 net7.n4144 0.007
R32161 net7.n4175 net7.n4174 0.007
R32162 net7.n4184 net7.n4183 0.007
R32163 net7.n4191 net7.n4190 0.007
R32164 net7.n4275 net7.n4274 0.007
R32165 net7.n4279 net7.n4276 0.007
R32166 net7.n4287 net7.n4282 0.007
R32167 net7.n4294 net7.n4293 0.007
R32168 net7.n4327 net7.n4325 0.007
R32169 net7.n3987 net7.n3986 0.007
R32170 net7.n3981 net7.n3980 0.007
R32171 net7.n4077 net7.n4076 0.007
R32172 net7.n4080 net7.n4079 0.007
R32173 net7.n4121 net7.n4120 0.007
R32174 net7.n4127 net7.n4126 0.007
R32175 net7.n4130 net7.n4129 0.007
R32176 net7.n4212 net7.n4211 0.007
R32177 net7.n4219 net7.n4218 0.007
R32178 net7.n4224 net7.n4223 0.007
R32179 net7.n4413 net7.n4412 0.007
R32180 net7.n4405 net7.n4404 0.007
R32181 net7.n4388 net7.n4387 0.007
R32182 net7.n4382 net7.n4381 0.007
R32183 net7.n4507 net7.n4506 0.007
R32184 net7.n4537 net7.n4536 0.007
R32185 net7.n4546 net7.n4545 0.007
R32186 net7.n4553 net7.n4552 0.007
R32187 net7.n4637 net7.n4636 0.007
R32188 net7.n4641 net7.n4638 0.007
R32189 net7.n4649 net7.n4644 0.007
R32190 net7.n4656 net7.n4655 0.007
R32191 net7.n4689 net7.n4687 0.007
R32192 net7.n4349 net7.n4348 0.007
R32193 net7.n4343 net7.n4342 0.007
R32194 net7.n4439 net7.n4438 0.007
R32195 net7.n4442 net7.n4441 0.007
R32196 net7.n4483 net7.n4482 0.007
R32197 net7.n4489 net7.n4488 0.007
R32198 net7.n4492 net7.n4491 0.007
R32199 net7.n4574 net7.n4573 0.007
R32200 net7.n4581 net7.n4580 0.007
R32201 net7.n4586 net7.n4585 0.007
R32202 net7.n4775 net7.n4774 0.007
R32203 net7.n4767 net7.n4766 0.007
R32204 net7.n4750 net7.n4749 0.007
R32205 net7.n4744 net7.n4743 0.007
R32206 net7.n4869 net7.n4868 0.007
R32207 net7.n4899 net7.n4898 0.007
R32208 net7.n4908 net7.n4907 0.007
R32209 net7.n4915 net7.n4914 0.007
R32210 net7.n4999 net7.n4998 0.007
R32211 net7.n5003 net7.n5000 0.007
R32212 net7.n5011 net7.n5006 0.007
R32213 net7.n5018 net7.n5017 0.007
R32214 net7.n5051 net7.n5049 0.007
R32215 net7.n4711 net7.n4710 0.007
R32216 net7.n4705 net7.n4704 0.007
R32217 net7.n4801 net7.n4800 0.007
R32218 net7.n4804 net7.n4803 0.007
R32219 net7.n4845 net7.n4844 0.007
R32220 net7.n4851 net7.n4850 0.007
R32221 net7.n4854 net7.n4853 0.007
R32222 net7.n4936 net7.n4935 0.007
R32223 net7.n4943 net7.n4942 0.007
R32224 net7.n4948 net7.n4947 0.007
R32225 net7.n5137 net7.n5136 0.007
R32226 net7.n5129 net7.n5128 0.007
R32227 net7.n5112 net7.n5111 0.007
R32228 net7.n5106 net7.n5105 0.007
R32229 net7.n5231 net7.n5230 0.007
R32230 net7.n5261 net7.n5260 0.007
R32231 net7.n5270 net7.n5269 0.007
R32232 net7.n5277 net7.n5276 0.007
R32233 net7.n5361 net7.n5360 0.007
R32234 net7.n5365 net7.n5362 0.007
R32235 net7.n5373 net7.n5368 0.007
R32236 net7.n5380 net7.n5379 0.007
R32237 net7.n5413 net7.n5411 0.007
R32238 net7.n5073 net7.n5072 0.007
R32239 net7.n5067 net7.n5066 0.007
R32240 net7.n5163 net7.n5162 0.007
R32241 net7.n5166 net7.n5165 0.007
R32242 net7.n5207 net7.n5206 0.007
R32243 net7.n5213 net7.n5212 0.007
R32244 net7.n5216 net7.n5215 0.007
R32245 net7.n5298 net7.n5297 0.007
R32246 net7.n5305 net7.n5304 0.007
R32247 net7.n5310 net7.n5309 0.007
R32248 net7.n5499 net7.n5498 0.007
R32249 net7.n5491 net7.n5490 0.007
R32250 net7.n5474 net7.n5473 0.007
R32251 net7.n5468 net7.n5467 0.007
R32252 net7.n5593 net7.n5592 0.007
R32253 net7.n5623 net7.n5622 0.007
R32254 net7.n5632 net7.n5631 0.007
R32255 net7.n5639 net7.n5638 0.007
R32256 net7.n5723 net7.n5722 0.007
R32257 net7.n5727 net7.n5724 0.007
R32258 net7.n5735 net7.n5730 0.007
R32259 net7.n5742 net7.n5741 0.007
R32260 net7.n5775 net7.n5773 0.007
R32261 net7.n5435 net7.n5434 0.007
R32262 net7.n5429 net7.n5428 0.007
R32263 net7.n5525 net7.n5524 0.007
R32264 net7.n5528 net7.n5527 0.007
R32265 net7.n5569 net7.n5568 0.007
R32266 net7.n5575 net7.n5574 0.007
R32267 net7.n5578 net7.n5577 0.007
R32268 net7.n5660 net7.n5659 0.007
R32269 net7.n5667 net7.n5666 0.007
R32270 net7.n5672 net7.n5671 0.007
R32271 net7.n5861 net7.n5860 0.007
R32272 net7.n5853 net7.n5852 0.007
R32273 net7.n5836 net7.n5835 0.007
R32274 net7.n5830 net7.n5829 0.007
R32275 net7.n5955 net7.n5954 0.007
R32276 net7.n5985 net7.n5984 0.007
R32277 net7.n5994 net7.n5993 0.007
R32278 net7.n6001 net7.n6000 0.007
R32279 net7.n6085 net7.n6084 0.007
R32280 net7.n6089 net7.n6086 0.007
R32281 net7.n6097 net7.n6092 0.007
R32282 net7.n6104 net7.n6103 0.007
R32283 net7.n6137 net7.n6135 0.007
R32284 net7.n5797 net7.n5796 0.007
R32285 net7.n5791 net7.n5790 0.007
R32286 net7.n5887 net7.n5886 0.007
R32287 net7.n5890 net7.n5889 0.007
R32288 net7.n5931 net7.n5930 0.007
R32289 net7.n5937 net7.n5936 0.007
R32290 net7.n5940 net7.n5939 0.007
R32291 net7.n6022 net7.n6021 0.007
R32292 net7.n6029 net7.n6028 0.007
R32293 net7.n6034 net7.n6033 0.007
R32294 net7.n6223 net7.n6222 0.007
R32295 net7.n6215 net7.n6214 0.007
R32296 net7.n6198 net7.n6197 0.007
R32297 net7.n6192 net7.n6191 0.007
R32298 net7.n6317 net7.n6316 0.007
R32299 net7.n6347 net7.n6346 0.007
R32300 net7.n6356 net7.n6355 0.007
R32301 net7.n6363 net7.n6362 0.007
R32302 net7.n6447 net7.n6446 0.007
R32303 net7.n6451 net7.n6448 0.007
R32304 net7.n6459 net7.n6454 0.007
R32305 net7.n6466 net7.n6465 0.007
R32306 net7.n6499 net7.n6497 0.007
R32307 net7.n6159 net7.n6158 0.007
R32308 net7.n6153 net7.n6152 0.007
R32309 net7.n6249 net7.n6248 0.007
R32310 net7.n6252 net7.n6251 0.007
R32311 net7.n6293 net7.n6292 0.007
R32312 net7.n6299 net7.n6298 0.007
R32313 net7.n6302 net7.n6301 0.007
R32314 net7.n6384 net7.n6383 0.007
R32315 net7.n6391 net7.n6390 0.007
R32316 net7.n6396 net7.n6395 0.007
R32317 net7.n6585 net7.n6584 0.007
R32318 net7.n6577 net7.n6576 0.007
R32319 net7.n6560 net7.n6559 0.007
R32320 net7.n6554 net7.n6553 0.007
R32321 net7.n6679 net7.n6678 0.007
R32322 net7.n6709 net7.n6708 0.007
R32323 net7.n6718 net7.n6717 0.007
R32324 net7.n6725 net7.n6724 0.007
R32325 net7.n6809 net7.n6808 0.007
R32326 net7.n6813 net7.n6810 0.007
R32327 net7.n6821 net7.n6816 0.007
R32328 net7.n6828 net7.n6827 0.007
R32329 net7.n6861 net7.n6859 0.007
R32330 net7.n6521 net7.n6520 0.007
R32331 net7.n6515 net7.n6514 0.007
R32332 net7.n6611 net7.n6610 0.007
R32333 net7.n6614 net7.n6613 0.007
R32334 net7.n6655 net7.n6654 0.007
R32335 net7.n6661 net7.n6660 0.007
R32336 net7.n6664 net7.n6663 0.007
R32337 net7.n6746 net7.n6745 0.007
R32338 net7.n6753 net7.n6752 0.007
R32339 net7.n6758 net7.n6757 0.007
R32340 net7.n6947 net7.n6946 0.007
R32341 net7.n6939 net7.n6938 0.007
R32342 net7.n6922 net7.n6921 0.007
R32343 net7.n6916 net7.n6915 0.007
R32344 net7.n7041 net7.n7040 0.007
R32345 net7.n7071 net7.n7070 0.007
R32346 net7.n7080 net7.n7079 0.007
R32347 net7.n7087 net7.n7086 0.007
R32348 net7.n7171 net7.n7170 0.007
R32349 net7.n7175 net7.n7172 0.007
R32350 net7.n7183 net7.n7178 0.007
R32351 net7.n7190 net7.n7189 0.007
R32352 net7.n7223 net7.n7221 0.007
R32353 net7.n6883 net7.n6882 0.007
R32354 net7.n6877 net7.n6876 0.007
R32355 net7.n6973 net7.n6972 0.007
R32356 net7.n6976 net7.n6975 0.007
R32357 net7.n7017 net7.n7016 0.007
R32358 net7.n7023 net7.n7022 0.007
R32359 net7.n7026 net7.n7025 0.007
R32360 net7.n7108 net7.n7107 0.007
R32361 net7.n7115 net7.n7114 0.007
R32362 net7.n7120 net7.n7119 0.007
R32363 net7.n3593 net7.n3592 0.005
R32364 net7.n3590 net7.n3588 0.005
R32365 net7.n3573 net7.n3572 0.005
R32366 net7.n3564 net7.n3563 0.005
R32367 net7.n3562 net7.n3561 0.005
R32368 net7.n3559 net7.n3558 0.005
R32369 net7.n3558 net7.n3555 0.005
R32370 net7.n3554 net7.n3553 0.005
R32371 net7.n3529 net7.n3528 0.005
R32372 net7.n3373 net7.n3372 0.005
R32373 net7.n3340 net7.n3339 0.005
R32374 net7.n3269 net7.n3268 0.005
R32375 net7.n3296 net7.n3295 0.005
R32376 net7.n3474 net7.n3468 0.005
R32377 net7.n3470 net7.n3469 0.005
R32378 net7.n3464 net7.n3461 0.005
R32379 net7.n3437 net7.n3436 0.005
R32380 net7.n3349 net7.n3348 0.005
R32381 net7.n3258 net7.n3257 0.005
R32382 net7.n3502 net7.n3501 0.005
R32383 net7.n3491 net7.n3490 0.005
R32384 net7.n3460 net7.n3459 0.005
R32385 net7.n3449 net7.n3448 0.005
R32386 net7.n3371 net7.n3370 0.005
R32387 net7.n3360 net7.n3359 0.005
R32388 net7.n3321 net7.n3320 0.005
R32389 net7.n3314 net7.n3313 0.005
R32390 net7.n3231 net7.n3230 0.005
R32391 net7.n3228 net7.n3226 0.005
R32392 net7.n3211 net7.n3210 0.005
R32393 net7.n3202 net7.n3201 0.005
R32394 net7.n3200 net7.n3199 0.005
R32395 net7.n3197 net7.n3196 0.005
R32396 net7.n3196 net7.n3193 0.005
R32397 net7.n3192 net7.n3191 0.005
R32398 net7.n3167 net7.n3166 0.005
R32399 net7.n3011 net7.n3010 0.005
R32400 net7.n2978 net7.n2977 0.005
R32401 net7.n2907 net7.n2906 0.005
R32402 net7.n2934 net7.n2933 0.005
R32403 net7.n3112 net7.n3106 0.005
R32404 net7.n3108 net7.n3107 0.005
R32405 net7.n3102 net7.n3099 0.005
R32406 net7.n3075 net7.n3074 0.005
R32407 net7.n2987 net7.n2986 0.005
R32408 net7.n2896 net7.n2895 0.005
R32409 net7.n3140 net7.n3139 0.005
R32410 net7.n3129 net7.n3128 0.005
R32411 net7.n3098 net7.n3097 0.005
R32412 net7.n3087 net7.n3086 0.005
R32413 net7.n3009 net7.n3008 0.005
R32414 net7.n2998 net7.n2997 0.005
R32415 net7.n2959 net7.n2958 0.005
R32416 net7.n2952 net7.n2951 0.005
R32417 net7.n2869 net7.n2868 0.005
R32418 net7.n2866 net7.n2864 0.005
R32419 net7.n2849 net7.n2848 0.005
R32420 net7.n2840 net7.n2839 0.005
R32421 net7.n2838 net7.n2837 0.005
R32422 net7.n2835 net7.n2834 0.005
R32423 net7.n2834 net7.n2831 0.005
R32424 net7.n2830 net7.n2829 0.005
R32425 net7.n2805 net7.n2804 0.005
R32426 net7.n2649 net7.n2648 0.005
R32427 net7.n2616 net7.n2615 0.005
R32428 net7.n2545 net7.n2544 0.005
R32429 net7.n2572 net7.n2571 0.005
R32430 net7.n2750 net7.n2744 0.005
R32431 net7.n2746 net7.n2745 0.005
R32432 net7.n2740 net7.n2737 0.005
R32433 net7.n2713 net7.n2712 0.005
R32434 net7.n2625 net7.n2624 0.005
R32435 net7.n2534 net7.n2533 0.005
R32436 net7.n2778 net7.n2777 0.005
R32437 net7.n2767 net7.n2766 0.005
R32438 net7.n2736 net7.n2735 0.005
R32439 net7.n2725 net7.n2724 0.005
R32440 net7.n2647 net7.n2646 0.005
R32441 net7.n2636 net7.n2635 0.005
R32442 net7.n2597 net7.n2596 0.005
R32443 net7.n2590 net7.n2589 0.005
R32444 net7.n2507 net7.n2506 0.005
R32445 net7.n2504 net7.n2502 0.005
R32446 net7.n2487 net7.n2486 0.005
R32447 net7.n2478 net7.n2477 0.005
R32448 net7.n2476 net7.n2475 0.005
R32449 net7.n2473 net7.n2472 0.005
R32450 net7.n2472 net7.n2469 0.005
R32451 net7.n2468 net7.n2467 0.005
R32452 net7.n2443 net7.n2442 0.005
R32453 net7.n2287 net7.n2286 0.005
R32454 net7.n2254 net7.n2253 0.005
R32455 net7.n2183 net7.n2182 0.005
R32456 net7.n2210 net7.n2209 0.005
R32457 net7.n2388 net7.n2382 0.005
R32458 net7.n2384 net7.n2383 0.005
R32459 net7.n2378 net7.n2375 0.005
R32460 net7.n2351 net7.n2350 0.005
R32461 net7.n2263 net7.n2262 0.005
R32462 net7.n2172 net7.n2171 0.005
R32463 net7.n2416 net7.n2415 0.005
R32464 net7.n2405 net7.n2404 0.005
R32465 net7.n2374 net7.n2373 0.005
R32466 net7.n2363 net7.n2362 0.005
R32467 net7.n2285 net7.n2284 0.005
R32468 net7.n2274 net7.n2273 0.005
R32469 net7.n2235 net7.n2234 0.005
R32470 net7.n2228 net7.n2227 0.005
R32471 net7.n2145 net7.n2144 0.005
R32472 net7.n2142 net7.n2140 0.005
R32473 net7.n2125 net7.n2124 0.005
R32474 net7.n2116 net7.n2115 0.005
R32475 net7.n2114 net7.n2113 0.005
R32476 net7.n2111 net7.n2110 0.005
R32477 net7.n2110 net7.n2107 0.005
R32478 net7.n2106 net7.n2105 0.005
R32479 net7.n2081 net7.n2080 0.005
R32480 net7.n1925 net7.n1924 0.005
R32481 net7.n1892 net7.n1891 0.005
R32482 net7.n1821 net7.n1820 0.005
R32483 net7.n1848 net7.n1847 0.005
R32484 net7.n2026 net7.n2020 0.005
R32485 net7.n2022 net7.n2021 0.005
R32486 net7.n2016 net7.n2013 0.005
R32487 net7.n1989 net7.n1988 0.005
R32488 net7.n1901 net7.n1900 0.005
R32489 net7.n1810 net7.n1809 0.005
R32490 net7.n2054 net7.n2053 0.005
R32491 net7.n2043 net7.n2042 0.005
R32492 net7.n2012 net7.n2011 0.005
R32493 net7.n2001 net7.n2000 0.005
R32494 net7.n1923 net7.n1922 0.005
R32495 net7.n1912 net7.n1911 0.005
R32496 net7.n1873 net7.n1872 0.005
R32497 net7.n1866 net7.n1865 0.005
R32498 net7.n1783 net7.n1782 0.005
R32499 net7.n1780 net7.n1778 0.005
R32500 net7.n1763 net7.n1762 0.005
R32501 net7.n1754 net7.n1753 0.005
R32502 net7.n1752 net7.n1751 0.005
R32503 net7.n1749 net7.n1748 0.005
R32504 net7.n1748 net7.n1745 0.005
R32505 net7.n1744 net7.n1743 0.005
R32506 net7.n1719 net7.n1718 0.005
R32507 net7.n1563 net7.n1562 0.005
R32508 net7.n1530 net7.n1529 0.005
R32509 net7.n1459 net7.n1458 0.005
R32510 net7.n1486 net7.n1485 0.005
R32511 net7.n1664 net7.n1658 0.005
R32512 net7.n1660 net7.n1659 0.005
R32513 net7.n1654 net7.n1651 0.005
R32514 net7.n1627 net7.n1626 0.005
R32515 net7.n1539 net7.n1538 0.005
R32516 net7.n1448 net7.n1447 0.005
R32517 net7.n1692 net7.n1691 0.005
R32518 net7.n1681 net7.n1680 0.005
R32519 net7.n1650 net7.n1649 0.005
R32520 net7.n1639 net7.n1638 0.005
R32521 net7.n1561 net7.n1560 0.005
R32522 net7.n1550 net7.n1549 0.005
R32523 net7.n1511 net7.n1510 0.005
R32524 net7.n1504 net7.n1503 0.005
R32525 net7.n1421 net7.n1420 0.005
R32526 net7.n1418 net7.n1416 0.005
R32527 net7.n1401 net7.n1400 0.005
R32528 net7.n1392 net7.n1391 0.005
R32529 net7.n1390 net7.n1389 0.005
R32530 net7.n1387 net7.n1386 0.005
R32531 net7.n1386 net7.n1383 0.005
R32532 net7.n1382 net7.n1381 0.005
R32533 net7.n1357 net7.n1356 0.005
R32534 net7.n1201 net7.n1200 0.005
R32535 net7.n1168 net7.n1167 0.005
R32536 net7.n1097 net7.n1096 0.005
R32537 net7.n1124 net7.n1123 0.005
R32538 net7.n1302 net7.n1296 0.005
R32539 net7.n1298 net7.n1297 0.005
R32540 net7.n1292 net7.n1289 0.005
R32541 net7.n1265 net7.n1264 0.005
R32542 net7.n1177 net7.n1176 0.005
R32543 net7.n1086 net7.n1085 0.005
R32544 net7.n1330 net7.n1329 0.005
R32545 net7.n1319 net7.n1318 0.005
R32546 net7.n1288 net7.n1287 0.005
R32547 net7.n1277 net7.n1276 0.005
R32548 net7.n1199 net7.n1198 0.005
R32549 net7.n1188 net7.n1187 0.005
R32550 net7.n1149 net7.n1148 0.005
R32551 net7.n1142 net7.n1141 0.005
R32552 net7.n1059 net7.n1058 0.005
R32553 net7.n1056 net7.n1054 0.005
R32554 net7.n1039 net7.n1038 0.005
R32555 net7.n1030 net7.n1029 0.005
R32556 net7.n1028 net7.n1027 0.005
R32557 net7.n1025 net7.n1024 0.005
R32558 net7.n1024 net7.n1021 0.005
R32559 net7.n1020 net7.n1019 0.005
R32560 net7.n995 net7.n994 0.005
R32561 net7.n839 net7.n838 0.005
R32562 net7.n806 net7.n805 0.005
R32563 net7.n735 net7.n734 0.005
R32564 net7.n762 net7.n761 0.005
R32565 net7.n940 net7.n934 0.005
R32566 net7.n936 net7.n935 0.005
R32567 net7.n930 net7.n927 0.005
R32568 net7.n903 net7.n902 0.005
R32569 net7.n815 net7.n814 0.005
R32570 net7.n724 net7.n723 0.005
R32571 net7.n968 net7.n967 0.005
R32572 net7.n957 net7.n956 0.005
R32573 net7.n926 net7.n925 0.005
R32574 net7.n915 net7.n914 0.005
R32575 net7.n837 net7.n836 0.005
R32576 net7.n826 net7.n825 0.005
R32577 net7.n787 net7.n786 0.005
R32578 net7.n780 net7.n779 0.005
R32579 net7.n697 net7.n696 0.005
R32580 net7.n694 net7.n692 0.005
R32581 net7.n677 net7.n676 0.005
R32582 net7.n668 net7.n667 0.005
R32583 net7.n666 net7.n665 0.005
R32584 net7.n663 net7.n662 0.005
R32585 net7.n662 net7.n659 0.005
R32586 net7.n658 net7.n657 0.005
R32587 net7.n633 net7.n632 0.005
R32588 net7.n477 net7.n476 0.005
R32589 net7.n444 net7.n443 0.005
R32590 net7.n373 net7.n372 0.005
R32591 net7.n400 net7.n399 0.005
R32592 net7.n578 net7.n572 0.005
R32593 net7.n574 net7.n573 0.005
R32594 net7.n568 net7.n565 0.005
R32595 net7.n541 net7.n540 0.005
R32596 net7.n453 net7.n452 0.005
R32597 net7.n362 net7.n361 0.005
R32598 net7.n606 net7.n605 0.005
R32599 net7.n595 net7.n594 0.005
R32600 net7.n564 net7.n563 0.005
R32601 net7.n553 net7.n552 0.005
R32602 net7.n475 net7.n474 0.005
R32603 net7.n464 net7.n463 0.005
R32604 net7.n425 net7.n424 0.005
R32605 net7.n418 net7.n417 0.005
R32606 net7.n336 net7.n335 0.005
R32607 net7.n333 net7.n331 0.005
R32608 net7.n316 net7.n315 0.005
R32609 net7.n307 net7.n306 0.005
R32610 net7.n305 net7.n304 0.005
R32611 net7.n302 net7.n301 0.005
R32612 net7.n301 net7.n298 0.005
R32613 net7.n297 net7.n296 0.005
R32614 net7.n272 net7.n271 0.005
R32615 net7.n116 net7.n115 0.005
R32616 net7.n83 net7.n82 0.005
R32617 net7.n12 net7.n11 0.005
R32618 net7.n39 net7.n38 0.005
R32619 net7.n217 net7.n211 0.005
R32620 net7.n213 net7.n212 0.005
R32621 net7.n207 net7.n204 0.005
R32622 net7.n180 net7.n179 0.005
R32623 net7.n92 net7.n91 0.005
R32624 net7.n1 net7.n0 0.005
R32625 net7.n245 net7.n244 0.005
R32626 net7.n234 net7.n233 0.005
R32627 net7.n203 net7.n202 0.005
R32628 net7.n192 net7.n191 0.005
R32629 net7.n114 net7.n113 0.005
R32630 net7.n103 net7.n102 0.005
R32631 net7.n64 net7.n63 0.005
R32632 net7.n57 net7.n56 0.005
R32633 net7.n3679 net7.n3678 0.005
R32634 net7.n3676 net7.n3674 0.005
R32635 net7.n3662 net7.n3661 0.005
R32636 net7.n3656 net7.n3655 0.005
R32637 net7.n3654 net7.n3653 0.005
R32638 net7.n3651 net7.n3650 0.005
R32639 net7.n3650 net7.n3647 0.005
R32640 net7.n3777 net7.n3776 0.005
R32641 net7.n3806 net7.n3803 0.005
R32642 net7.n3812 net7.n3811 0.005
R32643 net7.n3928 net7.n3927 0.005
R32644 net7.n3936 net7.n3935 0.005
R32645 net7.n3963 net7.n3962 0.005
R32646 net7.n3725 net7.n3722 0.005
R32647 net7.n3731 net7.n3730 0.005
R32648 net7.n3733 net7.n3732 0.005
R32649 net7.n3764 net7.n3763 0.005
R32650 net7.n3868 net7.n3867 0.005
R32651 net7.n3893 net7.n3892 0.005
R32652 net7.n3698 net7.n3697 0.005
R32653 net7.n3705 net7.n3704 0.005
R32654 net7.n3736 net7.n3735 0.005
R32655 net7.n3747 net7.n3746 0.005
R32656 net7.n3843 net7.n3842 0.005
R32657 net7.n3854 net7.n3853 0.005
R32658 net7.n3885 net7.n3884 0.005
R32659 net7.n3896 net7.n3895 0.005
R32660 net7.n4040 net7.n4039 0.005
R32661 net7.n4037 net7.n4035 0.005
R32662 net7.n4023 net7.n4022 0.005
R32663 net7.n4017 net7.n4016 0.005
R32664 net7.n4015 net7.n4014 0.005
R32665 net7.n4012 net7.n4011 0.005
R32666 net7.n4011 net7.n4008 0.005
R32667 net7.n4138 net7.n4137 0.005
R32668 net7.n4167 net7.n4164 0.005
R32669 net7.n4173 net7.n4172 0.005
R32670 net7.n4289 net7.n4288 0.005
R32671 net7.n4297 net7.n4296 0.005
R32672 net7.n4324 net7.n4323 0.005
R32673 net7.n4086 net7.n4083 0.005
R32674 net7.n4092 net7.n4091 0.005
R32675 net7.n4094 net7.n4093 0.005
R32676 net7.n4125 net7.n4124 0.005
R32677 net7.n4229 net7.n4228 0.005
R32678 net7.n4254 net7.n4253 0.005
R32679 net7.n4059 net7.n4058 0.005
R32680 net7.n4066 net7.n4065 0.005
R32681 net7.n4097 net7.n4096 0.005
R32682 net7.n4108 net7.n4107 0.005
R32683 net7.n4204 net7.n4203 0.005
R32684 net7.n4215 net7.n4214 0.005
R32685 net7.n4246 net7.n4245 0.005
R32686 net7.n4257 net7.n4256 0.005
R32687 net7.n4402 net7.n4401 0.005
R32688 net7.n4399 net7.n4397 0.005
R32689 net7.n4385 net7.n4384 0.005
R32690 net7.n4379 net7.n4378 0.005
R32691 net7.n4377 net7.n4376 0.005
R32692 net7.n4374 net7.n4373 0.005
R32693 net7.n4373 net7.n4370 0.005
R32694 net7.n4500 net7.n4499 0.005
R32695 net7.n4529 net7.n4526 0.005
R32696 net7.n4535 net7.n4534 0.005
R32697 net7.n4651 net7.n4650 0.005
R32698 net7.n4659 net7.n4658 0.005
R32699 net7.n4686 net7.n4685 0.005
R32700 net7.n4448 net7.n4445 0.005
R32701 net7.n4454 net7.n4453 0.005
R32702 net7.n4456 net7.n4455 0.005
R32703 net7.n4487 net7.n4486 0.005
R32704 net7.n4591 net7.n4590 0.005
R32705 net7.n4616 net7.n4615 0.005
R32706 net7.n4421 net7.n4420 0.005
R32707 net7.n4428 net7.n4427 0.005
R32708 net7.n4459 net7.n4458 0.005
R32709 net7.n4470 net7.n4469 0.005
R32710 net7.n4566 net7.n4565 0.005
R32711 net7.n4577 net7.n4576 0.005
R32712 net7.n4608 net7.n4607 0.005
R32713 net7.n4619 net7.n4618 0.005
R32714 net7.n4764 net7.n4763 0.005
R32715 net7.n4761 net7.n4759 0.005
R32716 net7.n4747 net7.n4746 0.005
R32717 net7.n4741 net7.n4740 0.005
R32718 net7.n4739 net7.n4738 0.005
R32719 net7.n4736 net7.n4735 0.005
R32720 net7.n4735 net7.n4732 0.005
R32721 net7.n4862 net7.n4861 0.005
R32722 net7.n4891 net7.n4888 0.005
R32723 net7.n4897 net7.n4896 0.005
R32724 net7.n5013 net7.n5012 0.005
R32725 net7.n5021 net7.n5020 0.005
R32726 net7.n5048 net7.n5047 0.005
R32727 net7.n4810 net7.n4807 0.005
R32728 net7.n4816 net7.n4815 0.005
R32729 net7.n4818 net7.n4817 0.005
R32730 net7.n4849 net7.n4848 0.005
R32731 net7.n4953 net7.n4952 0.005
R32732 net7.n4978 net7.n4977 0.005
R32733 net7.n4783 net7.n4782 0.005
R32734 net7.n4790 net7.n4789 0.005
R32735 net7.n4821 net7.n4820 0.005
R32736 net7.n4832 net7.n4831 0.005
R32737 net7.n4928 net7.n4927 0.005
R32738 net7.n4939 net7.n4938 0.005
R32739 net7.n4970 net7.n4969 0.005
R32740 net7.n4981 net7.n4980 0.005
R32741 net7.n5126 net7.n5125 0.005
R32742 net7.n5123 net7.n5121 0.005
R32743 net7.n5109 net7.n5108 0.005
R32744 net7.n5103 net7.n5102 0.005
R32745 net7.n5101 net7.n5100 0.005
R32746 net7.n5098 net7.n5097 0.005
R32747 net7.n5097 net7.n5094 0.005
R32748 net7.n5224 net7.n5223 0.005
R32749 net7.n5253 net7.n5250 0.005
R32750 net7.n5259 net7.n5258 0.005
R32751 net7.n5375 net7.n5374 0.005
R32752 net7.n5383 net7.n5382 0.005
R32753 net7.n5410 net7.n5409 0.005
R32754 net7.n5172 net7.n5169 0.005
R32755 net7.n5178 net7.n5177 0.005
R32756 net7.n5180 net7.n5179 0.005
R32757 net7.n5211 net7.n5210 0.005
R32758 net7.n5315 net7.n5314 0.005
R32759 net7.n5340 net7.n5339 0.005
R32760 net7.n5145 net7.n5144 0.005
R32761 net7.n5152 net7.n5151 0.005
R32762 net7.n5183 net7.n5182 0.005
R32763 net7.n5194 net7.n5193 0.005
R32764 net7.n5290 net7.n5289 0.005
R32765 net7.n5301 net7.n5300 0.005
R32766 net7.n5332 net7.n5331 0.005
R32767 net7.n5343 net7.n5342 0.005
R32768 net7.n5488 net7.n5487 0.005
R32769 net7.n5485 net7.n5483 0.005
R32770 net7.n5471 net7.n5470 0.005
R32771 net7.n5465 net7.n5464 0.005
R32772 net7.n5463 net7.n5462 0.005
R32773 net7.n5460 net7.n5459 0.005
R32774 net7.n5459 net7.n5456 0.005
R32775 net7.n5586 net7.n5585 0.005
R32776 net7.n5615 net7.n5612 0.005
R32777 net7.n5621 net7.n5620 0.005
R32778 net7.n5737 net7.n5736 0.005
R32779 net7.n5745 net7.n5744 0.005
R32780 net7.n5772 net7.n5771 0.005
R32781 net7.n5534 net7.n5531 0.005
R32782 net7.n5540 net7.n5539 0.005
R32783 net7.n5542 net7.n5541 0.005
R32784 net7.n5573 net7.n5572 0.005
R32785 net7.n5677 net7.n5676 0.005
R32786 net7.n5702 net7.n5701 0.005
R32787 net7.n5507 net7.n5506 0.005
R32788 net7.n5514 net7.n5513 0.005
R32789 net7.n5545 net7.n5544 0.005
R32790 net7.n5556 net7.n5555 0.005
R32791 net7.n5652 net7.n5651 0.005
R32792 net7.n5663 net7.n5662 0.005
R32793 net7.n5694 net7.n5693 0.005
R32794 net7.n5705 net7.n5704 0.005
R32795 net7.n5850 net7.n5849 0.005
R32796 net7.n5847 net7.n5845 0.005
R32797 net7.n5833 net7.n5832 0.005
R32798 net7.n5827 net7.n5826 0.005
R32799 net7.n5825 net7.n5824 0.005
R32800 net7.n5822 net7.n5821 0.005
R32801 net7.n5821 net7.n5818 0.005
R32802 net7.n5948 net7.n5947 0.005
R32803 net7.n5977 net7.n5974 0.005
R32804 net7.n5983 net7.n5982 0.005
R32805 net7.n6099 net7.n6098 0.005
R32806 net7.n6107 net7.n6106 0.005
R32807 net7.n6134 net7.n6133 0.005
R32808 net7.n5896 net7.n5893 0.005
R32809 net7.n5902 net7.n5901 0.005
R32810 net7.n5904 net7.n5903 0.005
R32811 net7.n5935 net7.n5934 0.005
R32812 net7.n6039 net7.n6038 0.005
R32813 net7.n6064 net7.n6063 0.005
R32814 net7.n5869 net7.n5868 0.005
R32815 net7.n5876 net7.n5875 0.005
R32816 net7.n5907 net7.n5906 0.005
R32817 net7.n5918 net7.n5917 0.005
R32818 net7.n6014 net7.n6013 0.005
R32819 net7.n6025 net7.n6024 0.005
R32820 net7.n6056 net7.n6055 0.005
R32821 net7.n6067 net7.n6066 0.005
R32822 net7.n6212 net7.n6211 0.005
R32823 net7.n6209 net7.n6207 0.005
R32824 net7.n6195 net7.n6194 0.005
R32825 net7.n6189 net7.n6188 0.005
R32826 net7.n6187 net7.n6186 0.005
R32827 net7.n6184 net7.n6183 0.005
R32828 net7.n6183 net7.n6180 0.005
R32829 net7.n6310 net7.n6309 0.005
R32830 net7.n6339 net7.n6336 0.005
R32831 net7.n6345 net7.n6344 0.005
R32832 net7.n6461 net7.n6460 0.005
R32833 net7.n6469 net7.n6468 0.005
R32834 net7.n6496 net7.n6495 0.005
R32835 net7.n6258 net7.n6255 0.005
R32836 net7.n6264 net7.n6263 0.005
R32837 net7.n6266 net7.n6265 0.005
R32838 net7.n6297 net7.n6296 0.005
R32839 net7.n6401 net7.n6400 0.005
R32840 net7.n6426 net7.n6425 0.005
R32841 net7.n6231 net7.n6230 0.005
R32842 net7.n6238 net7.n6237 0.005
R32843 net7.n6269 net7.n6268 0.005
R32844 net7.n6280 net7.n6279 0.005
R32845 net7.n6376 net7.n6375 0.005
R32846 net7.n6387 net7.n6386 0.005
R32847 net7.n6418 net7.n6417 0.005
R32848 net7.n6429 net7.n6428 0.005
R32849 net7.n6574 net7.n6573 0.005
R32850 net7.n6571 net7.n6569 0.005
R32851 net7.n6557 net7.n6556 0.005
R32852 net7.n6551 net7.n6550 0.005
R32853 net7.n6549 net7.n6548 0.005
R32854 net7.n6546 net7.n6545 0.005
R32855 net7.n6545 net7.n6542 0.005
R32856 net7.n6672 net7.n6671 0.005
R32857 net7.n6701 net7.n6698 0.005
R32858 net7.n6707 net7.n6706 0.005
R32859 net7.n6823 net7.n6822 0.005
R32860 net7.n6831 net7.n6830 0.005
R32861 net7.n6858 net7.n6857 0.005
R32862 net7.n6620 net7.n6617 0.005
R32863 net7.n6626 net7.n6625 0.005
R32864 net7.n6628 net7.n6627 0.005
R32865 net7.n6659 net7.n6658 0.005
R32866 net7.n6763 net7.n6762 0.005
R32867 net7.n6788 net7.n6787 0.005
R32868 net7.n6593 net7.n6592 0.005
R32869 net7.n6600 net7.n6599 0.005
R32870 net7.n6631 net7.n6630 0.005
R32871 net7.n6642 net7.n6641 0.005
R32872 net7.n6738 net7.n6737 0.005
R32873 net7.n6749 net7.n6748 0.005
R32874 net7.n6780 net7.n6779 0.005
R32875 net7.n6791 net7.n6790 0.005
R32876 net7.n6936 net7.n6935 0.005
R32877 net7.n6933 net7.n6931 0.005
R32878 net7.n6919 net7.n6918 0.005
R32879 net7.n6913 net7.n6912 0.005
R32880 net7.n6911 net7.n6910 0.005
R32881 net7.n6908 net7.n6907 0.005
R32882 net7.n6907 net7.n6904 0.005
R32883 net7.n7034 net7.n7033 0.005
R32884 net7.n7063 net7.n7060 0.005
R32885 net7.n7069 net7.n7068 0.005
R32886 net7.n7185 net7.n7184 0.005
R32887 net7.n7193 net7.n7192 0.005
R32888 net7.n7220 net7.n7219 0.005
R32889 net7.n6982 net7.n6979 0.005
R32890 net7.n6988 net7.n6987 0.005
R32891 net7.n6990 net7.n6989 0.005
R32892 net7.n7021 net7.n7020 0.005
R32893 net7.n7125 net7.n7124 0.005
R32894 net7.n7150 net7.n7149 0.005
R32895 net7.n6955 net7.n6954 0.005
R32896 net7.n6962 net7.n6961 0.005
R32897 net7.n6993 net7.n6992 0.005
R32898 net7.n7004 net7.n7003 0.005
R32899 net7.n7100 net7.n7099 0.005
R32900 net7.n7111 net7.n7110 0.005
R32901 net7.n7142 net7.n7141 0.005
R32902 net7.n7153 net7.n7152 0.005
R32903 net7.n3604 net7.n3603 0.003
R32904 net7.n3417 net7.n3386 0.003
R32905 net7.n3414 net7.n3412 0.003
R32906 net7.n3398 net7.n3397 0.003
R32907 net7.n3273 net7.n3269 0.003
R32908 net7.n3287 net7.n3285 0.003
R32909 net7.n3293 net7.n3292 0.003
R32910 net7.n3304 net7.n3303 0.003
R32911 net7.n3617 net7.n3509 0.003
R32912 net7.n3484 net7.n3483 0.003
R32913 net7.n3475 net7.n3467 0.003
R32914 net7.n3440 net7.n3439 0.003
R32915 net7.n3430 net7.n3423 0.003
R32916 net7.n3351 net7.n3350 0.003
R32917 net7.n3335 net7.n3328 0.003
R32918 net7.n3242 net7.n3241 0.003
R32919 net7.n3055 net7.n3024 0.003
R32920 net7.n3052 net7.n3050 0.003
R32921 net7.n3036 net7.n3035 0.003
R32922 net7.n2911 net7.n2907 0.003
R32923 net7.n2925 net7.n2923 0.003
R32924 net7.n2931 net7.n2930 0.003
R32925 net7.n2942 net7.n2941 0.003
R32926 net7.n3255 net7.n3147 0.003
R32927 net7.n3122 net7.n3121 0.003
R32928 net7.n3113 net7.n3105 0.003
R32929 net7.n3078 net7.n3077 0.003
R32930 net7.n3068 net7.n3061 0.003
R32931 net7.n2989 net7.n2988 0.003
R32932 net7.n2973 net7.n2966 0.003
R32933 net7.n2880 net7.n2879 0.003
R32934 net7.n2693 net7.n2662 0.003
R32935 net7.n2690 net7.n2688 0.003
R32936 net7.n2674 net7.n2673 0.003
R32937 net7.n2549 net7.n2545 0.003
R32938 net7.n2563 net7.n2561 0.003
R32939 net7.n2569 net7.n2568 0.003
R32940 net7.n2580 net7.n2579 0.003
R32941 net7.n2893 net7.n2785 0.003
R32942 net7.n2760 net7.n2759 0.003
R32943 net7.n2751 net7.n2743 0.003
R32944 net7.n2716 net7.n2715 0.003
R32945 net7.n2706 net7.n2699 0.003
R32946 net7.n2627 net7.n2626 0.003
R32947 net7.n2611 net7.n2604 0.003
R32948 net7.n2518 net7.n2517 0.003
R32949 net7.n2331 net7.n2300 0.003
R32950 net7.n2328 net7.n2326 0.003
R32951 net7.n2312 net7.n2311 0.003
R32952 net7.n2187 net7.n2183 0.003
R32953 net7.n2201 net7.n2199 0.003
R32954 net7.n2207 net7.n2206 0.003
R32955 net7.n2218 net7.n2217 0.003
R32956 net7.n2531 net7.n2423 0.003
R32957 net7.n2398 net7.n2397 0.003
R32958 net7.n2389 net7.n2381 0.003
R32959 net7.n2354 net7.n2353 0.003
R32960 net7.n2344 net7.n2337 0.003
R32961 net7.n2265 net7.n2264 0.003
R32962 net7.n2249 net7.n2242 0.003
R32963 net7.n2156 net7.n2155 0.003
R32964 net7.n1969 net7.n1938 0.003
R32965 net7.n1966 net7.n1964 0.003
R32966 net7.n1950 net7.n1949 0.003
R32967 net7.n1825 net7.n1821 0.003
R32968 net7.n1839 net7.n1837 0.003
R32969 net7.n1845 net7.n1844 0.003
R32970 net7.n1856 net7.n1855 0.003
R32971 net7.n2169 net7.n2061 0.003
R32972 net7.n2036 net7.n2035 0.003
R32973 net7.n2027 net7.n2019 0.003
R32974 net7.n1992 net7.n1991 0.003
R32975 net7.n1982 net7.n1975 0.003
R32976 net7.n1903 net7.n1902 0.003
R32977 net7.n1887 net7.n1880 0.003
R32978 net7.n1794 net7.n1793 0.003
R32979 net7.n1607 net7.n1576 0.003
R32980 net7.n1604 net7.n1602 0.003
R32981 net7.n1588 net7.n1587 0.003
R32982 net7.n1463 net7.n1459 0.003
R32983 net7.n1477 net7.n1475 0.003
R32984 net7.n1483 net7.n1482 0.003
R32985 net7.n1494 net7.n1493 0.003
R32986 net7.n1807 net7.n1699 0.003
R32987 net7.n1674 net7.n1673 0.003
R32988 net7.n1665 net7.n1657 0.003
R32989 net7.n1630 net7.n1629 0.003
R32990 net7.n1620 net7.n1613 0.003
R32991 net7.n1541 net7.n1540 0.003
R32992 net7.n1525 net7.n1518 0.003
R32993 net7.n1432 net7.n1431 0.003
R32994 net7.n1245 net7.n1214 0.003
R32995 net7.n1242 net7.n1240 0.003
R32996 net7.n1226 net7.n1225 0.003
R32997 net7.n1101 net7.n1097 0.003
R32998 net7.n1115 net7.n1113 0.003
R32999 net7.n1121 net7.n1120 0.003
R33000 net7.n1132 net7.n1131 0.003
R33001 net7.n1445 net7.n1337 0.003
R33002 net7.n1312 net7.n1311 0.003
R33003 net7.n1303 net7.n1295 0.003
R33004 net7.n1268 net7.n1267 0.003
R33005 net7.n1258 net7.n1251 0.003
R33006 net7.n1179 net7.n1178 0.003
R33007 net7.n1163 net7.n1156 0.003
R33008 net7.n1070 net7.n1069 0.003
R33009 net7.n883 net7.n852 0.003
R33010 net7.n880 net7.n878 0.003
R33011 net7.n864 net7.n863 0.003
R33012 net7.n739 net7.n735 0.003
R33013 net7.n753 net7.n751 0.003
R33014 net7.n759 net7.n758 0.003
R33015 net7.n770 net7.n769 0.003
R33016 net7.n1083 net7.n975 0.003
R33017 net7.n950 net7.n949 0.003
R33018 net7.n941 net7.n933 0.003
R33019 net7.n906 net7.n905 0.003
R33020 net7.n896 net7.n889 0.003
R33021 net7.n817 net7.n816 0.003
R33022 net7.n801 net7.n794 0.003
R33023 net7.n708 net7.n707 0.003
R33024 net7.n521 net7.n490 0.003
R33025 net7.n518 net7.n516 0.003
R33026 net7.n502 net7.n501 0.003
R33027 net7.n377 net7.n373 0.003
R33028 net7.n391 net7.n389 0.003
R33029 net7.n397 net7.n396 0.003
R33030 net7.n408 net7.n407 0.003
R33031 net7.n721 net7.n613 0.003
R33032 net7.n588 net7.n587 0.003
R33033 net7.n579 net7.n571 0.003
R33034 net7.n544 net7.n543 0.003
R33035 net7.n534 net7.n527 0.003
R33036 net7.n455 net7.n454 0.003
R33037 net7.n439 net7.n432 0.003
R33038 net7.n347 net7.n346 0.003
R33039 net7.n160 net7.n129 0.003
R33040 net7.n157 net7.n155 0.003
R33041 net7.n141 net7.n140 0.003
R33042 net7.n16 net7.n12 0.003
R33043 net7.n30 net7.n28 0.003
R33044 net7.n36 net7.n35 0.003
R33045 net7.n47 net7.n46 0.003
R33046 net7.n360 net7.n252 0.003
R33047 net7.n227 net7.n226 0.003
R33048 net7.n218 net7.n210 0.003
R33049 net7.n183 net7.n182 0.003
R33050 net7.n173 net7.n166 0.003
R33051 net7.n94 net7.n93 0.003
R33052 net7.n78 net7.n71 0.003
R33053 net7.n3688 net7.n3687 0.003
R33054 net7.n3839 net7.n3825 0.003
R33055 net7.n3838 net7.n3836 0.003
R33056 net7.n3919 net7.n3918 0.003
R33057 net7.n3940 net7.n3936 0.003
R33058 net7.n3954 net7.n3952 0.003
R33059 net7.n3960 net7.n3959 0.003
R33060 net7.n3971 net7.n3970 0.003
R33061 net7.n3717 net7.n3711 0.003
R33062 net7.n3727 net7.n3726 0.003
R33063 net7.n3762 net7.n3754 0.003
R33064 net7.n3772 net7.n3771 0.003
R33065 net7.n3869 net7.n3861 0.003
R33066 net7.n3876 net7.n3875 0.003
R33067 net7.n3979 net7.n3904 0.003
R33068 net7.n4049 net7.n4048 0.003
R33069 net7.n4200 net7.n4186 0.003
R33070 net7.n4199 net7.n4197 0.003
R33071 net7.n4280 net7.n4279 0.003
R33072 net7.n4301 net7.n4297 0.003
R33073 net7.n4315 net7.n4313 0.003
R33074 net7.n4321 net7.n4320 0.003
R33075 net7.n4332 net7.n4331 0.003
R33076 net7.n4078 net7.n4072 0.003
R33077 net7.n4088 net7.n4087 0.003
R33078 net7.n4123 net7.n4115 0.003
R33079 net7.n4133 net7.n4132 0.003
R33080 net7.n4230 net7.n4222 0.003
R33081 net7.n4237 net7.n4236 0.003
R33082 net7.n4340 net7.n4265 0.003
R33083 net7.n4411 net7.n4410 0.003
R33084 net7.n4562 net7.n4548 0.003
R33085 net7.n4561 net7.n4559 0.003
R33086 net7.n4642 net7.n4641 0.003
R33087 net7.n4663 net7.n4659 0.003
R33088 net7.n4677 net7.n4675 0.003
R33089 net7.n4683 net7.n4682 0.003
R33090 net7.n4694 net7.n4693 0.003
R33091 net7.n4440 net7.n4434 0.003
R33092 net7.n4450 net7.n4449 0.003
R33093 net7.n4485 net7.n4477 0.003
R33094 net7.n4495 net7.n4494 0.003
R33095 net7.n4592 net7.n4584 0.003
R33096 net7.n4599 net7.n4598 0.003
R33097 net7.n4702 net7.n4627 0.003
R33098 net7.n4773 net7.n4772 0.003
R33099 net7.n4924 net7.n4910 0.003
R33100 net7.n4923 net7.n4921 0.003
R33101 net7.n5004 net7.n5003 0.003
R33102 net7.n5025 net7.n5021 0.003
R33103 net7.n5039 net7.n5037 0.003
R33104 net7.n5045 net7.n5044 0.003
R33105 net7.n5056 net7.n5055 0.003
R33106 net7.n4802 net7.n4796 0.003
R33107 net7.n4812 net7.n4811 0.003
R33108 net7.n4847 net7.n4839 0.003
R33109 net7.n4857 net7.n4856 0.003
R33110 net7.n4954 net7.n4946 0.003
R33111 net7.n4961 net7.n4960 0.003
R33112 net7.n5064 net7.n4989 0.003
R33113 net7.n5135 net7.n5134 0.003
R33114 net7.n5286 net7.n5272 0.003
R33115 net7.n5285 net7.n5283 0.003
R33116 net7.n5366 net7.n5365 0.003
R33117 net7.n5387 net7.n5383 0.003
R33118 net7.n5401 net7.n5399 0.003
R33119 net7.n5407 net7.n5406 0.003
R33120 net7.n5418 net7.n5417 0.003
R33121 net7.n5164 net7.n5158 0.003
R33122 net7.n5174 net7.n5173 0.003
R33123 net7.n5209 net7.n5201 0.003
R33124 net7.n5219 net7.n5218 0.003
R33125 net7.n5316 net7.n5308 0.003
R33126 net7.n5323 net7.n5322 0.003
R33127 net7.n5426 net7.n5351 0.003
R33128 net7.n5497 net7.n5496 0.003
R33129 net7.n5648 net7.n5634 0.003
R33130 net7.n5647 net7.n5645 0.003
R33131 net7.n5728 net7.n5727 0.003
R33132 net7.n5749 net7.n5745 0.003
R33133 net7.n5763 net7.n5761 0.003
R33134 net7.n5769 net7.n5768 0.003
R33135 net7.n5780 net7.n5779 0.003
R33136 net7.n5526 net7.n5520 0.003
R33137 net7.n5536 net7.n5535 0.003
R33138 net7.n5571 net7.n5563 0.003
R33139 net7.n5581 net7.n5580 0.003
R33140 net7.n5678 net7.n5670 0.003
R33141 net7.n5685 net7.n5684 0.003
R33142 net7.n5788 net7.n5713 0.003
R33143 net7.n5859 net7.n5858 0.003
R33144 net7.n6010 net7.n5996 0.003
R33145 net7.n6009 net7.n6007 0.003
R33146 net7.n6090 net7.n6089 0.003
R33147 net7.n6111 net7.n6107 0.003
R33148 net7.n6125 net7.n6123 0.003
R33149 net7.n6131 net7.n6130 0.003
R33150 net7.n6142 net7.n6141 0.003
R33151 net7.n5888 net7.n5882 0.003
R33152 net7.n5898 net7.n5897 0.003
R33153 net7.n5933 net7.n5925 0.003
R33154 net7.n5943 net7.n5942 0.003
R33155 net7.n6040 net7.n6032 0.003
R33156 net7.n6047 net7.n6046 0.003
R33157 net7.n6150 net7.n6075 0.003
R33158 net7.n6221 net7.n6220 0.003
R33159 net7.n6372 net7.n6358 0.003
R33160 net7.n6371 net7.n6369 0.003
R33161 net7.n6452 net7.n6451 0.003
R33162 net7.n6473 net7.n6469 0.003
R33163 net7.n6487 net7.n6485 0.003
R33164 net7.n6493 net7.n6492 0.003
R33165 net7.n6504 net7.n6503 0.003
R33166 net7.n6250 net7.n6244 0.003
R33167 net7.n6260 net7.n6259 0.003
R33168 net7.n6295 net7.n6287 0.003
R33169 net7.n6305 net7.n6304 0.003
R33170 net7.n6402 net7.n6394 0.003
R33171 net7.n6409 net7.n6408 0.003
R33172 net7.n6512 net7.n6437 0.003
R33173 net7.n6583 net7.n6582 0.003
R33174 net7.n6734 net7.n6720 0.003
R33175 net7.n6733 net7.n6731 0.003
R33176 net7.n6814 net7.n6813 0.003
R33177 net7.n6835 net7.n6831 0.003
R33178 net7.n6849 net7.n6847 0.003
R33179 net7.n6855 net7.n6854 0.003
R33180 net7.n6866 net7.n6865 0.003
R33181 net7.n6612 net7.n6606 0.003
R33182 net7.n6622 net7.n6621 0.003
R33183 net7.n6657 net7.n6649 0.003
R33184 net7.n6667 net7.n6666 0.003
R33185 net7.n6764 net7.n6756 0.003
R33186 net7.n6771 net7.n6770 0.003
R33187 net7.n6874 net7.n6799 0.003
R33188 net7.n6945 net7.n6944 0.003
R33189 net7.n7096 net7.n7082 0.003
R33190 net7.n7095 net7.n7093 0.003
R33191 net7.n7176 net7.n7175 0.003
R33192 net7.n7197 net7.n7193 0.003
R33193 net7.n7211 net7.n7209 0.003
R33194 net7.n7217 net7.n7216 0.003
R33195 net7.n7228 net7.n7227 0.003
R33196 net7.n6974 net7.n6968 0.003
R33197 net7.n6984 net7.n6983 0.003
R33198 net7.n7019 net7.n7011 0.003
R33199 net7.n7029 net7.n7028 0.003
R33200 net7.n7126 net7.n7118 0.003
R33201 net7.n7133 net7.n7132 0.003
R33202 net7.n7236 net7.n7161 0.003
R33203 net7.n3585 net7.n3584 0.001
R33204 net7.n3580 net7.n3578 0.001
R33205 net7.n3574 net7.n3573 0.001
R33206 net7.n3569 net7.n3568 0.001
R33207 net7.n3552 net7.n3549 0.001
R33208 net7.n3546 net7.n3545 0.001
R33209 net7.n3541 net7.n3538 0.001
R33210 net7.n3536 net7.n3535 0.001
R33211 net7.n3535 net7.n3532 0.001
R33212 net7.n3531 net7.n3530 0.001
R33213 net7.n3525 net7.n3524 0.001
R33214 net7.n3380 net7.n3376 0.001
R33215 net7.n3281 net7.n3278 0.001
R33216 net7.n3283 net7.n3282 0.001
R33217 net7.n3477 net7.n3476 0.001
R33218 net7.n3479 net7.n3478 0.001
R33219 net7.n3446 net7.n3445 0.001
R33220 net7.n3444 net7.n3443 0.001
R33221 net7.n3438 net7.n3433 0.001
R33222 net7.n3429 net7.n3428 0.001
R33223 net7.n3331 net7.n3330 0.001
R33224 net7.n3325 net7.n3324 0.001
R33225 net7.n3261 net7.n3260 0.001
R33226 net7.n3223 net7.n3222 0.001
R33227 net7.n3218 net7.n3216 0.001
R33228 net7.n3212 net7.n3211 0.001
R33229 net7.n3207 net7.n3206 0.001
R33230 net7.n3190 net7.n3187 0.001
R33231 net7.n3184 net7.n3183 0.001
R33232 net7.n3179 net7.n3176 0.001
R33233 net7.n3174 net7.n3173 0.001
R33234 net7.n3173 net7.n3170 0.001
R33235 net7.n3169 net7.n3168 0.001
R33236 net7.n3163 net7.n3162 0.001
R33237 net7.n3018 net7.n3014 0.001
R33238 net7.n2919 net7.n2916 0.001
R33239 net7.n2921 net7.n2920 0.001
R33240 net7.n3115 net7.n3114 0.001
R33241 net7.n3117 net7.n3116 0.001
R33242 net7.n3084 net7.n3083 0.001
R33243 net7.n3082 net7.n3081 0.001
R33244 net7.n3076 net7.n3071 0.001
R33245 net7.n3067 net7.n3066 0.001
R33246 net7.n2969 net7.n2968 0.001
R33247 net7.n2963 net7.n2962 0.001
R33248 net7.n2899 net7.n2898 0.001
R33249 net7.n2861 net7.n2860 0.001
R33250 net7.n2856 net7.n2854 0.001
R33251 net7.n2850 net7.n2849 0.001
R33252 net7.n2845 net7.n2844 0.001
R33253 net7.n2828 net7.n2825 0.001
R33254 net7.n2822 net7.n2821 0.001
R33255 net7.n2817 net7.n2814 0.001
R33256 net7.n2812 net7.n2811 0.001
R33257 net7.n2811 net7.n2808 0.001
R33258 net7.n2807 net7.n2806 0.001
R33259 net7.n2801 net7.n2800 0.001
R33260 net7.n2656 net7.n2652 0.001
R33261 net7.n2557 net7.n2554 0.001
R33262 net7.n2559 net7.n2558 0.001
R33263 net7.n2753 net7.n2752 0.001
R33264 net7.n2755 net7.n2754 0.001
R33265 net7.n2722 net7.n2721 0.001
R33266 net7.n2720 net7.n2719 0.001
R33267 net7.n2714 net7.n2709 0.001
R33268 net7.n2705 net7.n2704 0.001
R33269 net7.n2607 net7.n2606 0.001
R33270 net7.n2601 net7.n2600 0.001
R33271 net7.n2537 net7.n2536 0.001
R33272 net7.n2499 net7.n2498 0.001
R33273 net7.n2494 net7.n2492 0.001
R33274 net7.n2488 net7.n2487 0.001
R33275 net7.n2483 net7.n2482 0.001
R33276 net7.n2466 net7.n2463 0.001
R33277 net7.n2460 net7.n2459 0.001
R33278 net7.n2455 net7.n2452 0.001
R33279 net7.n2450 net7.n2449 0.001
R33280 net7.n2449 net7.n2446 0.001
R33281 net7.n2445 net7.n2444 0.001
R33282 net7.n2439 net7.n2438 0.001
R33283 net7.n2294 net7.n2290 0.001
R33284 net7.n2195 net7.n2192 0.001
R33285 net7.n2197 net7.n2196 0.001
R33286 net7.n2391 net7.n2390 0.001
R33287 net7.n2393 net7.n2392 0.001
R33288 net7.n2360 net7.n2359 0.001
R33289 net7.n2358 net7.n2357 0.001
R33290 net7.n2352 net7.n2347 0.001
R33291 net7.n2343 net7.n2342 0.001
R33292 net7.n2245 net7.n2244 0.001
R33293 net7.n2239 net7.n2238 0.001
R33294 net7.n2175 net7.n2174 0.001
R33295 net7.n2137 net7.n2136 0.001
R33296 net7.n2132 net7.n2130 0.001
R33297 net7.n2126 net7.n2125 0.001
R33298 net7.n2121 net7.n2120 0.001
R33299 net7.n2104 net7.n2101 0.001
R33300 net7.n2098 net7.n2097 0.001
R33301 net7.n2093 net7.n2090 0.001
R33302 net7.n2088 net7.n2087 0.001
R33303 net7.n2087 net7.n2084 0.001
R33304 net7.n2083 net7.n2082 0.001
R33305 net7.n2077 net7.n2076 0.001
R33306 net7.n1932 net7.n1928 0.001
R33307 net7.n1833 net7.n1830 0.001
R33308 net7.n1835 net7.n1834 0.001
R33309 net7.n2029 net7.n2028 0.001
R33310 net7.n2031 net7.n2030 0.001
R33311 net7.n1998 net7.n1997 0.001
R33312 net7.n1996 net7.n1995 0.001
R33313 net7.n1990 net7.n1985 0.001
R33314 net7.n1981 net7.n1980 0.001
R33315 net7.n1883 net7.n1882 0.001
R33316 net7.n1877 net7.n1876 0.001
R33317 net7.n1813 net7.n1812 0.001
R33318 net7.n1775 net7.n1774 0.001
R33319 net7.n1770 net7.n1768 0.001
R33320 net7.n1764 net7.n1763 0.001
R33321 net7.n1759 net7.n1758 0.001
R33322 net7.n1742 net7.n1739 0.001
R33323 net7.n1736 net7.n1735 0.001
R33324 net7.n1731 net7.n1728 0.001
R33325 net7.n1726 net7.n1725 0.001
R33326 net7.n1725 net7.n1722 0.001
R33327 net7.n1721 net7.n1720 0.001
R33328 net7.n1715 net7.n1714 0.001
R33329 net7.n1570 net7.n1566 0.001
R33330 net7.n1471 net7.n1468 0.001
R33331 net7.n1473 net7.n1472 0.001
R33332 net7.n1667 net7.n1666 0.001
R33333 net7.n1669 net7.n1668 0.001
R33334 net7.n1636 net7.n1635 0.001
R33335 net7.n1634 net7.n1633 0.001
R33336 net7.n1628 net7.n1623 0.001
R33337 net7.n1619 net7.n1618 0.001
R33338 net7.n1521 net7.n1520 0.001
R33339 net7.n1515 net7.n1514 0.001
R33340 net7.n1451 net7.n1450 0.001
R33341 net7.n1413 net7.n1412 0.001
R33342 net7.n1408 net7.n1406 0.001
R33343 net7.n1402 net7.n1401 0.001
R33344 net7.n1397 net7.n1396 0.001
R33345 net7.n1380 net7.n1377 0.001
R33346 net7.n1374 net7.n1373 0.001
R33347 net7.n1369 net7.n1366 0.001
R33348 net7.n1364 net7.n1363 0.001
R33349 net7.n1363 net7.n1360 0.001
R33350 net7.n1359 net7.n1358 0.001
R33351 net7.n1353 net7.n1352 0.001
R33352 net7.n1208 net7.n1204 0.001
R33353 net7.n1109 net7.n1106 0.001
R33354 net7.n1111 net7.n1110 0.001
R33355 net7.n1305 net7.n1304 0.001
R33356 net7.n1307 net7.n1306 0.001
R33357 net7.n1274 net7.n1273 0.001
R33358 net7.n1272 net7.n1271 0.001
R33359 net7.n1266 net7.n1261 0.001
R33360 net7.n1257 net7.n1256 0.001
R33361 net7.n1159 net7.n1158 0.001
R33362 net7.n1153 net7.n1152 0.001
R33363 net7.n1089 net7.n1088 0.001
R33364 net7.n1051 net7.n1050 0.001
R33365 net7.n1046 net7.n1044 0.001
R33366 net7.n1040 net7.n1039 0.001
R33367 net7.n1035 net7.n1034 0.001
R33368 net7.n1018 net7.n1015 0.001
R33369 net7.n1012 net7.n1011 0.001
R33370 net7.n1007 net7.n1004 0.001
R33371 net7.n1002 net7.n1001 0.001
R33372 net7.n1001 net7.n998 0.001
R33373 net7.n997 net7.n996 0.001
R33374 net7.n991 net7.n990 0.001
R33375 net7.n846 net7.n842 0.001
R33376 net7.n747 net7.n744 0.001
R33377 net7.n749 net7.n748 0.001
R33378 net7.n943 net7.n942 0.001
R33379 net7.n945 net7.n944 0.001
R33380 net7.n912 net7.n911 0.001
R33381 net7.n910 net7.n909 0.001
R33382 net7.n904 net7.n899 0.001
R33383 net7.n895 net7.n894 0.001
R33384 net7.n797 net7.n796 0.001
R33385 net7.n791 net7.n790 0.001
R33386 net7.n727 net7.n726 0.001
R33387 net7.n689 net7.n688 0.001
R33388 net7.n684 net7.n682 0.001
R33389 net7.n678 net7.n677 0.001
R33390 net7.n673 net7.n672 0.001
R33391 net7.n656 net7.n653 0.001
R33392 net7.n650 net7.n649 0.001
R33393 net7.n645 net7.n642 0.001
R33394 net7.n640 net7.n639 0.001
R33395 net7.n639 net7.n636 0.001
R33396 net7.n635 net7.n634 0.001
R33397 net7.n629 net7.n628 0.001
R33398 net7.n484 net7.n480 0.001
R33399 net7.n385 net7.n382 0.001
R33400 net7.n387 net7.n386 0.001
R33401 net7.n581 net7.n580 0.001
R33402 net7.n583 net7.n582 0.001
R33403 net7.n550 net7.n549 0.001
R33404 net7.n548 net7.n547 0.001
R33405 net7.n542 net7.n537 0.001
R33406 net7.n533 net7.n532 0.001
R33407 net7.n435 net7.n434 0.001
R33408 net7.n429 net7.n428 0.001
R33409 net7.n365 net7.n364 0.001
R33410 net7.n328 net7.n327 0.001
R33411 net7.n323 net7.n321 0.001
R33412 net7.n317 net7.n316 0.001
R33413 net7.n312 net7.n311 0.001
R33414 net7.n295 net7.n292 0.001
R33415 net7.n289 net7.n288 0.001
R33416 net7.n284 net7.n281 0.001
R33417 net7.n279 net7.n278 0.001
R33418 net7.n278 net7.n275 0.001
R33419 net7.n274 net7.n273 0.001
R33420 net7.n268 net7.n267 0.001
R33421 net7.n123 net7.n119 0.001
R33422 net7.n24 net7.n21 0.001
R33423 net7.n26 net7.n25 0.001
R33424 net7.n220 net7.n219 0.001
R33425 net7.n222 net7.n221 0.001
R33426 net7.n189 net7.n188 0.001
R33427 net7.n187 net7.n186 0.001
R33428 net7.n181 net7.n176 0.001
R33429 net7.n172 net7.n171 0.001
R33430 net7.n74 net7.n73 0.001
R33431 net7.n68 net7.n67 0.001
R33432 net7.n4 net7.n3 0.001
R33433 net7.n3671 net7.n3670 0.001
R33434 net7.n3669 net7.n3667 0.001
R33435 net7.n3663 net7.n3662 0.001
R33436 net7.n3658 net7.n3657 0.001
R33437 net7.n3782 net7.n3780 0.001
R33438 net7.n3787 net7.n3784 0.001
R33439 net7.n3795 net7.n3793 0.001
R33440 net7.n3799 net7.n3796 0.001
R33441 net7.n3800 net7.n3799 0.001
R33442 net7.n3802 net7.n3801 0.001
R33443 net7.n3810 net7.n3809 0.001
R33444 net7.n3819 net7.n3815 0.001
R33445 net7.n3948 net7.n3945 0.001
R33446 net7.n3950 net7.n3949 0.001
R33447 net7.n3715 net7.n3714 0.001
R33448 net7.n3721 net7.n3720 0.001
R33449 net7.n3751 net7.n3750 0.001
R33450 net7.n3756 net7.n3755 0.001
R33451 net7.n3761 net7.n3760 0.001
R33452 net7.n3770 net7.n3769 0.001
R33453 net7.n3880 net7.n3879 0.001
R33454 net7.n3882 net7.n3881 0.001
R33455 net7.n3899 net7.n3898 0.001
R33456 net7.n4032 net7.n4031 0.001
R33457 net7.n4030 net7.n4028 0.001
R33458 net7.n4024 net7.n4023 0.001
R33459 net7.n4019 net7.n4018 0.001
R33460 net7.n4143 net7.n4141 0.001
R33461 net7.n4148 net7.n4145 0.001
R33462 net7.n4156 net7.n4154 0.001
R33463 net7.n4160 net7.n4157 0.001
R33464 net7.n4161 net7.n4160 0.001
R33465 net7.n4163 net7.n4162 0.001
R33466 net7.n4171 net7.n4170 0.001
R33467 net7.n4180 net7.n4176 0.001
R33468 net7.n4309 net7.n4306 0.001
R33469 net7.n4311 net7.n4310 0.001
R33470 net7.n4076 net7.n4075 0.001
R33471 net7.n4082 net7.n4081 0.001
R33472 net7.n4112 net7.n4111 0.001
R33473 net7.n4117 net7.n4116 0.001
R33474 net7.n4122 net7.n4121 0.001
R33475 net7.n4131 net7.n4130 0.001
R33476 net7.n4241 net7.n4240 0.001
R33477 net7.n4243 net7.n4242 0.001
R33478 net7.n4260 net7.n4259 0.001
R33479 net7.n4394 net7.n4393 0.001
R33480 net7.n4392 net7.n4390 0.001
R33481 net7.n4386 net7.n4385 0.001
R33482 net7.n4381 net7.n4380 0.001
R33483 net7.n4505 net7.n4503 0.001
R33484 net7.n4510 net7.n4507 0.001
R33485 net7.n4518 net7.n4516 0.001
R33486 net7.n4522 net7.n4519 0.001
R33487 net7.n4523 net7.n4522 0.001
R33488 net7.n4525 net7.n4524 0.001
R33489 net7.n4533 net7.n4532 0.001
R33490 net7.n4542 net7.n4538 0.001
R33491 net7.n4671 net7.n4668 0.001
R33492 net7.n4673 net7.n4672 0.001
R33493 net7.n4438 net7.n4437 0.001
R33494 net7.n4444 net7.n4443 0.001
R33495 net7.n4474 net7.n4473 0.001
R33496 net7.n4479 net7.n4478 0.001
R33497 net7.n4484 net7.n4483 0.001
R33498 net7.n4493 net7.n4492 0.001
R33499 net7.n4603 net7.n4602 0.001
R33500 net7.n4605 net7.n4604 0.001
R33501 net7.n4622 net7.n4621 0.001
R33502 net7.n4756 net7.n4755 0.001
R33503 net7.n4754 net7.n4752 0.001
R33504 net7.n4748 net7.n4747 0.001
R33505 net7.n4743 net7.n4742 0.001
R33506 net7.n4867 net7.n4865 0.001
R33507 net7.n4872 net7.n4869 0.001
R33508 net7.n4880 net7.n4878 0.001
R33509 net7.n4884 net7.n4881 0.001
R33510 net7.n4885 net7.n4884 0.001
R33511 net7.n4887 net7.n4886 0.001
R33512 net7.n4895 net7.n4894 0.001
R33513 net7.n4904 net7.n4900 0.001
R33514 net7.n5033 net7.n5030 0.001
R33515 net7.n5035 net7.n5034 0.001
R33516 net7.n4800 net7.n4799 0.001
R33517 net7.n4806 net7.n4805 0.001
R33518 net7.n4836 net7.n4835 0.001
R33519 net7.n4841 net7.n4840 0.001
R33520 net7.n4846 net7.n4845 0.001
R33521 net7.n4855 net7.n4854 0.001
R33522 net7.n4965 net7.n4964 0.001
R33523 net7.n4967 net7.n4966 0.001
R33524 net7.n4984 net7.n4983 0.001
R33525 net7.n5118 net7.n5117 0.001
R33526 net7.n5116 net7.n5114 0.001
R33527 net7.n5110 net7.n5109 0.001
R33528 net7.n5105 net7.n5104 0.001
R33529 net7.n5229 net7.n5227 0.001
R33530 net7.n5234 net7.n5231 0.001
R33531 net7.n5242 net7.n5240 0.001
R33532 net7.n5246 net7.n5243 0.001
R33533 net7.n5247 net7.n5246 0.001
R33534 net7.n5249 net7.n5248 0.001
R33535 net7.n5257 net7.n5256 0.001
R33536 net7.n5266 net7.n5262 0.001
R33537 net7.n5395 net7.n5392 0.001
R33538 net7.n5397 net7.n5396 0.001
R33539 net7.n5162 net7.n5161 0.001
R33540 net7.n5168 net7.n5167 0.001
R33541 net7.n5198 net7.n5197 0.001
R33542 net7.n5203 net7.n5202 0.001
R33543 net7.n5208 net7.n5207 0.001
R33544 net7.n5217 net7.n5216 0.001
R33545 net7.n5327 net7.n5326 0.001
R33546 net7.n5329 net7.n5328 0.001
R33547 net7.n5346 net7.n5345 0.001
R33548 net7.n5480 net7.n5479 0.001
R33549 net7.n5478 net7.n5476 0.001
R33550 net7.n5472 net7.n5471 0.001
R33551 net7.n5467 net7.n5466 0.001
R33552 net7.n5591 net7.n5589 0.001
R33553 net7.n5596 net7.n5593 0.001
R33554 net7.n5604 net7.n5602 0.001
R33555 net7.n5608 net7.n5605 0.001
R33556 net7.n5609 net7.n5608 0.001
R33557 net7.n5611 net7.n5610 0.001
R33558 net7.n5619 net7.n5618 0.001
R33559 net7.n5628 net7.n5624 0.001
R33560 net7.n5757 net7.n5754 0.001
R33561 net7.n5759 net7.n5758 0.001
R33562 net7.n5524 net7.n5523 0.001
R33563 net7.n5530 net7.n5529 0.001
R33564 net7.n5560 net7.n5559 0.001
R33565 net7.n5565 net7.n5564 0.001
R33566 net7.n5570 net7.n5569 0.001
R33567 net7.n5579 net7.n5578 0.001
R33568 net7.n5689 net7.n5688 0.001
R33569 net7.n5691 net7.n5690 0.001
R33570 net7.n5708 net7.n5707 0.001
R33571 net7.n5842 net7.n5841 0.001
R33572 net7.n5840 net7.n5838 0.001
R33573 net7.n5834 net7.n5833 0.001
R33574 net7.n5829 net7.n5828 0.001
R33575 net7.n5953 net7.n5951 0.001
R33576 net7.n5958 net7.n5955 0.001
R33577 net7.n5966 net7.n5964 0.001
R33578 net7.n5970 net7.n5967 0.001
R33579 net7.n5971 net7.n5970 0.001
R33580 net7.n5973 net7.n5972 0.001
R33581 net7.n5981 net7.n5980 0.001
R33582 net7.n5990 net7.n5986 0.001
R33583 net7.n6119 net7.n6116 0.001
R33584 net7.n6121 net7.n6120 0.001
R33585 net7.n5886 net7.n5885 0.001
R33586 net7.n5892 net7.n5891 0.001
R33587 net7.n5922 net7.n5921 0.001
R33588 net7.n5927 net7.n5926 0.001
R33589 net7.n5932 net7.n5931 0.001
R33590 net7.n5941 net7.n5940 0.001
R33591 net7.n6051 net7.n6050 0.001
R33592 net7.n6053 net7.n6052 0.001
R33593 net7.n6070 net7.n6069 0.001
R33594 net7.n6204 net7.n6203 0.001
R33595 net7.n6202 net7.n6200 0.001
R33596 net7.n6196 net7.n6195 0.001
R33597 net7.n6191 net7.n6190 0.001
R33598 net7.n6315 net7.n6313 0.001
R33599 net7.n6320 net7.n6317 0.001
R33600 net7.n6328 net7.n6326 0.001
R33601 net7.n6332 net7.n6329 0.001
R33602 net7.n6333 net7.n6332 0.001
R33603 net7.n6335 net7.n6334 0.001
R33604 net7.n6343 net7.n6342 0.001
R33605 net7.n6352 net7.n6348 0.001
R33606 net7.n6481 net7.n6478 0.001
R33607 net7.n6483 net7.n6482 0.001
R33608 net7.n6248 net7.n6247 0.001
R33609 net7.n6254 net7.n6253 0.001
R33610 net7.n6284 net7.n6283 0.001
R33611 net7.n6289 net7.n6288 0.001
R33612 net7.n6294 net7.n6293 0.001
R33613 net7.n6303 net7.n6302 0.001
R33614 net7.n6413 net7.n6412 0.001
R33615 net7.n6415 net7.n6414 0.001
R33616 net7.n6432 net7.n6431 0.001
R33617 net7.n6566 net7.n6565 0.001
R33618 net7.n6564 net7.n6562 0.001
R33619 net7.n6558 net7.n6557 0.001
R33620 net7.n6553 net7.n6552 0.001
R33621 net7.n6677 net7.n6675 0.001
R33622 net7.n6682 net7.n6679 0.001
R33623 net7.n6690 net7.n6688 0.001
R33624 net7.n6694 net7.n6691 0.001
R33625 net7.n6695 net7.n6694 0.001
R33626 net7.n6697 net7.n6696 0.001
R33627 net7.n6705 net7.n6704 0.001
R33628 net7.n6714 net7.n6710 0.001
R33629 net7.n6843 net7.n6840 0.001
R33630 net7.n6845 net7.n6844 0.001
R33631 net7.n6610 net7.n6609 0.001
R33632 net7.n6616 net7.n6615 0.001
R33633 net7.n6646 net7.n6645 0.001
R33634 net7.n6651 net7.n6650 0.001
R33635 net7.n6656 net7.n6655 0.001
R33636 net7.n6665 net7.n6664 0.001
R33637 net7.n6775 net7.n6774 0.001
R33638 net7.n6777 net7.n6776 0.001
R33639 net7.n6794 net7.n6793 0.001
R33640 net7.n6928 net7.n6927 0.001
R33641 net7.n6926 net7.n6924 0.001
R33642 net7.n6920 net7.n6919 0.001
R33643 net7.n6915 net7.n6914 0.001
R33644 net7.n7039 net7.n7037 0.001
R33645 net7.n7044 net7.n7041 0.001
R33646 net7.n7052 net7.n7050 0.001
R33647 net7.n7056 net7.n7053 0.001
R33648 net7.n7057 net7.n7056 0.001
R33649 net7.n7059 net7.n7058 0.001
R33650 net7.n7067 net7.n7066 0.001
R33651 net7.n7076 net7.n7072 0.001
R33652 net7.n7205 net7.n7202 0.001
R33653 net7.n7207 net7.n7206 0.001
R33654 net7.n6972 net7.n6971 0.001
R33655 net7.n6978 net7.n6977 0.001
R33656 net7.n7008 net7.n7007 0.001
R33657 net7.n7013 net7.n7012 0.001
R33658 net7.n7018 net7.n7017 0.001
R33659 net7.n7027 net7.n7026 0.001
R33660 net7.n7137 net7.n7136 0.001
R33661 net7.n7139 net7.n7138 0.001
R33662 net7.n7156 net7.n7155 0.001
R33663 UP.n1 UP.t2 1702.33
R33664 UP.n0 UP.t0 411.601
R33665 UP.n0 UP.t1 236.477
R33666 UP.n1 UP.n0 2.8
R33667 UP UP.n1 0.818
R33668 a_16669_n8264.n20 a_16669_n8264.t2 124.695
R33669 a_16669_n8264.n6 a_16669_n8264.t3 124.695
R33670 a_16669_n8264.n19 a_16669_n8264.n18 92.5
R33671 a_16669_n8264.n5 a_16669_n8264.n4 92.5
R33672 a_16669_n8264.n27 a_16669_n8264.n26 31.034
R33673 a_16669_n8264.n13 a_16669_n8264.n12 31.034
R33674 a_16669_n8264.n33 a_16669_n8264.t1 27.462
R33675 a_16669_n8264.t0 a_16669_n8264.n33 27.245
R33676 a_16669_n8264.n20 a_16669_n8264.n19 15.431
R33677 a_16669_n8264.n6 a_16669_n8264.n5 15.431
R33678 a_16669_n8264.n3 a_16669_n8264.n30 9.3
R33679 a_16669_n8264.n1 a_16669_n8264.n22 9.3
R33680 a_16669_n8264.n1 a_16669_n8264.n21 9.3
R33681 a_16669_n8264.n1 a_16669_n8264.n28 9.3
R33682 a_16669_n8264.n28 a_16669_n8264.n27 9.3
R33683 a_16669_n8264.n3 a_16669_n8264.n29 9.3
R33684 a_16669_n8264.n3 a_16669_n8264.n31 9.3
R33685 a_16669_n8264.n2 a_16669_n8264.n16 9.3
R33686 a_16669_n8264.n0 a_16669_n8264.n8 9.3
R33687 a_16669_n8264.n0 a_16669_n8264.n7 9.3
R33688 a_16669_n8264.n0 a_16669_n8264.n14 9.3
R33689 a_16669_n8264.n14 a_16669_n8264.n13 9.3
R33690 a_16669_n8264.n2 a_16669_n8264.n15 9.3
R33691 a_16669_n8264.n2 a_16669_n8264.n17 9.3
R33692 a_16669_n8264.n28 a_16669_n8264.n24 5.647
R33693 a_16669_n8264.n14 a_16669_n8264.n10 5.647
R33694 a_16669_n8264.n33 a_16669_n8264.n32 5.289
R33695 a_16669_n8264.n32 a_16669_n8264.n2 4.854
R33696 a_16669_n8264.n32 a_16669_n8264.n3 4.839
R33697 a_16669_n8264.n26 a_16669_n8264.n25 4.137
R33698 a_16669_n8264.n12 a_16669_n8264.n11 4.137
R33699 a_16669_n8264.n1 a_16669_n8264.n20 1.57
R33700 a_16669_n8264.n0 a_16669_n8264.n6 1.57
R33701 a_16669_n8264.n24 a_16669_n8264.n23 0.752
R33702 a_16669_n8264.n10 a_16669_n8264.n9 0.752
R33703 a_16669_n8264.n3 a_16669_n8264.n1 0.234
R33704 a_16669_n8264.n2 a_16669_n8264.n0 0.234
R33705 net3.n121 net3.n120 13.176
R33706 net3.n482 net3.n481 13.176
R33707 net3.n921 net3.n920 13.176
R33708 net3.n1282 net3.n1281 13.176
R33709 net3.n155 net3.n154 9.3
R33710 net3.n281 net3.n280 9.3
R33711 net3.n284 net3.n283 9.3
R33712 net3.n292 net3.n291 9.3
R33713 net3.n331 net3.n330 9.3
R33714 net3.n342 net3.n341 9.3
R33715 net3.n333 net3.n332 9.3
R33716 net3.n321 net3.n320 9.3
R33717 net3.n323 net3.n322 9.3
R33718 net3.n295 net3.n294 9.3
R33719 net3.n271 net3.n270 9.3
R33720 net3.n126 net3.n125 9.3
R33721 net3.n157 net3.n156 9.3
R33722 net3.n42 net3.n41 9.3
R33723 net3.n30 net3.n29 9.3
R33724 net3.n28 net3.n27 9.3
R33725 net3.n703 net3.n702 9.3
R33726 net3.n516 net3.n515 9.3
R33727 net3.n642 net3.n641 9.3
R33728 net3.n645 net3.n644 9.3
R33729 net3.n653 net3.n652 9.3
R33730 net3.n692 net3.n691 9.3
R33731 net3.n694 net3.n693 9.3
R33732 net3.n682 net3.n681 9.3
R33733 net3.n684 net3.n683 9.3
R33734 net3.n656 net3.n655 9.3
R33735 net3.n632 net3.n631 9.3
R33736 net3.n487 net3.n486 9.3
R33737 net3.n518 net3.n517 9.3
R33738 net3.n403 net3.n402 9.3
R33739 net3.n391 net3.n390 9.3
R33740 net3.n389 net3.n388 9.3
R33741 net3.n897 net3.n896 9.3
R33742 net3.n778 net3.n777 9.3
R33743 net3.n780 net3.n779 9.3
R33744 net3.n789 net3.n788 9.3
R33745 net3.n771 net3.n770 9.3
R33746 net3.n773 net3.n772 9.3
R33747 net3.n884 net3.n883 9.3
R33748 net3.n926 net3.n925 9.3
R33749 net3.n910 net3.n909 9.3
R33750 net3.n899 net3.n898 9.3
R33751 net3.n886 net3.n885 9.3
R33752 net3.n940 net3.n939 9.3
R33753 net3.n942 net3.n941 9.3
R33754 net3.n1070 net3.n1069 9.3
R33755 net3.n1058 net3.n1057 9.3
R33756 net3.n1056 net3.n1055 9.3
R33757 net3.n1258 net3.n1257 9.3
R33758 net3.n1139 net3.n1138 9.3
R33759 net3.n1141 net3.n1140 9.3
R33760 net3.n1150 net3.n1149 9.3
R33761 net3.n1132 net3.n1131 9.3
R33762 net3.n1134 net3.n1133 9.3
R33763 net3.n1245 net3.n1244 9.3
R33764 net3.n1287 net3.n1286 9.3
R33765 net3.n1271 net3.n1270 9.3
R33766 net3.n1260 net3.n1259 9.3
R33767 net3.n1247 net3.n1246 9.3
R33768 net3.n1301 net3.n1300 9.3
R33769 net3.n1303 net3.n1302 9.3
R33770 net3.n1431 net3.n1430 9.3
R33771 net3.n1419 net3.n1418 9.3
R33772 net3.n1417 net3.n1416 9.3
R33773 net3.n797 net3.n796 8.454
R33774 net3.n1158 net3.n1157 8.454
R33775 net3.n52 net3.n51 8.454
R33776 net3.n413 net3.n412 8.454
R33777 net3.n353 net3.n352 8.454
R33778 net3.n714 net3.n713 8.454
R33779 net3.n1081 net3.n1080 8.453
R33780 net3.n1442 net3.n1441 8.453
R33781 net3.n283 net3.n282 5.458
R33782 net3.n644 net3.n643 5.458
R33783 net3.n896 net3.n895 5.458
R33784 net3.n1257 net3.n1256 5.458
R33785 net3.n154 net3.n153 5.081
R33786 net3.n515 net3.n514 5.081
R33787 net3.n939 net3.n938 5.081
R33788 net3.n1300 net3.n1299 5.081
R33789 net3.n20 net3.n19 4.65
R33790 net3.n147 net3.n146 4.65
R33791 net3.n381 net3.n380 4.65
R33792 net3.n508 net3.n507 4.65
R33793 net3.n1048 net3.n1047 4.65
R33794 net3.n1016 net3.n1015 4.65
R33795 net3.n1409 net3.n1408 4.65
R33796 net3.n1377 net3.n1376 4.65
R33797 net3.n35 net3.n34 4.5
R33798 net3.n311 net3.n310 4.5
R33799 net3.n305 net3.n262 4.5
R33800 net3.n317 net3.n258 4.5
R33801 net3.n327 net3.n326 4.5
R33802 net3.n346 net3.n345 4.5
R33803 net3.n335 net3.n255 4.5
R33804 net3.n301 net3.n300 4.5
R33805 net3.n288 net3.n264 4.5
R33806 net3.n278 net3.n277 4.5
R33807 net3.n268 net3.n266 4.5
R33808 net3.n123 net3.n122 4.5
R33809 net3.n160 net3.n159 4.5
R33810 net3.n141 net3.n132 4.5
R33811 net3.n89 net3.n86 4.5
R33812 net3.n137 net3.n136 4.5
R33813 net3.n16 net3.n15 4.5
R33814 net3.n46 net3.n45 4.5
R33815 net3.n396 net3.n395 4.5
R33816 net3.n672 net3.n671 4.5
R33817 net3.n666 net3.n623 4.5
R33818 net3.n678 net3.n619 4.5
R33819 net3.n688 net3.n687 4.5
R33820 net3.n696 net3.n616 4.5
R33821 net3.n662 net3.n661 4.5
R33822 net3.n649 net3.n625 4.5
R33823 net3.n639 net3.n638 4.5
R33824 net3.n629 net3.n627 4.5
R33825 net3.n484 net3.n483 4.5
R33826 net3.n521 net3.n520 4.5
R33827 net3.n502 net3.n493 4.5
R33828 net3.n450 net3.n447 4.5
R33829 net3.n498 net3.n497 4.5
R33830 net3.n377 net3.n376 4.5
R33831 net3.n407 net3.n406 4.5
R33832 net3.n707 net3.n706 4.5
R33833 net3.n1063 net3.n1062 4.5
R33834 net3.n1044 net3.n1043 4.5
R33835 net3.n1036 net3.n1035 4.5
R33836 net3.n1022 net3.n1021 4.5
R33837 net3.n943 net3.n931 4.5
R33838 net3.n923 net3.n922 4.5
R33839 net3.n913 net3.n912 4.5
R33840 net3.n903 net3.n902 4.5
R33841 net3.n891 net3.n890 4.5
R33842 net3.n774 net3.n740 4.5
R33843 net3.n767 net3.n743 4.5
R33844 net3.n782 net3.n737 4.5
R33845 net3.n791 net3.n734 4.5
R33846 net3.n761 net3.n746 4.5
R33847 net3.n758 net3.n750 4.5
R33848 net3.n754 net3.n753 4.5
R33849 net3.n1030 net3.n1029 4.5
R33850 net3.n1074 net3.n1073 4.5
R33851 net3.n1424 net3.n1423 4.5
R33852 net3.n1405 net3.n1404 4.5
R33853 net3.n1397 net3.n1396 4.5
R33854 net3.n1383 net3.n1382 4.5
R33855 net3.n1304 net3.n1292 4.5
R33856 net3.n1284 net3.n1283 4.5
R33857 net3.n1274 net3.n1273 4.5
R33858 net3.n1264 net3.n1263 4.5
R33859 net3.n1252 net3.n1251 4.5
R33860 net3.n1135 net3.n1101 4.5
R33861 net3.n1128 net3.n1104 4.5
R33862 net3.n1143 net3.n1098 4.5
R33863 net3.n1152 net3.n1095 4.5
R33864 net3.n1122 net3.n1107 4.5
R33865 net3.n1119 net3.n1111 4.5
R33866 net3.n1115 net3.n1114 4.5
R33867 net3.n1391 net3.n1390 4.5
R33868 net3.n1435 net3.n1434 4.5
R33869 net3.n258 net3.n256 4.325
R33870 net3.n619 net3.n617 4.325
R33871 net3.n743 net3.n741 4.325
R33872 net3.n1104 net3.n1102 4.325
R33873 net3.n351 net3.t1 4.289
R33874 net3.n712 net3.t0 4.289
R33875 net3.n1079 net3.t3 4.289
R33876 net3.n1440 net3.t2 4.289
R33877 net3.n262 net3.n259 3.95
R33878 net3.n623 net3.n620 3.95
R33879 net3.n750 net3.n747 3.95
R33880 net3.n1111 net3.n1108 3.95
R33881 net3.n15 net3.n14 3.948
R33882 net3.n376 net3.n375 3.948
R33883 net3.n1043 net3.n1042 3.948
R33884 net3.n1404 net3.n1403 3.948
R33885 net3.n136 net3.n135 3.573
R33886 net3.n497 net3.n496 3.573
R33887 net3.n1029 net3.n1028 3.573
R33888 net3.n1390 net3.n1389 3.573
R33889 net3.n722 net3.n360 3.343
R33890 net3.n149 net3.n130 3.033
R33891 net3.n24 net3.n23 3.033
R33892 net3.n510 net3.n491 3.033
R33893 net3.n385 net3.n384 3.033
R33894 net3.n934 net3.n932 3.033
R33895 net3.n1052 net3.n1051 3.033
R33896 net3.n1295 net3.n1293 3.033
R33897 net3.n1413 net3.n1412 3.033
R33898 net3.n722 net3.n721 2.795
R33899 net3 net3.n722 2.662
R33900 net3.n261 net3.n260 2.258
R33901 net3.n134 net3.n133 2.258
R33902 net3.n622 net3.n621 2.258
R33903 net3.n495 net3.n494 2.258
R33904 net3.n749 net3.n748 2.258
R33905 net3.n1027 net3.n1026 2.258
R33906 net3.n1110 net3.n1109 2.258
R33907 net3.n1388 net3.n1387 2.258
R33908 net3.n309 net3.n308 1.882
R33909 net3.n310 net3.n309 1.882
R33910 net3.n85 net3.n84 1.882
R33911 net3.n670 net3.n669 1.882
R33912 net3.n671 net3.n670 1.882
R33913 net3.n446 net3.n445 1.882
R33914 net3.n745 net3.n744 1.882
R33915 net3.n746 net3.n745 1.882
R33916 net3.n1034 net3.n1033 1.882
R33917 net3.n1106 net3.n1105 1.882
R33918 net3.n1107 net3.n1106 1.882
R33919 net3.n1395 net3.n1394 1.882
R33920 net3.n352 net3.n351 1.844
R33921 net3.n713 net3.n712 1.844
R33922 net3.n1080 net3.n1079 1.844
R33923 net3.n1441 net3.n1440 1.844
R33924 net3.n1445 net3.n1083 1.612
R33925 net3.n136 net3.n134 1.505
R33926 net3.n86 net3.n85 1.505
R33927 net3.n497 net3.n495 1.505
R33928 net3.n447 net3.n446 1.505
R33929 net3.n1029 net3.n1027 1.505
R33930 net3.n1035 net3.n1034 1.505
R33931 net3.n1390 net3.n1388 1.505
R33932 net3.n1396 net3.n1395 1.505
R33933 net3.n1445 net3.n1444 1.292
R33934 net3.n112 net3.n111 1.137
R33935 net3.n190 net3.n189 1.137
R33936 net3.n197 net3.n196 1.137
R33937 net3.n201 net3.n200 1.137
R33938 net3.n208 net3.n207 1.137
R33939 net3.n226 net3.n225 1.137
R33940 net3.n243 net3.n242 1.137
R33941 net3.n250 net3.n249 1.137
R33942 net3.n239 net3.n238 1.137
R33943 net3.n232 net3.n231 1.137
R33944 net3.n218 net3.n217 1.137
R33945 net3.n182 net3.n181 1.137
R33946 net3.n173 net3.n172 1.137
R33947 net3.n164 net3.n163 1.137
R33948 net3.n101 net3.n100 1.137
R33949 net3.n108 net3.n107 1.137
R33950 net3.n93 net3.n92 1.137
R33951 net3.n78 net3.n77 1.137
R33952 net3.n62 net3.n61 1.137
R33953 net3.n69 net3.n68 1.137
R33954 net3.n360 net3.n359 1.137
R33955 net3.n721 net3.n720 1.137
R33956 net3.n473 net3.n472 1.137
R33957 net3.n551 net3.n550 1.137
R33958 net3.n558 net3.n557 1.137
R33959 net3.n562 net3.n561 1.137
R33960 net3.n569 net3.n568 1.137
R33961 net3.n587 net3.n586 1.137
R33962 net3.n604 net3.n603 1.137
R33963 net3.n600 net3.n599 1.137
R33964 net3.n593 net3.n592 1.137
R33965 net3.n579 net3.n578 1.137
R33966 net3.n543 net3.n542 1.137
R33967 net3.n534 net3.n533 1.137
R33968 net3.n525 net3.n524 1.137
R33969 net3.n462 net3.n461 1.137
R33970 net3.n469 net3.n468 1.137
R33971 net3.n454 net3.n453 1.137
R33972 net3.n439 net3.n438 1.137
R33973 net3.n423 net3.n422 1.137
R33974 net3.n430 net3.n429 1.137
R33975 net3.n611 net3.n610 1.137
R33976 net3.n998 net3.n997 1.137
R33977 net3.n1006 net3.n1005 1.137
R33978 net3.n956 net3.n955 1.137
R33979 net3.n849 net3.n848 1.137
R33980 net3.n821 net3.n820 1.137
R33981 net3.n807 net3.n806 1.137
R33982 net3.n813 net3.n812 1.137
R33983 net3.n830 net3.n829 1.137
R33984 net3.n845 net3.n844 1.137
R33985 net3.n838 net3.n837 1.137
R33986 net3.n856 net3.n855 1.137
R33987 net3.n866 net3.n865 1.137
R33988 net3.n952 net3.n951 1.137
R33989 net3.n875 net3.n874 1.137
R33990 net3.n945 net3.n944 1.137
R33991 net3.n963 net3.n962 1.137
R33992 net3.n973 net3.n972 1.137
R33993 net3.n979 net3.n978 1.137
R33994 net3.n994 net3.n993 1.137
R33995 net3.n987 net3.n986 1.137
R33996 net3.n1083 net3.n1082 1.137
R33997 net3.n1359 net3.n1358 1.137
R33998 net3.n1367 net3.n1366 1.137
R33999 net3.n1317 net3.n1316 1.137
R34000 net3.n1210 net3.n1209 1.137
R34001 net3.n1182 net3.n1181 1.137
R34002 net3.n1168 net3.n1167 1.137
R34003 net3.n1174 net3.n1173 1.137
R34004 net3.n1191 net3.n1190 1.137
R34005 net3.n1206 net3.n1205 1.137
R34006 net3.n1199 net3.n1198 1.137
R34007 net3.n1217 net3.n1216 1.137
R34008 net3.n1227 net3.n1226 1.137
R34009 net3.n1313 net3.n1312 1.137
R34010 net3.n1236 net3.n1235 1.137
R34011 net3.n1306 net3.n1305 1.137
R34012 net3.n1324 net3.n1323 1.137
R34013 net3.n1334 net3.n1333 1.137
R34014 net3.n1340 net3.n1339 1.137
R34015 net3.n1355 net3.n1354 1.137
R34016 net3.n1348 net3.n1347 1.137
R34017 net3.n1444 net3.n1443 1.137
R34018 net3.n255 net3.n254 1.129
R34019 net3.n262 net3.n261 1.129
R34020 net3.n300 net3.n299 1.129
R34021 net3.n616 net3.n615 1.129
R34022 net3.n623 net3.n622 1.129
R34023 net3.n661 net3.n660 1.129
R34024 net3.n737 net3.n736 1.129
R34025 net3.n750 net3.n749 1.129
R34026 net3.n753 net3.n752 1.129
R34027 net3.n1098 net3.n1097 1.129
R34028 net3.n1111 net3.n1110 1.129
R34029 net3.n1114 net3.n1113 1.129
R34030 net3.n90 net3.n89 1.125
R34031 net3.n451 net3.n450 1.125
R34032 net3.n163 net3.n160 1.042
R34033 net3.n524 net3.n521 1.042
R34034 net3.n944 net3.n943 1.042
R34035 net3.n1305 net3.n1304 1.042
R34036 net3.n54 net3.n53 0.869
R34037 net3.n415 net3.n414 0.869
R34038 net3.n799 net3.n798 0.869
R34039 net3.n1160 net3.n1159 0.869
R34040 net3.n345 net3.n344 0.752
R34041 net3.n159 net3.n158 0.752
R34042 net3.n132 net3.n131 0.752
R34043 net3.n15 net3.n13 0.752
R34044 net3.n34 net3.n33 0.752
R34045 net3.n45 net3.n44 0.752
R34046 net3.n706 net3.n705 0.752
R34047 net3.n520 net3.n519 0.752
R34048 net3.n493 net3.n492 0.752
R34049 net3.n376 net3.n374 0.752
R34050 net3.n395 net3.n394 0.752
R34051 net3.n406 net3.n405 0.752
R34052 net3.n734 net3.n733 0.752
R34053 net3.n931 net3.n930 0.752
R34054 net3.n1021 net3.n1020 0.752
R34055 net3.n1043 net3.n1041 0.752
R34056 net3.n1062 net3.n1061 0.752
R34057 net3.n1073 net3.n1072 0.752
R34058 net3.n1095 net3.n1094 0.752
R34059 net3.n1292 net3.n1291 0.752
R34060 net3.n1382 net3.n1381 0.752
R34061 net3.n1404 net3.n1402 0.752
R34062 net3.n1423 net3.n1422 0.752
R34063 net3.n1434 net3.n1433 0.752
R34064 net3.n798 net3.n797 0.729
R34065 net3.n1159 net3.n1158 0.729
R34066 net3.n53 net3.n52 0.728
R34067 net3.n414 net3.n413 0.728
R34068 net3.n1082 net3.n1081 0.725
R34069 net3.n1443 net3.n1442 0.725
R34070 net3.n359 net3.n353 0.725
R34071 net3.n720 net3.n714 0.725
R34072 net3.n326 net3.n325 0.376
R34073 net3.n258 net3.n257 0.376
R34074 net3.n264 net3.n263 0.376
R34075 net3.n277 net3.n276 0.376
R34076 net3.n266 net3.n265 0.376
R34077 net3.n122 net3.n121 0.376
R34078 net3.n687 net3.n686 0.376
R34079 net3.n619 net3.n618 0.376
R34080 net3.n625 net3.n624 0.376
R34081 net3.n638 net3.n637 0.376
R34082 net3.n627 net3.n626 0.376
R34083 net3.n483 net3.n482 0.376
R34084 net3.n740 net3.n739 0.376
R34085 net3.n743 net3.n742 0.376
R34086 net3.n890 net3.n889 0.376
R34087 net3.n902 net3.n901 0.376
R34088 net3.n912 net3.n911 0.376
R34089 net3.n922 net3.n921 0.376
R34090 net3.n1101 net3.n1100 0.376
R34091 net3.n1104 net3.n1103 0.376
R34092 net3.n1251 net3.n1250 0.376
R34093 net3.n1263 net3.n1262 0.376
R34094 net3.n1273 net3.n1272 0.376
R34095 net3.n1283 net3.n1282 0.376
R34096 net3 net3.n1445 0.317
R34097 net3.n125 net3.n124 0.189
R34098 net3.n486 net3.n485 0.189
R34099 net3.n909 net3.n908 0.189
R34100 net3.n925 net3.n924 0.189
R34101 net3.n1270 net3.n1269 0.189
R34102 net3.n1286 net3.n1285 0.189
R34103 net3.n270 net3.n269 0.188
R34104 net3.n631 net3.n630 0.188
R34105 net3.n146 net3.n145 0.166
R34106 net3.n507 net3.n506 0.166
R34107 net3.n883 net3.n882 0.166
R34108 net3.n1015 net3.n1014 0.166
R34109 net3.n1244 net3.n1243 0.166
R34110 net3.n1376 net3.n1375 0.166
R34111 net3.n294 net3.n293 0.166
R34112 net3.n655 net3.n654 0.166
R34113 net3.n23 net3.n22 0.133
R34114 net3.n384 net3.n383 0.133
R34115 net3.n325 net3.n324 0.132
R34116 net3.n686 net3.n685 0.132
R34117 net3.n739 net3.n738 0.132
R34118 net3.n1051 net3.n1050 0.132
R34119 net3.n1100 net3.n1099 0.132
R34120 net3.n1412 net3.n1411 0.132
R34121 net3.n33 net3.n32 0.121
R34122 net3.n394 net3.n393 0.121
R34123 net3.n736 net3.n735 0.121
R34124 net3.n1061 net3.n1060 0.121
R34125 net3.n1097 net3.n1096 0.121
R34126 net3.n1422 net3.n1421 0.121
R34127 net3.n254 net3.n253 0.121
R34128 net3.n615 net3.n614 0.121
R34129 net3.n231 net3.n230 0.049
R34130 net3.n226 net3.n218 0.049
R34131 net3.n182 net3.n173 0.049
R34132 net3.n93 net3.n78 0.049
R34133 net3.n592 net3.n591 0.049
R34134 net3.n587 net3.n579 0.049
R34135 net3.n543 net3.n534 0.049
R34136 net3.n454 net3.n439 0.049
R34137 net3.n944 net3.n879 0.049
R34138 net3.n830 net3.n821 0.049
R34139 net3.n875 net3.n866 0.049
R34140 net3.n979 net3.n973 0.049
R34141 net3.n1305 net3.n1240 0.049
R34142 net3.n1191 net3.n1182 0.049
R34143 net3.n1236 net3.n1227 0.049
R34144 net3.n1340 net3.n1334 0.049
R34145 net3.n350 net3.n349 0.047
R34146 net3.n331 net3.n329 0.047
R34147 net3.n329 net3.n328 0.047
R34148 net3.n321 net3.n319 0.047
R34149 net3.n273 net3.n272 0.047
R34150 net3.n128 net3.n127 0.047
R34151 net3.n20 net3.n18 0.047
R34152 net3.n25 net3.n24 0.047
R34153 net3.n28 net3.n26 0.047
R34154 net3.n50 net3.n49 0.047
R34155 net3.n188 net3.n187 0.047
R34156 net3.n711 net3.n710 0.047
R34157 net3.n692 net3.n690 0.047
R34158 net3.n690 net3.n689 0.047
R34159 net3.n682 net3.n680 0.047
R34160 net3.n634 net3.n633 0.047
R34161 net3.n489 net3.n488 0.047
R34162 net3.n381 net3.n379 0.047
R34163 net3.n386 net3.n385 0.047
R34164 net3.n389 net3.n387 0.047
R34165 net3.n411 net3.n410 0.047
R34166 net3.n549 net3.n548 0.047
R34167 net3.n795 net3.n794 0.047
R34168 net3.n778 net3.n776 0.047
R34169 net3.n776 net3.n775 0.047
R34170 net3.n771 net3.n769 0.047
R34171 net3.n907 net3.n906 0.047
R34172 net3.n928 net3.n927 0.047
R34173 net3.n1048 net3.n1046 0.047
R34174 net3.n1053 net3.n1052 0.047
R34175 net3.n1056 net3.n1054 0.047
R34176 net3.n1078 net3.n1077 0.047
R34177 net3.n986 net3.n984 0.047
R34178 net3.n1156 net3.n1155 0.047
R34179 net3.n1139 net3.n1137 0.047
R34180 net3.n1137 net3.n1136 0.047
R34181 net3.n1132 net3.n1130 0.047
R34182 net3.n1268 net3.n1267 0.047
R34183 net3.n1289 net3.n1288 0.047
R34184 net3.n1409 net3.n1407 0.047
R34185 net3.n1414 net3.n1413 0.047
R34186 net3.n1417 net3.n1415 0.047
R34187 net3.n1439 net3.n1438 0.047
R34188 net3.n1347 net3.n1345 0.047
R34189 net3.n275 net3.n274 0.045
R34190 net3.n129 net3.n128 0.045
R34191 net3.n636 net3.n635 0.045
R34192 net3.n490 net3.n489 0.045
R34193 net3.n905 net3.n904 0.045
R34194 net3.n929 net3.n928 0.045
R34195 net3.n1266 net3.n1265 0.045
R34196 net3.n1290 net3.n1289 0.045
R34197 net3.n298 net3.n297 0.043
R34198 net3.n89 net3.n83 0.043
R34199 net3.n181 net3.n180 0.043
R34200 net3.n91 net3.n90 0.043
R34201 net3.n76 net3.n75 0.043
R34202 net3.n659 net3.n658 0.043
R34203 net3.n450 net3.n444 0.043
R34204 net3.n542 net3.n541 0.043
R34205 net3.n452 net3.n451 0.043
R34206 net3.n437 net3.n436 0.043
R34207 net3.n915 net3.n914 0.043
R34208 net3.n1036 net3.n1032 0.043
R34209 net3.n818 net3.n817 0.043
R34210 net3.n836 net3.n835 0.043
R34211 net3.n1276 net3.n1275 0.043
R34212 net3.n1397 net3.n1393 0.043
R34213 net3.n1179 net3.n1178 0.043
R34214 net3.n1197 net3.n1196 0.043
R34215 net3.n353 net3.n350 0.043
R34216 net3.n714 net3.n711 0.043
R34217 net3.n797 net3.n795 0.043
R34218 net3.n1158 net3.n1156 0.043
R34219 net3.n318 net3.n317 0.041
R34220 net3.n311 net3.n307 0.041
R34221 net3.n119 net3.n118 0.041
R34222 net3.n143 net3.n142 0.041
R34223 net3.n40 net3.n39 0.041
R34224 net3.n225 net3.n224 0.041
R34225 net3.n99 net3.n98 0.041
R34226 net3.n679 net3.n678 0.041
R34227 net3.n672 net3.n668 0.041
R34228 net3.n480 net3.n479 0.041
R34229 net3.n504 net3.n503 0.041
R34230 net3.n401 net3.n400 0.041
R34231 net3.n586 net3.n585 0.041
R34232 net3.n460 net3.n459 0.041
R34233 net3.n768 net3.n767 0.041
R34234 net3.n761 net3.n760 0.041
R34235 net3.n919 net3.n918 0.041
R34236 net3.n1019 net3.n1018 0.041
R34237 net3.n1068 net3.n1067 0.041
R34238 net3.n826 net3.n825 0.041
R34239 net3.n874 net3.n870 0.041
R34240 net3.n1129 net3.n1128 0.041
R34241 net3.n1122 net3.n1121 0.041
R34242 net3.n1280 net3.n1279 0.041
R34243 net3.n1380 net3.n1379 0.041
R34244 net3.n1429 net3.n1428 0.041
R34245 net3.n1187 net3.n1186 0.041
R34246 net3.n1235 net3.n1231 0.041
R34247 net3.n1081 net3.n1078 0.041
R34248 net3.n1442 net3.n1439 0.041
R34249 net3.n52 net3.n50 0.041
R34250 net3.n413 net3.n411 0.041
R34251 net3.n340 net3.n339 0.039
R34252 net3.n296 net3.n295 0.039
R34253 net3.n147 net3.n144 0.039
R34254 net3.n17 net3.n16 0.039
R34255 net3.n77 net3.n72 0.039
R34256 net3.n701 net3.n700 0.039
R34257 net3.n657 net3.n656 0.039
R34258 net3.n508 net3.n505 0.039
R34259 net3.n378 net3.n377 0.039
R34260 net3.n438 net3.n433 0.039
R34261 net3.n787 net3.n786 0.039
R34262 net3.n884 net3.n881 0.039
R34263 net3.n1017 net3.n1016 0.039
R34264 net3.n1045 net3.n1044 0.039
R34265 net3.n978 net3.n976 0.039
R34266 net3.n1148 net3.n1147 0.039
R34267 net3.n1245 net3.n1242 0.039
R34268 net3.n1378 net3.n1377 0.039
R34269 net3.n1406 net3.n1405 0.039
R34270 net3.n1339 net3.n1337 0.039
R34271 net3.n306 net3.n305 0.037
R34272 net3.n667 net3.n666 0.037
R34273 net3.n759 net3.n758 0.037
R34274 net3.n1120 net3.n1119 0.037
R34275 net3.n7 net3.n6 0.035
R34276 net3.n368 net3.n367 0.035
R34277 net3.n1031 net3.n1030 0.035
R34278 net3.n729 net3.n728 0.035
R34279 net3.n1392 net3.n1391 0.035
R34280 net3.n1090 net3.n1089 0.035
R34281 net3.n285 net3.n284 0.034
R34282 net3.n117 net3.n116 0.034
R34283 net3.n230 net3.n229 0.034
R34284 net3.n223 net3.n222 0.034
R34285 net3.n179 net3.n178 0.034
R34286 net3.n168 net3.n167 0.034
R34287 net3.n90 net3.n81 0.034
R34288 net3.n75 net3.n74 0.034
R34289 net3.n646 net3.n645 0.034
R34290 net3.n478 net3.n477 0.034
R34291 net3.n591 net3.n590 0.034
R34292 net3.n584 net3.n583 0.034
R34293 net3.n540 net3.n539 0.034
R34294 net3.n529 net3.n528 0.034
R34295 net3.n451 net3.n442 0.034
R34296 net3.n436 net3.n435 0.034
R34297 net3.n897 net3.n894 0.034
R34298 net3.n917 net3.n916 0.034
R34299 net3.n817 net3.n816 0.034
R34300 net3.n824 net3.n823 0.034
R34301 net3.n869 net3.n868 0.034
R34302 net3.n879 net3.n878 0.034
R34303 net3.n975 net3.n974 0.034
R34304 net3.n983 net3.n982 0.034
R34305 net3.n1258 net3.n1255 0.034
R34306 net3.n1278 net3.n1277 0.034
R34307 net3.n1178 net3.n1177 0.034
R34308 net3.n1185 net3.n1184 0.034
R34309 net3.n1230 net3.n1229 0.034
R34310 net3.n1240 net3.n1239 0.034
R34311 net3.n1336 net3.n1335 0.034
R34312 net3.n1344 net3.n1343 0.034
R34313 net3.n348 net3.n347 0.032
R34314 net3.n155 net3.n152 0.032
R34315 net3.n48 net3.n47 0.032
R34316 net3.n186 net3.n185 0.032
R34317 net3.n709 net3.n708 0.032
R34318 net3.n516 net3.n513 0.032
R34319 net3.n409 net3.n408 0.032
R34320 net3.n547 net3.n546 0.032
R34321 net3.n793 net3.n792 0.032
R34322 net3.n940 net3.n937 0.032
R34323 net3.n1076 net3.n1075 0.032
R34324 net3.n861 net3.n860 0.032
R34325 net3.n1154 net3.n1153 0.032
R34326 net3.n1301 net3.n1298 0.032
R34327 net3.n1437 net3.n1436 0.032
R34328 net3.n1222 net3.n1221 0.032
R34329 net3.n251 net3.n250 0.031
R34330 net3.n232 net3.n228 0.031
R34331 net3.n209 net3.n208 0.031
R34332 net3.n190 net3.n184 0.031
R34333 net3.n165 net3.n164 0.031
R34334 net3.n101 net3.n95 0.031
R34335 net3.n70 net3.n69 0.031
R34336 net3.n55 net3.n54 0.031
R34337 net3.n612 net3.n611 0.031
R34338 net3.n593 net3.n589 0.031
R34339 net3.n570 net3.n569 0.031
R34340 net3.n551 net3.n545 0.031
R34341 net3.n526 net3.n525 0.031
R34342 net3.n462 net3.n456 0.031
R34343 net3.n431 net3.n430 0.031
R34344 net3.n416 net3.n415 0.031
R34345 net3.n800 net3.n799 0.031
R34346 net3.n814 net3.n813 0.031
R34347 net3.n838 net3.n832 0.031
R34348 net3.n857 net3.n856 0.031
R34349 net3.n945 net3.n877 0.031
R34350 net3.n964 net3.n963 0.031
R34351 net3.n987 net3.n981 0.031
R34352 net3.n1007 net3.n1006 0.031
R34353 net3.n1161 net3.n1160 0.031
R34354 net3.n1175 net3.n1174 0.031
R34355 net3.n1199 net3.n1193 0.031
R34356 net3.n1218 net3.n1217 0.031
R34357 net3.n1306 net3.n1238 0.031
R34358 net3.n1325 net3.n1324 0.031
R34359 net3.n1348 net3.n1342 0.031
R34360 net3.n1368 net3.n1367 0.031
R34361 net3.n327 net3.n323 0.03
R34362 net3.n271 net3.n268 0.03
R34363 net3.n126 net3.n123 0.03
R34364 net3.n21 net3.n20 0.03
R34365 net3.n38 net3.n37 0.03
R34366 net3.n170 net3.n169 0.03
R34367 net3.n688 net3.n684 0.03
R34368 net3.n632 net3.n629 0.03
R34369 net3.n487 net3.n484 0.03
R34370 net3.n382 net3.n381 0.03
R34371 net3.n399 net3.n398 0.03
R34372 net3.n531 net3.n530 0.03
R34373 net3.n774 net3.n773 0.03
R34374 net3.n913 net3.n910 0.03
R34375 net3.n926 net3.n923 0.03
R34376 net3.n1049 net3.n1048 0.03
R34377 net3.n1066 net3.n1065 0.03
R34378 net3.n872 net3.n871 0.03
R34379 net3.n996 net3.n995 0.03
R34380 net3.n1135 net3.n1134 0.03
R34381 net3.n1274 net3.n1271 0.03
R34382 net3.n1287 net3.n1284 0.03
R34383 net3.n1410 net3.n1409 0.03
R34384 net3.n1427 net3.n1426 0.03
R34385 net3.n1233 net3.n1232 0.03
R34386 net3.n1357 net3.n1356 0.03
R34387 net3.n798 net3.n732 0.029
R34388 net3.n1159 net3.n1093 0.029
R34389 net3.n338 net3.n337 0.028
R34390 net3.n281 net3.n279 0.028
R34391 net3.n160 net3.n157 0.028
R34392 net3.n150 net3.n149 0.028
R34393 net3.n241 net3.n240 0.028
R34394 net3.n216 net3.n215 0.028
R34395 net3.n214 net3.n213 0.028
R34396 net3.n175 net3.n174 0.028
R34397 net3.n699 net3.n698 0.028
R34398 net3.n642 net3.n640 0.028
R34399 net3.n521 net3.n518 0.028
R34400 net3.n511 net3.n510 0.028
R34401 net3.n602 net3.n601 0.028
R34402 net3.n577 net3.n576 0.028
R34403 net3.n575 net3.n574 0.028
R34404 net3.n536 net3.n535 0.028
R34405 net3.n785 net3.n784 0.028
R34406 net3.n900 net3.n899 0.028
R34407 net3.n943 net3.n942 0.028
R34408 net3.n935 net3.n934 0.028
R34409 net3.n828 net3.n827 0.028
R34410 net3.n834 net3.n833 0.028
R34411 net3.n863 net3.n862 0.028
R34412 net3.n954 net3.n953 0.028
R34413 net3.n1146 net3.n1145 0.028
R34414 net3.n1261 net3.n1260 0.028
R34415 net3.n1304 net3.n1303 0.028
R34416 net3.n1296 net3.n1295 0.028
R34417 net3.n1189 net3.n1188 0.028
R34418 net3.n1195 net3.n1194 0.028
R34419 net3.n1224 net3.n1223 0.028
R34420 net3.n1315 net3.n1314 0.028
R34421 net3.n53 net3.n10 0.027
R34422 net3.n414 net3.n371 0.027
R34423 net3.n243 net3.n239 0.027
R34424 net3.n201 net3.n197 0.027
R34425 net3.n112 net3.n108 0.027
R34426 net3.n62 net3.n58 0.027
R34427 net3.n604 net3.n600 0.027
R34428 net3.n562 net3.n558 0.027
R34429 net3.n473 net3.n469 0.027
R34430 net3.n423 net3.n419 0.027
R34431 net3.n807 net3.n803 0.027
R34432 net3.n849 net3.n845 0.027
R34433 net3.n956 net3.n952 0.027
R34434 net3.n998 net3.n994 0.027
R34435 net3.n1168 net3.n1164 0.027
R34436 net3.n1210 net3.n1206 0.027
R34437 net3.n1317 net3.n1313 0.027
R34438 net3.n1359 net3.n1355 0.027
R34439 net3.n288 net3.n287 0.026
R34440 net3.n356 net3.n355 0.026
R34441 net3.n199 net3.n198 0.026
R34442 net3.n97 net3.n96 0.026
R34443 net3.n80 net3.n79 0.026
R34444 net3.n649 net3.n648 0.026
R34445 net3.n717 net3.n716 0.026
R34446 net3.n560 net3.n559 0.026
R34447 net3.n458 net3.n457 0.026
R34448 net3.n441 net3.n440 0.026
R34449 net3.n892 net3.n891 0.026
R34450 net3.n731 net3.n730 0.026
R34451 net3.n968 net3.n967 0.026
R34452 net3.n970 net3.n969 0.026
R34453 net3.n1253 net3.n1252 0.026
R34454 net3.n1092 net3.n1091 0.026
R34455 net3.n1329 net3.n1328 0.026
R34456 net3.n1331 net3.n1330 0.026
R34457 net3.n148 net3.n147 0.024
R34458 net3.n249 net3.n248 0.024
R34459 net3.n238 net3.n237 0.024
R34460 net3.n207 net3.n206 0.024
R34461 net3.n196 net3.n195 0.024
R34462 net3.n163 net3.n162 0.024
R34463 net3.n107 net3.n106 0.024
R34464 net3.n2 net3.n1 0.024
R34465 net3.n9 net3.n8 0.024
R34466 net3.n509 net3.n508 0.024
R34467 net3.n610 net3.n609 0.024
R34468 net3.n599 net3.n598 0.024
R34469 net3.n568 net3.n567 0.024
R34470 net3.n557 net3.n556 0.024
R34471 net3.n524 net3.n523 0.024
R34472 net3.n468 net3.n467 0.024
R34473 net3.n363 net3.n362 0.024
R34474 net3.n370 net3.n369 0.024
R34475 net3.n727 net3.n726 0.024
R34476 net3.n725 net3.n724 0.024
R34477 net3.n812 net3.n811 0.024
R34478 net3.n844 net3.n842 0.024
R34479 net3.n855 net3.n853 0.024
R34480 net3.n951 net3.n949 0.024
R34481 net3.n962 net3.n960 0.024
R34482 net3.n993 net3.n991 0.024
R34483 net3.n1011 net3.n1010 0.024
R34484 net3.n1088 net3.n1087 0.024
R34485 net3.n1086 net3.n1085 0.024
R34486 net3.n1173 net3.n1172 0.024
R34487 net3.n1205 net3.n1203 0.024
R34488 net3.n1216 net3.n1214 0.024
R34489 net3.n1312 net3.n1310 0.024
R34490 net3.n1323 net3.n1321 0.024
R34491 net3.n1354 net3.n1352 0.024
R34492 net3.n1372 net3.n1371 0.024
R34493 net3.n292 net3.n290 0.022
R34494 net3.n287 net3.n286 0.022
R34495 net3.n358 net3.n357 0.022
R34496 net3.n67 net3.n66 0.022
R34497 net3.n5 net3.n4 0.022
R34498 net3.n10 net3.n9 0.022
R34499 net3.n653 net3.n651 0.022
R34500 net3.n648 net3.n647 0.022
R34501 net3.n719 net3.n718 0.022
R34502 net3.n428 net3.n427 0.022
R34503 net3.n366 net3.n365 0.022
R34504 net3.n371 net3.n370 0.022
R34505 net3.n887 net3.n886 0.022
R34506 net3.n893 net3.n892 0.022
R34507 net3.n847 net3.n846 0.022
R34508 net3.n1005 net3.n1003 0.022
R34509 net3.n1012 net3.n1011 0.022
R34510 net3.n1248 net3.n1247 0.022
R34511 net3.n1254 net3.n1253 0.022
R34512 net3.n1208 net3.n1207 0.022
R34513 net3.n1366 net3.n1364 0.022
R34514 net3.n1373 net3.n1372 0.022
R34515 net3.n303 net3.n302 0.02
R34516 net3.n151 net3.n150 0.02
R34517 net3.n140 net3.n139 0.02
R34518 net3.n357 net3.n356 0.02
R34519 net3.n110 net3.n109 0.02
R34520 net3.n664 net3.n663 0.02
R34521 net3.n512 net3.n511 0.02
R34522 net3.n501 net3.n500 0.02
R34523 net3.n718 net3.n717 0.02
R34524 net3.n471 net3.n470 0.02
R34525 net3.n756 net3.n755 0.02
R34526 net3.n936 net3.n935 0.02
R34527 net3.n1024 net3.n1023 0.02
R34528 net3.n732 net3.n731 0.02
R34529 net3.n805 net3.n804 0.02
R34530 net3.n1013 net3.n1012 0.02
R34531 net3.n1117 net3.n1116 0.02
R34532 net3.n1297 net3.n1296 0.02
R34533 net3.n1385 net3.n1384 0.02
R34534 net3.n1093 net3.n1092 0.02
R34535 net3.n1166 net3.n1165 0.02
R34536 net3.n1374 net3.n1373 0.02
R34537 net3.n60 net3.n59 0.018
R34538 net3.n421 net3.n420 0.018
R34539 net3.n315 net3.n314 0.017
R34540 net3.n35 net3.n31 0.017
R34541 net3.n61 net3.n60 0.017
R34542 net3.n676 net3.n675 0.017
R34543 net3.n396 net3.n392 0.017
R34544 net3.n422 net3.n421 0.017
R34545 net3.n765 net3.n764 0.017
R34546 net3.n1039 net3.n1038 0.017
R34547 net3.n1063 net3.n1059 0.017
R34548 net3.n969 net3.n968 0.017
R34549 net3.n993 net3.n992 0.017
R34550 net3.n1126 net3.n1125 0.017
R34551 net3.n1400 net3.n1399 0.017
R34552 net3.n1424 net3.n1420 0.017
R34553 net3.n1330 net3.n1329 0.017
R34554 net3.n1354 net3.n1353 0.017
R34555 net3.n252 net3.n251 0.016
R34556 net3.n228 net3.n227 0.016
R34557 net3.n210 net3.n209 0.016
R34558 net3.n184 net3.n183 0.016
R34559 net3.n166 net3.n165 0.016
R34560 net3.n95 net3.n94 0.016
R34561 net3.n71 net3.n70 0.016
R34562 net3.n613 net3.n612 0.016
R34563 net3.n589 net3.n588 0.016
R34564 net3.n571 net3.n570 0.016
R34565 net3.n545 net3.n544 0.016
R34566 net3.n527 net3.n526 0.016
R34567 net3.n456 net3.n455 0.016
R34568 net3.n432 net3.n431 0.016
R34569 net3.n815 net3.n814 0.016
R34570 net3.n832 net3.n831 0.016
R34571 net3.n858 net3.n857 0.016
R34572 net3.n877 net3.n876 0.016
R34573 net3.n965 net3.n964 0.016
R34574 net3.n981 net3.n980 0.016
R34575 net3.n1008 net3.n1007 0.016
R34576 net3.n1176 net3.n1175 0.016
R34577 net3.n1193 net3.n1192 0.016
R34578 net3.n1219 net3.n1218 0.016
R34579 net3.n1238 net3.n1237 0.016
R34580 net3.n1326 net3.n1325 0.016
R34581 net3.n1342 net3.n1341 0.016
R34582 net3.n1369 net3.n1368 0.016
R34583 net3.n343 net3.n342 0.015
R34584 net3.n337 net3.n336 0.015
R34585 net3.n335 net3.n334 0.015
R34586 net3.n152 net3.n151 0.015
R34587 net3.n37 net3.n36 0.015
R34588 net3.n43 net3.n42 0.015
R34589 net3.n248 net3.n247 0.015
R34590 net3.n238 net3.n235 0.015
R34591 net3.n237 net3.n236 0.015
R34592 net3.n215 net3.n214 0.015
R34593 net3.n206 net3.n205 0.015
R34594 net3.n195 net3.n194 0.015
R34595 net3.n162 net3.n161 0.015
R34596 net3.n111 net3.n110 0.015
R34597 net3.n106 net3.n105 0.015
R34598 net3.n66 net3.n65 0.015
R34599 net3.n3 net3.n2 0.015
R34600 net3.n704 net3.n703 0.015
R34601 net3.n698 net3.n697 0.015
R34602 net3.n696 net3.n695 0.015
R34603 net3.n513 net3.n512 0.015
R34604 net3.n398 net3.n397 0.015
R34605 net3.n404 net3.n403 0.015
R34606 net3.n609 net3.n608 0.015
R34607 net3.n599 net3.n596 0.015
R34608 net3.n598 net3.n597 0.015
R34609 net3.n576 net3.n575 0.015
R34610 net3.n567 net3.n566 0.015
R34611 net3.n556 net3.n555 0.015
R34612 net3.n523 net3.n522 0.015
R34613 net3.n472 net3.n471 0.015
R34614 net3.n467 net3.n466 0.015
R34615 net3.n427 net3.n426 0.015
R34616 net3.n364 net3.n363 0.015
R34617 net3.n790 net3.n789 0.015
R34618 net3.n784 net3.n783 0.015
R34619 net3.n782 net3.n781 0.015
R34620 net3.n937 net3.n936 0.015
R34621 net3.n1065 net3.n1064 0.015
R34622 net3.n1071 net3.n1070 0.015
R34623 net3.n726 net3.n725 0.015
R34624 net3.n806 net3.n805 0.015
R34625 net3.n811 net3.n810 0.015
R34626 net3.n842 net3.n841 0.015
R34627 net3.n853 net3.n852 0.015
R34628 net3.n862 net3.n861 0.015
R34629 net3.n949 net3.n948 0.015
R34630 net3.n951 net3.n950 0.015
R34631 net3.n960 net3.n959 0.015
R34632 net3.n991 net3.n990 0.015
R34633 net3.n1002 net3.n1001 0.015
R34634 net3.n1151 net3.n1150 0.015
R34635 net3.n1145 net3.n1144 0.015
R34636 net3.n1143 net3.n1142 0.015
R34637 net3.n1298 net3.n1297 0.015
R34638 net3.n1426 net3.n1425 0.015
R34639 net3.n1432 net3.n1431 0.015
R34640 net3.n1087 net3.n1086 0.015
R34641 net3.n1167 net3.n1166 0.015
R34642 net3.n1172 net3.n1171 0.015
R34643 net3.n1203 net3.n1202 0.015
R34644 net3.n1214 net3.n1213 0.015
R34645 net3.n1223 net3.n1222 0.015
R34646 net3.n1310 net3.n1309 0.015
R34647 net3.n1312 net3.n1311 0.015
R34648 net3.n1321 net3.n1320 0.015
R34649 net3.n1352 net3.n1351 0.015
R34650 net3.n1363 net3.n1362 0.015
R34651 net3.n346 net3.n343 0.013
R34652 net3.n286 net3.n285 0.013
R34653 net3.n46 net3.n43 0.013
R34654 net3.n249 net3.n246 0.013
R34655 net3.n196 net3.n193 0.013
R34656 net3.n169 net3.n168 0.013
R34657 net3.n6 net3.n5 0.013
R34658 net3.n707 net3.n704 0.013
R34659 net3.n647 net3.n646 0.013
R34660 net3.n407 net3.n404 0.013
R34661 net3.n610 net3.n607 0.013
R34662 net3.n557 net3.n554 0.013
R34663 net3.n530 net3.n529 0.013
R34664 net3.n367 net3.n366 0.013
R34665 net3.n791 net3.n790 0.013
R34666 net3.n894 net3.n893 0.013
R34667 net3.n1074 net3.n1071 0.013
R34668 net3.n728 net3.n727 0.013
R34669 net3.n848 net3.n847 0.013
R34670 net3.n1005 net3.n1004 0.013
R34671 net3.n1152 net3.n1151 0.013
R34672 net3.n1255 net3.n1254 0.013
R34673 net3.n1435 net3.n1432 0.013
R34674 net3.n1089 net3.n1088 0.013
R34675 net3.n1209 net3.n1208 0.013
R34676 net3.n1366 net3.n1365 0.013
R34677 net3.n334 net3.n333 0.011
R34678 net3.n304 net3.n303 0.011
R34679 net3.n139 net3.n138 0.011
R34680 net3.n31 net3.n30 0.011
R34681 net3.n695 net3.n694 0.011
R34682 net3.n665 net3.n664 0.011
R34683 net3.n500 net3.n499 0.011
R34684 net3.n392 net3.n391 0.011
R34685 net3.n781 net3.n780 0.011
R34686 net3.n757 net3.n756 0.011
R34687 net3.n1025 net3.n1024 0.011
R34688 net3.n1059 net3.n1058 0.011
R34689 net3.n1142 net3.n1141 0.011
R34690 net3.n1118 net3.n1117 0.011
R34691 net3.n1386 net3.n1385 0.011
R34692 net3.n1420 net3.n1419 0.011
R34693 net3.n342 net3.n340 0.009
R34694 net3.n314 net3.n313 0.009
R34695 net3.n88 net3.n87 0.009
R34696 net3.n18 net3.n17 0.009
R34697 net3.n49 net3.n48 0.009
R34698 net3.n359 net3.n358 0.009
R34699 net3.n217 net3.n216 0.009
R34700 net3.n200 net3.n199 0.009
R34701 net3.n92 net3.n80 0.009
R34702 net3.n77 net3.n76 0.009
R34703 net3.n8 net3.n7 0.009
R34704 net3.n250 net3.n245 0.009
R34705 net3.n244 net3.n243 0.009
R34706 net3.n239 net3.n234 0.009
R34707 net3.n233 net3.n232 0.009
R34708 net3.n208 net3.n203 0.009
R34709 net3.n202 net3.n201 0.009
R34710 net3.n197 net3.n192 0.009
R34711 net3.n191 net3.n190 0.009
R34712 net3.n164 net3.n114 0.009
R34713 net3.n113 net3.n112 0.009
R34714 net3.n108 net3.n103 0.009
R34715 net3.n102 net3.n101 0.009
R34716 net3.n69 net3.n64 0.009
R34717 net3.n63 net3.n62 0.009
R34718 net3.n58 net3.n57 0.009
R34719 net3.n56 net3.n55 0.009
R34720 net3.n703 net3.n701 0.009
R34721 net3.n675 net3.n674 0.009
R34722 net3.n449 net3.n448 0.009
R34723 net3.n379 net3.n378 0.009
R34724 net3.n410 net3.n409 0.009
R34725 net3.n720 net3.n719 0.009
R34726 net3.n578 net3.n577 0.009
R34727 net3.n561 net3.n560 0.009
R34728 net3.n453 net3.n441 0.009
R34729 net3.n438 net3.n437 0.009
R34730 net3.n369 net3.n368 0.009
R34731 net3.n611 net3.n606 0.009
R34732 net3.n605 net3.n604 0.009
R34733 net3.n600 net3.n595 0.009
R34734 net3.n594 net3.n593 0.009
R34735 net3.n569 net3.n564 0.009
R34736 net3.n563 net3.n562 0.009
R34737 net3.n558 net3.n553 0.009
R34738 net3.n552 net3.n551 0.009
R34739 net3.n525 net3.n475 0.009
R34740 net3.n474 net3.n473 0.009
R34741 net3.n469 net3.n464 0.009
R34742 net3.n463 net3.n462 0.009
R34743 net3.n430 net3.n425 0.009
R34744 net3.n424 net3.n423 0.009
R34745 net3.n419 net3.n418 0.009
R34746 net3.n417 net3.n416 0.009
R34747 net3.n789 net3.n787 0.009
R34748 net3.n764 net3.n763 0.009
R34749 net3.n1038 net3.n1037 0.009
R34750 net3.n1046 net3.n1045 0.009
R34751 net3.n1077 net3.n1076 0.009
R34752 net3.n829 net3.n828 0.009
R34753 net3.n844 net3.n843 0.009
R34754 net3.n972 net3.n970 0.009
R34755 net3.n976 net3.n975 0.009
R34756 net3.n978 net3.n977 0.009
R34757 net3.n1010 net3.n1009 0.009
R34758 net3.n1082 net3.n1013 0.009
R34759 net3.n801 net3.n800 0.009
R34760 net3.n803 net3.n802 0.009
R34761 net3.n808 net3.n807 0.009
R34762 net3.n813 net3.n809 0.009
R34763 net3.n839 net3.n838 0.009
R34764 net3.n845 net3.n840 0.009
R34765 net3.n850 net3.n849 0.009
R34766 net3.n856 net3.n851 0.009
R34767 net3.n946 net3.n945 0.009
R34768 net3.n952 net3.n947 0.009
R34769 net3.n957 net3.n956 0.009
R34770 net3.n963 net3.n958 0.009
R34771 net3.n988 net3.n987 0.009
R34772 net3.n994 net3.n989 0.009
R34773 net3.n999 net3.n998 0.009
R34774 net3.n1006 net3.n1000 0.009
R34775 net3.n1150 net3.n1148 0.009
R34776 net3.n1125 net3.n1124 0.009
R34777 net3.n1399 net3.n1398 0.009
R34778 net3.n1407 net3.n1406 0.009
R34779 net3.n1438 net3.n1437 0.009
R34780 net3.n1190 net3.n1189 0.009
R34781 net3.n1205 net3.n1204 0.009
R34782 net3.n1333 net3.n1331 0.009
R34783 net3.n1337 net3.n1336 0.009
R34784 net3.n1339 net3.n1338 0.009
R34785 net3.n1371 net3.n1370 0.009
R34786 net3.n1443 net3.n1374 0.009
R34787 net3.n1162 net3.n1161 0.009
R34788 net3.n1164 net3.n1163 0.009
R34789 net3.n1169 net3.n1168 0.009
R34790 net3.n1174 net3.n1170 0.009
R34791 net3.n1200 net3.n1199 0.009
R34792 net3.n1206 net3.n1201 0.009
R34793 net3.n1211 net3.n1210 0.009
R34794 net3.n1217 net3.n1212 0.009
R34795 net3.n1307 net3.n1306 0.009
R34796 net3.n1313 net3.n1308 0.009
R34797 net3.n1318 net3.n1317 0.009
R34798 net3.n1324 net3.n1319 0.009
R34799 net3.n1349 net3.n1348 0.009
R34800 net3.n1355 net3.n1350 0.009
R34801 net3.n1360 net3.n1359 0.009
R34802 net3.n1367 net3.n1361 0.009
R34803 net3.n349 net3.n348 0.007
R34804 net3.n339 net3.n338 0.007
R34805 net3.n319 net3.n318 0.007
R34806 net3.n313 net3.n312 0.007
R34807 net3.n290 net3.n289 0.007
R34808 net3.n118 net3.n117 0.007
R34809 net3.n127 net3.n126 0.007
R34810 net3.n149 net3.n148 0.007
R34811 net3.n144 net3.n143 0.007
R34812 net3.n142 net3.n141 0.007
R34813 net3.n138 net3.n137 0.007
R34814 net3.n89 net3.n88 0.007
R34815 net3.n42 net3.n40 0.007
R34816 net3.n355 net3.n354 0.007
R34817 net3.n242 net3.n241 0.007
R34818 net3.n225 net3.n220 0.007
R34819 net3.n224 net3.n223 0.007
R34820 net3.n176 net3.n175 0.007
R34821 net3.n178 net3.n177 0.007
R34822 net3.n171 net3.n170 0.007
R34823 net3.n107 net3.n104 0.007
R34824 net3.n100 net3.n99 0.007
R34825 net3.n98 net3.n97 0.007
R34826 net3.n710 net3.n709 0.007
R34827 net3.n700 net3.n699 0.007
R34828 net3.n680 net3.n679 0.007
R34829 net3.n674 net3.n673 0.007
R34830 net3.n651 net3.n650 0.007
R34831 net3.n479 net3.n478 0.007
R34832 net3.n488 net3.n487 0.007
R34833 net3.n510 net3.n509 0.007
R34834 net3.n505 net3.n504 0.007
R34835 net3.n503 net3.n502 0.007
R34836 net3.n499 net3.n498 0.007
R34837 net3.n450 net3.n449 0.007
R34838 net3.n403 net3.n401 0.007
R34839 net3.n716 net3.n715 0.007
R34840 net3.n603 net3.n602 0.007
R34841 net3.n586 net3.n581 0.007
R34842 net3.n585 net3.n584 0.007
R34843 net3.n537 net3.n536 0.007
R34844 net3.n539 net3.n538 0.007
R34845 net3.n532 net3.n531 0.007
R34846 net3.n468 net3.n465 0.007
R34847 net3.n461 net3.n460 0.007
R34848 net3.n459 net3.n458 0.007
R34849 net3.n794 net3.n793 0.007
R34850 net3.n786 net3.n785 0.007
R34851 net3.n769 net3.n768 0.007
R34852 net3.n763 net3.n762 0.007
R34853 net3.n888 net3.n887 0.007
R34854 net3.n918 net3.n917 0.007
R34855 net3.n927 net3.n926 0.007
R34856 net3.n934 net3.n933 0.007
R34857 net3.n1018 net3.n1017 0.007
R34858 net3.n1022 net3.n1019 0.007
R34859 net3.n1030 net3.n1025 0.007
R34860 net3.n1037 net3.n1036 0.007
R34861 net3.n1070 net3.n1068 0.007
R34862 net3.n730 net3.n729 0.007
R34863 net3.n724 net3.n723 0.007
R34864 net3.n820 net3.n819 0.007
R34865 net3.n823 net3.n822 0.007
R34866 net3.n864 net3.n863 0.007
R34867 net3.n870 net3.n869 0.007
R34868 net3.n873 net3.n872 0.007
R34869 net3.n955 net3.n954 0.007
R34870 net3.n962 net3.n961 0.007
R34871 net3.n967 net3.n966 0.007
R34872 net3.n1155 net3.n1154 0.007
R34873 net3.n1147 net3.n1146 0.007
R34874 net3.n1130 net3.n1129 0.007
R34875 net3.n1124 net3.n1123 0.007
R34876 net3.n1249 net3.n1248 0.007
R34877 net3.n1279 net3.n1278 0.007
R34878 net3.n1288 net3.n1287 0.007
R34879 net3.n1295 net3.n1294 0.007
R34880 net3.n1379 net3.n1378 0.007
R34881 net3.n1383 net3.n1380 0.007
R34882 net3.n1391 net3.n1386 0.007
R34883 net3.n1398 net3.n1397 0.007
R34884 net3.n1431 net3.n1429 0.007
R34885 net3.n1091 net3.n1090 0.007
R34886 net3.n1085 net3.n1084 0.007
R34887 net3.n1181 net3.n1180 0.007
R34888 net3.n1184 net3.n1183 0.007
R34889 net3.n1225 net3.n1224 0.007
R34890 net3.n1231 net3.n1230 0.007
R34891 net3.n1234 net3.n1233 0.007
R34892 net3.n1316 net3.n1315 0.007
R34893 net3.n1323 net3.n1322 0.007
R34894 net3.n1328 net3.n1327 0.007
R34895 net3.n336 net3.n335 0.005
R34896 net3.n333 net3.n331 0.005
R34897 net3.n316 net3.n315 0.005
R34898 net3.n307 net3.n306 0.005
R34899 net3.n305 net3.n304 0.005
R34900 net3.n302 net3.n301 0.005
R34901 net3.n301 net3.n298 0.005
R34902 net3.n297 net3.n296 0.005
R34903 net3.n272 net3.n271 0.005
R34904 net3.n116 net3.n115 0.005
R34905 net3.n83 net3.n82 0.005
R34906 net3.n12 net3.n11 0.005
R34907 net3.n39 net3.n38 0.005
R34908 net3.n217 net3.n211 0.005
R34909 net3.n213 net3.n212 0.005
R34910 net3.n207 net3.n204 0.005
R34911 net3.n180 net3.n179 0.005
R34912 net3.n92 net3.n91 0.005
R34913 net3.n1 net3.n0 0.005
R34914 net3.n245 net3.n244 0.005
R34915 net3.n234 net3.n233 0.005
R34916 net3.n203 net3.n202 0.005
R34917 net3.n192 net3.n191 0.005
R34918 net3.n114 net3.n113 0.005
R34919 net3.n103 net3.n102 0.005
R34920 net3.n64 net3.n63 0.005
R34921 net3.n57 net3.n56 0.005
R34922 net3.n697 net3.n696 0.005
R34923 net3.n694 net3.n692 0.005
R34924 net3.n677 net3.n676 0.005
R34925 net3.n668 net3.n667 0.005
R34926 net3.n666 net3.n665 0.005
R34927 net3.n663 net3.n662 0.005
R34928 net3.n662 net3.n659 0.005
R34929 net3.n658 net3.n657 0.005
R34930 net3.n633 net3.n632 0.005
R34931 net3.n477 net3.n476 0.005
R34932 net3.n444 net3.n443 0.005
R34933 net3.n373 net3.n372 0.005
R34934 net3.n400 net3.n399 0.005
R34935 net3.n578 net3.n572 0.005
R34936 net3.n574 net3.n573 0.005
R34937 net3.n568 net3.n565 0.005
R34938 net3.n541 net3.n540 0.005
R34939 net3.n453 net3.n452 0.005
R34940 net3.n362 net3.n361 0.005
R34941 net3.n606 net3.n605 0.005
R34942 net3.n595 net3.n594 0.005
R34943 net3.n564 net3.n563 0.005
R34944 net3.n553 net3.n552 0.005
R34945 net3.n475 net3.n474 0.005
R34946 net3.n464 net3.n463 0.005
R34947 net3.n425 net3.n424 0.005
R34948 net3.n418 net3.n417 0.005
R34949 net3.n783 net3.n782 0.005
R34950 net3.n780 net3.n778 0.005
R34951 net3.n766 net3.n765 0.005
R34952 net3.n760 net3.n759 0.005
R34953 net3.n758 net3.n757 0.005
R34954 net3.n755 net3.n754 0.005
R34955 net3.n754 net3.n751 0.005
R34956 net3.n881 net3.n880 0.005
R34957 net3.n910 net3.n907 0.005
R34958 net3.n916 net3.n915 0.005
R34959 net3.n1032 net3.n1031 0.005
R34960 net3.n1040 net3.n1039 0.005
R34961 net3.n1067 net3.n1066 0.005
R34962 net3.n829 net3.n826 0.005
R34963 net3.n835 net3.n834 0.005
R34964 net3.n837 net3.n836 0.005
R34965 net3.n868 net3.n867 0.005
R34966 net3.n972 net3.n971 0.005
R34967 net3.n997 net3.n996 0.005
R34968 net3.n802 net3.n801 0.005
R34969 net3.n809 net3.n808 0.005
R34970 net3.n840 net3.n839 0.005
R34971 net3.n851 net3.n850 0.005
R34972 net3.n947 net3.n946 0.005
R34973 net3.n958 net3.n957 0.005
R34974 net3.n989 net3.n988 0.005
R34975 net3.n1000 net3.n999 0.005
R34976 net3.n1144 net3.n1143 0.005
R34977 net3.n1141 net3.n1139 0.005
R34978 net3.n1127 net3.n1126 0.005
R34979 net3.n1121 net3.n1120 0.005
R34980 net3.n1119 net3.n1118 0.005
R34981 net3.n1116 net3.n1115 0.005
R34982 net3.n1115 net3.n1112 0.005
R34983 net3.n1242 net3.n1241 0.005
R34984 net3.n1271 net3.n1268 0.005
R34985 net3.n1277 net3.n1276 0.005
R34986 net3.n1393 net3.n1392 0.005
R34987 net3.n1401 net3.n1400 0.005
R34988 net3.n1428 net3.n1427 0.005
R34989 net3.n1190 net3.n1187 0.005
R34990 net3.n1196 net3.n1195 0.005
R34991 net3.n1198 net3.n1197 0.005
R34992 net3.n1229 net3.n1228 0.005
R34993 net3.n1333 net3.n1332 0.005
R34994 net3.n1358 net3.n1357 0.005
R34995 net3.n1163 net3.n1162 0.005
R34996 net3.n1170 net3.n1169 0.005
R34997 net3.n1201 net3.n1200 0.005
R34998 net3.n1212 net3.n1211 0.005
R34999 net3.n1308 net3.n1307 0.005
R35000 net3.n1319 net3.n1318 0.005
R35001 net3.n1350 net3.n1349 0.005
R35002 net3.n1361 net3.n1360 0.005
R35003 net3.n347 net3.n346 0.003
R35004 net3.n160 net3.n129 0.003
R35005 net3.n157 net3.n155 0.003
R35006 net3.n141 net3.n140 0.003
R35007 net3.n16 net3.n12 0.003
R35008 net3.n30 net3.n28 0.003
R35009 net3.n36 net3.n35 0.003
R35010 net3.n47 net3.n46 0.003
R35011 net3.n360 net3.n252 0.003
R35012 net3.n227 net3.n226 0.003
R35013 net3.n218 net3.n210 0.003
R35014 net3.n183 net3.n182 0.003
R35015 net3.n173 net3.n166 0.003
R35016 net3.n94 net3.n93 0.003
R35017 net3.n78 net3.n71 0.003
R35018 net3.n708 net3.n707 0.003
R35019 net3.n521 net3.n490 0.003
R35020 net3.n518 net3.n516 0.003
R35021 net3.n502 net3.n501 0.003
R35022 net3.n377 net3.n373 0.003
R35023 net3.n391 net3.n389 0.003
R35024 net3.n397 net3.n396 0.003
R35025 net3.n408 net3.n407 0.003
R35026 net3.n721 net3.n613 0.003
R35027 net3.n588 net3.n587 0.003
R35028 net3.n579 net3.n571 0.003
R35029 net3.n544 net3.n543 0.003
R35030 net3.n534 net3.n527 0.003
R35031 net3.n455 net3.n454 0.003
R35032 net3.n439 net3.n432 0.003
R35033 net3.n792 net3.n791 0.003
R35034 net3.n943 net3.n929 0.003
R35035 net3.n942 net3.n940 0.003
R35036 net3.n1023 net3.n1022 0.003
R35037 net3.n1044 net3.n1040 0.003
R35038 net3.n1058 net3.n1056 0.003
R35039 net3.n1064 net3.n1063 0.003
R35040 net3.n1075 net3.n1074 0.003
R35041 net3.n821 net3.n815 0.003
R35042 net3.n831 net3.n830 0.003
R35043 net3.n866 net3.n858 0.003
R35044 net3.n876 net3.n875 0.003
R35045 net3.n973 net3.n965 0.003
R35046 net3.n980 net3.n979 0.003
R35047 net3.n1083 net3.n1008 0.003
R35048 net3.n1153 net3.n1152 0.003
R35049 net3.n1304 net3.n1290 0.003
R35050 net3.n1303 net3.n1301 0.003
R35051 net3.n1384 net3.n1383 0.003
R35052 net3.n1405 net3.n1401 0.003
R35053 net3.n1419 net3.n1417 0.003
R35054 net3.n1425 net3.n1424 0.003
R35055 net3.n1436 net3.n1435 0.003
R35056 net3.n1182 net3.n1176 0.003
R35057 net3.n1192 net3.n1191 0.003
R35058 net3.n1227 net3.n1219 0.003
R35059 net3.n1237 net3.n1236 0.003
R35060 net3.n1334 net3.n1326 0.003
R35061 net3.n1341 net3.n1340 0.003
R35062 net3.n1444 net3.n1369 0.003
R35063 net3.n328 net3.n327 0.001
R35064 net3.n323 net3.n321 0.001
R35065 net3.n317 net3.n316 0.001
R35066 net3.n312 net3.n311 0.001
R35067 net3.n295 net3.n292 0.001
R35068 net3.n289 net3.n288 0.001
R35069 net3.n284 net3.n281 0.001
R35070 net3.n279 net3.n278 0.001
R35071 net3.n278 net3.n275 0.001
R35072 net3.n274 net3.n273 0.001
R35073 net3.n268 net3.n267 0.001
R35074 net3.n123 net3.n119 0.001
R35075 net3.n24 net3.n21 0.001
R35076 net3.n26 net3.n25 0.001
R35077 net3.n220 net3.n219 0.001
R35078 net3.n222 net3.n221 0.001
R35079 net3.n189 net3.n188 0.001
R35080 net3.n187 net3.n186 0.001
R35081 net3.n181 net3.n176 0.001
R35082 net3.n172 net3.n171 0.001
R35083 net3.n74 net3.n73 0.001
R35084 net3.n68 net3.n67 0.001
R35085 net3.n4 net3.n3 0.001
R35086 net3.n689 net3.n688 0.001
R35087 net3.n684 net3.n682 0.001
R35088 net3.n678 net3.n677 0.001
R35089 net3.n673 net3.n672 0.001
R35090 net3.n656 net3.n653 0.001
R35091 net3.n650 net3.n649 0.001
R35092 net3.n645 net3.n642 0.001
R35093 net3.n640 net3.n639 0.001
R35094 net3.n639 net3.n636 0.001
R35095 net3.n635 net3.n634 0.001
R35096 net3.n629 net3.n628 0.001
R35097 net3.n484 net3.n480 0.001
R35098 net3.n385 net3.n382 0.001
R35099 net3.n387 net3.n386 0.001
R35100 net3.n581 net3.n580 0.001
R35101 net3.n583 net3.n582 0.001
R35102 net3.n550 net3.n549 0.001
R35103 net3.n548 net3.n547 0.001
R35104 net3.n542 net3.n537 0.001
R35105 net3.n533 net3.n532 0.001
R35106 net3.n435 net3.n434 0.001
R35107 net3.n429 net3.n428 0.001
R35108 net3.n365 net3.n364 0.001
R35109 net3.n775 net3.n774 0.001
R35110 net3.n773 net3.n771 0.001
R35111 net3.n767 net3.n766 0.001
R35112 net3.n762 net3.n761 0.001
R35113 net3.n886 net3.n884 0.001
R35114 net3.n891 net3.n888 0.001
R35115 net3.n899 net3.n897 0.001
R35116 net3.n903 net3.n900 0.001
R35117 net3.n904 net3.n903 0.001
R35118 net3.n906 net3.n905 0.001
R35119 net3.n914 net3.n913 0.001
R35120 net3.n923 net3.n919 0.001
R35121 net3.n1052 net3.n1049 0.001
R35122 net3.n1054 net3.n1053 0.001
R35123 net3.n819 net3.n818 0.001
R35124 net3.n825 net3.n824 0.001
R35125 net3.n855 net3.n854 0.001
R35126 net3.n860 net3.n859 0.001
R35127 net3.n865 net3.n864 0.001
R35128 net3.n874 net3.n873 0.001
R35129 net3.n984 net3.n983 0.001
R35130 net3.n986 net3.n985 0.001
R35131 net3.n1003 net3.n1002 0.001
R35132 net3.n1136 net3.n1135 0.001
R35133 net3.n1134 net3.n1132 0.001
R35134 net3.n1128 net3.n1127 0.001
R35135 net3.n1123 net3.n1122 0.001
R35136 net3.n1247 net3.n1245 0.001
R35137 net3.n1252 net3.n1249 0.001
R35138 net3.n1260 net3.n1258 0.001
R35139 net3.n1264 net3.n1261 0.001
R35140 net3.n1265 net3.n1264 0.001
R35141 net3.n1267 net3.n1266 0.001
R35142 net3.n1275 net3.n1274 0.001
R35143 net3.n1284 net3.n1280 0.001
R35144 net3.n1413 net3.n1410 0.001
R35145 net3.n1415 net3.n1414 0.001
R35146 net3.n1180 net3.n1179 0.001
R35147 net3.n1186 net3.n1185 0.001
R35148 net3.n1216 net3.n1215 0.001
R35149 net3.n1221 net3.n1220 0.001
R35150 net3.n1226 net3.n1225 0.001
R35151 net3.n1235 net3.n1234 0.001
R35152 net3.n1345 net3.n1344 0.001
R35153 net3.n1347 net3.n1346 0.001
R35154 net3.n1364 net3.n1363 0.001
R35155 net6_ota.n122 net6_ota.n121 13.176
R35156 net6_ota.n0 net6_ota.t2 12.018
R35157 net6_ota.n0 net6_ota.t0 11.988
R35158 net6_ota.n343 net6_ota.n342 9.3
R35159 net6_ota.n156 net6_ota.n155 9.3
R35160 net6_ota.n282 net6_ota.n281 9.3
R35161 net6_ota.n285 net6_ota.n284 9.3
R35162 net6_ota.n293 net6_ota.n292 9.3
R35163 net6_ota.n332 net6_ota.n331 9.3
R35164 net6_ota.n334 net6_ota.n333 9.3
R35165 net6_ota.n322 net6_ota.n321 9.3
R35166 net6_ota.n324 net6_ota.n323 9.3
R35167 net6_ota.n296 net6_ota.n295 9.3
R35168 net6_ota.n272 net6_ota.n271 9.3
R35169 net6_ota.n127 net6_ota.n126 9.3
R35170 net6_ota.n158 net6_ota.n157 9.3
R35171 net6_ota.n43 net6_ota.n42 9.3
R35172 net6_ota.n31 net6_ota.n30 9.3
R35173 net6_ota.n29 net6_ota.n28 9.3
R35174 net6_ota.n53 net6_ota.n52 8.454
R35175 net6_ota.n354 net6_ota.n353 8.454
R35176 net6_ota net6_ota.n361 6.851
R35177 net6_ota.n284 net6_ota.n283 5.458
R35178 net6_ota.n155 net6_ota.n154 5.081
R35179 net6_ota.n21 net6_ota.n20 4.65
R35180 net6_ota.n148 net6_ota.n147 4.65
R35181 net6_ota.n36 net6_ota.n35 4.5
R35182 net6_ota.n312 net6_ota.n311 4.5
R35183 net6_ota.n306 net6_ota.n263 4.5
R35184 net6_ota.n318 net6_ota.n259 4.5
R35185 net6_ota.n328 net6_ota.n327 4.5
R35186 net6_ota.n336 net6_ota.n256 4.5
R35187 net6_ota.n302 net6_ota.n301 4.5
R35188 net6_ota.n289 net6_ota.n265 4.5
R35189 net6_ota.n279 net6_ota.n278 4.5
R35190 net6_ota.n269 net6_ota.n267 4.5
R35191 net6_ota.n124 net6_ota.n123 4.5
R35192 net6_ota.n161 net6_ota.n160 4.5
R35193 net6_ota.n142 net6_ota.n133 4.5
R35194 net6_ota.n90 net6_ota.n87 4.5
R35195 net6_ota.n138 net6_ota.n137 4.5
R35196 net6_ota.n17 net6_ota.n16 4.5
R35197 net6_ota.n47 net6_ota.n46 4.5
R35198 net6_ota.n347 net6_ota.n346 4.5
R35199 net6_ota.n259 net6_ota.n257 4.325
R35200 net6_ota.n352 net6_ota.t1 4.289
R35201 net6_ota.n263 net6_ota.n260 3.95
R35202 net6_ota.n16 net6_ota.n15 3.948
R35203 net6_ota.n137 net6_ota.n136 3.573
R35204 net6_ota net6_ota.n0 3.353
R35205 net6_ota.n150 net6_ota.n131 3.033
R35206 net6_ota.n25 net6_ota.n24 3.033
R35207 net6_ota.n262 net6_ota.n261 2.258
R35208 net6_ota.n135 net6_ota.n134 2.258
R35209 net6_ota.n310 net6_ota.n309 1.882
R35210 net6_ota.n311 net6_ota.n310 1.882
R35211 net6_ota.n86 net6_ota.n85 1.882
R35212 net6_ota.n353 net6_ota.n352 1.844
R35213 net6_ota.n137 net6_ota.n135 1.505
R35214 net6_ota.n87 net6_ota.n86 1.505
R35215 net6_ota.n361 net6_ota.n360 1.137
R35216 net6_ota.n113 net6_ota.n112 1.137
R35217 net6_ota.n191 net6_ota.n190 1.137
R35218 net6_ota.n198 net6_ota.n197 1.137
R35219 net6_ota.n202 net6_ota.n201 1.137
R35220 net6_ota.n209 net6_ota.n208 1.137
R35221 net6_ota.n227 net6_ota.n226 1.137
R35222 net6_ota.n244 net6_ota.n243 1.137
R35223 net6_ota.n240 net6_ota.n239 1.137
R35224 net6_ota.n233 net6_ota.n232 1.137
R35225 net6_ota.n219 net6_ota.n218 1.137
R35226 net6_ota.n183 net6_ota.n182 1.137
R35227 net6_ota.n174 net6_ota.n173 1.137
R35228 net6_ota.n165 net6_ota.n164 1.137
R35229 net6_ota.n102 net6_ota.n101 1.137
R35230 net6_ota.n109 net6_ota.n108 1.137
R35231 net6_ota.n94 net6_ota.n93 1.137
R35232 net6_ota.n79 net6_ota.n78 1.137
R35233 net6_ota.n63 net6_ota.n62 1.137
R35234 net6_ota.n70 net6_ota.n69 1.137
R35235 net6_ota.n251 net6_ota.n250 1.137
R35236 net6_ota.n256 net6_ota.n255 1.129
R35237 net6_ota.n263 net6_ota.n262 1.129
R35238 net6_ota.n301 net6_ota.n300 1.129
R35239 net6_ota.n91 net6_ota.n90 1.125
R35240 net6_ota.n164 net6_ota.n161 1.042
R35241 net6_ota.n55 net6_ota.n54 0.869
R35242 net6_ota.n346 net6_ota.n345 0.752
R35243 net6_ota.n160 net6_ota.n159 0.752
R35244 net6_ota.n133 net6_ota.n132 0.752
R35245 net6_ota.n16 net6_ota.n14 0.752
R35246 net6_ota.n35 net6_ota.n34 0.752
R35247 net6_ota.n46 net6_ota.n45 0.752
R35248 net6_ota.n54 net6_ota.n53 0.728
R35249 net6_ota.n360 net6_ota.n354 0.725
R35250 net6_ota.n327 net6_ota.n326 0.376
R35251 net6_ota.n259 net6_ota.n258 0.376
R35252 net6_ota.n265 net6_ota.n264 0.376
R35253 net6_ota.n278 net6_ota.n277 0.376
R35254 net6_ota.n267 net6_ota.n266 0.376
R35255 net6_ota.n123 net6_ota.n122 0.376
R35256 net6_ota.n126 net6_ota.n125 0.189
R35257 net6_ota.n271 net6_ota.n270 0.188
R35258 net6_ota.n147 net6_ota.n146 0.166
R35259 net6_ota.n295 net6_ota.n294 0.166
R35260 net6_ota.n24 net6_ota.n23 0.133
R35261 net6_ota.n326 net6_ota.n325 0.132
R35262 net6_ota.n34 net6_ota.n33 0.121
R35263 net6_ota.n255 net6_ota.n254 0.121
R35264 net6_ota.n232 net6_ota.n231 0.049
R35265 net6_ota.n227 net6_ota.n219 0.049
R35266 net6_ota.n183 net6_ota.n174 0.049
R35267 net6_ota.n94 net6_ota.n79 0.049
R35268 net6_ota.n351 net6_ota.n350 0.047
R35269 net6_ota.n332 net6_ota.n330 0.047
R35270 net6_ota.n330 net6_ota.n329 0.047
R35271 net6_ota.n322 net6_ota.n320 0.047
R35272 net6_ota.n274 net6_ota.n273 0.047
R35273 net6_ota.n129 net6_ota.n128 0.047
R35274 net6_ota.n21 net6_ota.n19 0.047
R35275 net6_ota.n26 net6_ota.n25 0.047
R35276 net6_ota.n29 net6_ota.n27 0.047
R35277 net6_ota.n51 net6_ota.n50 0.047
R35278 net6_ota.n189 net6_ota.n188 0.047
R35279 net6_ota.n276 net6_ota.n275 0.045
R35280 net6_ota.n130 net6_ota.n129 0.045
R35281 net6_ota.n299 net6_ota.n298 0.043
R35282 net6_ota.n90 net6_ota.n84 0.043
R35283 net6_ota.n182 net6_ota.n181 0.043
R35284 net6_ota.n92 net6_ota.n91 0.043
R35285 net6_ota.n77 net6_ota.n76 0.043
R35286 net6_ota.n354 net6_ota.n351 0.043
R35287 net6_ota.n319 net6_ota.n318 0.041
R35288 net6_ota.n312 net6_ota.n308 0.041
R35289 net6_ota.n120 net6_ota.n119 0.041
R35290 net6_ota.n144 net6_ota.n143 0.041
R35291 net6_ota.n41 net6_ota.n40 0.041
R35292 net6_ota.n226 net6_ota.n225 0.041
R35293 net6_ota.n100 net6_ota.n99 0.041
R35294 net6_ota.n53 net6_ota.n51 0.041
R35295 net6_ota.n341 net6_ota.n340 0.039
R35296 net6_ota.n297 net6_ota.n296 0.039
R35297 net6_ota.n148 net6_ota.n145 0.039
R35298 net6_ota.n18 net6_ota.n17 0.039
R35299 net6_ota.n78 net6_ota.n73 0.039
R35300 net6_ota.n307 net6_ota.n306 0.037
R35301 net6_ota.n8 net6_ota.n7 0.035
R35302 net6_ota.n286 net6_ota.n285 0.034
R35303 net6_ota.n118 net6_ota.n117 0.034
R35304 net6_ota.n231 net6_ota.n230 0.034
R35305 net6_ota.n224 net6_ota.n223 0.034
R35306 net6_ota.n180 net6_ota.n179 0.034
R35307 net6_ota.n169 net6_ota.n168 0.034
R35308 net6_ota.n91 net6_ota.n82 0.034
R35309 net6_ota.n76 net6_ota.n75 0.034
R35310 net6_ota.n349 net6_ota.n348 0.032
R35311 net6_ota.n156 net6_ota.n153 0.032
R35312 net6_ota.n49 net6_ota.n48 0.032
R35313 net6_ota.n187 net6_ota.n186 0.032
R35314 net6_ota.n252 net6_ota.n251 0.031
R35315 net6_ota.n233 net6_ota.n229 0.031
R35316 net6_ota.n210 net6_ota.n209 0.031
R35317 net6_ota.n191 net6_ota.n185 0.031
R35318 net6_ota.n166 net6_ota.n165 0.031
R35319 net6_ota.n102 net6_ota.n96 0.031
R35320 net6_ota.n71 net6_ota.n70 0.031
R35321 net6_ota.n56 net6_ota.n55 0.031
R35322 net6_ota.n328 net6_ota.n324 0.03
R35323 net6_ota.n272 net6_ota.n269 0.03
R35324 net6_ota.n127 net6_ota.n124 0.03
R35325 net6_ota.n22 net6_ota.n21 0.03
R35326 net6_ota.n39 net6_ota.n38 0.03
R35327 net6_ota.n171 net6_ota.n170 0.03
R35328 net6_ota.n339 net6_ota.n338 0.028
R35329 net6_ota.n282 net6_ota.n280 0.028
R35330 net6_ota.n161 net6_ota.n158 0.028
R35331 net6_ota.n151 net6_ota.n150 0.028
R35332 net6_ota.n242 net6_ota.n241 0.028
R35333 net6_ota.n217 net6_ota.n216 0.028
R35334 net6_ota.n215 net6_ota.n214 0.028
R35335 net6_ota.n176 net6_ota.n175 0.028
R35336 net6_ota.n54 net6_ota.n11 0.027
R35337 net6_ota.n244 net6_ota.n240 0.027
R35338 net6_ota.n202 net6_ota.n198 0.027
R35339 net6_ota.n113 net6_ota.n109 0.027
R35340 net6_ota.n63 net6_ota.n59 0.027
R35341 net6_ota.n289 net6_ota.n288 0.026
R35342 net6_ota.n357 net6_ota.n356 0.026
R35343 net6_ota.n200 net6_ota.n199 0.026
R35344 net6_ota.n98 net6_ota.n97 0.026
R35345 net6_ota.n81 net6_ota.n80 0.026
R35346 net6_ota.n149 net6_ota.n148 0.024
R35347 net6_ota.n250 net6_ota.n249 0.024
R35348 net6_ota.n239 net6_ota.n238 0.024
R35349 net6_ota.n208 net6_ota.n207 0.024
R35350 net6_ota.n197 net6_ota.n196 0.024
R35351 net6_ota.n164 net6_ota.n163 0.024
R35352 net6_ota.n108 net6_ota.n107 0.024
R35353 net6_ota.n3 net6_ota.n2 0.024
R35354 net6_ota.n10 net6_ota.n9 0.024
R35355 net6_ota.n293 net6_ota.n291 0.022
R35356 net6_ota.n288 net6_ota.n287 0.022
R35357 net6_ota.n359 net6_ota.n358 0.022
R35358 net6_ota.n68 net6_ota.n67 0.022
R35359 net6_ota.n6 net6_ota.n5 0.022
R35360 net6_ota.n11 net6_ota.n10 0.022
R35361 net6_ota.n304 net6_ota.n303 0.02
R35362 net6_ota.n152 net6_ota.n151 0.02
R35363 net6_ota.n141 net6_ota.n140 0.02
R35364 net6_ota.n358 net6_ota.n357 0.02
R35365 net6_ota.n111 net6_ota.n110 0.02
R35366 net6_ota.n61 net6_ota.n60 0.018
R35367 net6_ota.n316 net6_ota.n315 0.017
R35368 net6_ota.n36 net6_ota.n32 0.017
R35369 net6_ota.n62 net6_ota.n61 0.017
R35370 net6_ota.n253 net6_ota.n252 0.016
R35371 net6_ota.n229 net6_ota.n228 0.016
R35372 net6_ota.n211 net6_ota.n210 0.016
R35373 net6_ota.n185 net6_ota.n184 0.016
R35374 net6_ota.n167 net6_ota.n166 0.016
R35375 net6_ota.n96 net6_ota.n95 0.016
R35376 net6_ota.n72 net6_ota.n71 0.016
R35377 net6_ota.n344 net6_ota.n343 0.015
R35378 net6_ota.n338 net6_ota.n337 0.015
R35379 net6_ota.n336 net6_ota.n335 0.015
R35380 net6_ota.n153 net6_ota.n152 0.015
R35381 net6_ota.n38 net6_ota.n37 0.015
R35382 net6_ota.n44 net6_ota.n43 0.015
R35383 net6_ota.n249 net6_ota.n248 0.015
R35384 net6_ota.n239 net6_ota.n236 0.015
R35385 net6_ota.n238 net6_ota.n237 0.015
R35386 net6_ota.n216 net6_ota.n215 0.015
R35387 net6_ota.n207 net6_ota.n206 0.015
R35388 net6_ota.n196 net6_ota.n195 0.015
R35389 net6_ota.n163 net6_ota.n162 0.015
R35390 net6_ota.n112 net6_ota.n111 0.015
R35391 net6_ota.n107 net6_ota.n106 0.015
R35392 net6_ota.n67 net6_ota.n66 0.015
R35393 net6_ota.n4 net6_ota.n3 0.015
R35394 net6_ota.n347 net6_ota.n344 0.013
R35395 net6_ota.n287 net6_ota.n286 0.013
R35396 net6_ota.n47 net6_ota.n44 0.013
R35397 net6_ota.n250 net6_ota.n247 0.013
R35398 net6_ota.n197 net6_ota.n194 0.013
R35399 net6_ota.n170 net6_ota.n169 0.013
R35400 net6_ota.n7 net6_ota.n6 0.013
R35401 net6_ota.n335 net6_ota.n334 0.011
R35402 net6_ota.n305 net6_ota.n304 0.011
R35403 net6_ota.n140 net6_ota.n139 0.011
R35404 net6_ota.n32 net6_ota.n31 0.011
R35405 net6_ota.n343 net6_ota.n341 0.009
R35406 net6_ota.n315 net6_ota.n314 0.009
R35407 net6_ota.n89 net6_ota.n88 0.009
R35408 net6_ota.n19 net6_ota.n18 0.009
R35409 net6_ota.n50 net6_ota.n49 0.009
R35410 net6_ota.n360 net6_ota.n359 0.009
R35411 net6_ota.n218 net6_ota.n217 0.009
R35412 net6_ota.n201 net6_ota.n200 0.009
R35413 net6_ota.n93 net6_ota.n81 0.009
R35414 net6_ota.n78 net6_ota.n77 0.009
R35415 net6_ota.n9 net6_ota.n8 0.009
R35416 net6_ota.n251 net6_ota.n246 0.009
R35417 net6_ota.n245 net6_ota.n244 0.009
R35418 net6_ota.n240 net6_ota.n235 0.009
R35419 net6_ota.n234 net6_ota.n233 0.009
R35420 net6_ota.n209 net6_ota.n204 0.009
R35421 net6_ota.n203 net6_ota.n202 0.009
R35422 net6_ota.n198 net6_ota.n193 0.009
R35423 net6_ota.n192 net6_ota.n191 0.009
R35424 net6_ota.n165 net6_ota.n115 0.009
R35425 net6_ota.n114 net6_ota.n113 0.009
R35426 net6_ota.n109 net6_ota.n104 0.009
R35427 net6_ota.n103 net6_ota.n102 0.009
R35428 net6_ota.n70 net6_ota.n65 0.009
R35429 net6_ota.n64 net6_ota.n63 0.009
R35430 net6_ota.n59 net6_ota.n58 0.009
R35431 net6_ota.n57 net6_ota.n56 0.009
R35432 net6_ota.n350 net6_ota.n349 0.007
R35433 net6_ota.n340 net6_ota.n339 0.007
R35434 net6_ota.n320 net6_ota.n319 0.007
R35435 net6_ota.n314 net6_ota.n313 0.007
R35436 net6_ota.n291 net6_ota.n290 0.007
R35437 net6_ota.n119 net6_ota.n118 0.007
R35438 net6_ota.n128 net6_ota.n127 0.007
R35439 net6_ota.n150 net6_ota.n149 0.007
R35440 net6_ota.n145 net6_ota.n144 0.007
R35441 net6_ota.n143 net6_ota.n142 0.007
R35442 net6_ota.n139 net6_ota.n138 0.007
R35443 net6_ota.n90 net6_ota.n89 0.007
R35444 net6_ota.n43 net6_ota.n41 0.007
R35445 net6_ota.n356 net6_ota.n355 0.007
R35446 net6_ota.n243 net6_ota.n242 0.007
R35447 net6_ota.n226 net6_ota.n221 0.007
R35448 net6_ota.n225 net6_ota.n224 0.007
R35449 net6_ota.n177 net6_ota.n176 0.007
R35450 net6_ota.n179 net6_ota.n178 0.007
R35451 net6_ota.n172 net6_ota.n171 0.007
R35452 net6_ota.n108 net6_ota.n105 0.007
R35453 net6_ota.n101 net6_ota.n100 0.007
R35454 net6_ota.n99 net6_ota.n98 0.007
R35455 net6_ota.n337 net6_ota.n336 0.005
R35456 net6_ota.n334 net6_ota.n332 0.005
R35457 net6_ota.n317 net6_ota.n316 0.005
R35458 net6_ota.n308 net6_ota.n307 0.005
R35459 net6_ota.n306 net6_ota.n305 0.005
R35460 net6_ota.n303 net6_ota.n302 0.005
R35461 net6_ota.n302 net6_ota.n299 0.005
R35462 net6_ota.n298 net6_ota.n297 0.005
R35463 net6_ota.n273 net6_ota.n272 0.005
R35464 net6_ota.n117 net6_ota.n116 0.005
R35465 net6_ota.n84 net6_ota.n83 0.005
R35466 net6_ota.n13 net6_ota.n12 0.005
R35467 net6_ota.n40 net6_ota.n39 0.005
R35468 net6_ota.n218 net6_ota.n212 0.005
R35469 net6_ota.n214 net6_ota.n213 0.005
R35470 net6_ota.n208 net6_ota.n205 0.005
R35471 net6_ota.n181 net6_ota.n180 0.005
R35472 net6_ota.n93 net6_ota.n92 0.005
R35473 net6_ota.n2 net6_ota.n1 0.005
R35474 net6_ota.n246 net6_ota.n245 0.005
R35475 net6_ota.n235 net6_ota.n234 0.005
R35476 net6_ota.n204 net6_ota.n203 0.005
R35477 net6_ota.n193 net6_ota.n192 0.005
R35478 net6_ota.n115 net6_ota.n114 0.005
R35479 net6_ota.n104 net6_ota.n103 0.005
R35480 net6_ota.n65 net6_ota.n64 0.005
R35481 net6_ota.n58 net6_ota.n57 0.005
R35482 net6_ota.n348 net6_ota.n347 0.003
R35483 net6_ota.n161 net6_ota.n130 0.003
R35484 net6_ota.n158 net6_ota.n156 0.003
R35485 net6_ota.n142 net6_ota.n141 0.003
R35486 net6_ota.n17 net6_ota.n13 0.003
R35487 net6_ota.n31 net6_ota.n29 0.003
R35488 net6_ota.n37 net6_ota.n36 0.003
R35489 net6_ota.n48 net6_ota.n47 0.003
R35490 net6_ota.n361 net6_ota.n253 0.003
R35491 net6_ota.n228 net6_ota.n227 0.003
R35492 net6_ota.n219 net6_ota.n211 0.003
R35493 net6_ota.n184 net6_ota.n183 0.003
R35494 net6_ota.n174 net6_ota.n167 0.003
R35495 net6_ota.n95 net6_ota.n94 0.003
R35496 net6_ota.n79 net6_ota.n72 0.003
R35497 net6_ota.n329 net6_ota.n328 0.001
R35498 net6_ota.n324 net6_ota.n322 0.001
R35499 net6_ota.n318 net6_ota.n317 0.001
R35500 net6_ota.n313 net6_ota.n312 0.001
R35501 net6_ota.n296 net6_ota.n293 0.001
R35502 net6_ota.n290 net6_ota.n289 0.001
R35503 net6_ota.n285 net6_ota.n282 0.001
R35504 net6_ota.n280 net6_ota.n279 0.001
R35505 net6_ota.n279 net6_ota.n276 0.001
R35506 net6_ota.n275 net6_ota.n274 0.001
R35507 net6_ota.n269 net6_ota.n268 0.001
R35508 net6_ota.n124 net6_ota.n120 0.001
R35509 net6_ota.n25 net6_ota.n22 0.001
R35510 net6_ota.n27 net6_ota.n26 0.001
R35511 net6_ota.n221 net6_ota.n220 0.001
R35512 net6_ota.n223 net6_ota.n222 0.001
R35513 net6_ota.n190 net6_ota.n189 0.001
R35514 net6_ota.n188 net6_ota.n187 0.001
R35515 net6_ota.n182 net6_ota.n177 0.001
R35516 net6_ota.n173 net6_ota.n172 0.001
R35517 net6_ota.n75 net6_ota.n74 0.001
R35518 net6_ota.n69 net6_ota.n68 0.001
R35519 net6_ota.n5 net6_ota.n4 0.001
R35520 net2.n118 net2.t1 124.695
R35521 net2.n15 net2.n14 92.5
R35522 net2.n78 net2.n77 92.5
R35523 net2.n117 net2.n116 92.5
R35524 net2.n14 net2.t0 70.344
R35525 net2.n28 net2.n27 31.034
R35526 net2.n95 net2.n94 31.034
R35527 net2.n127 net2.n126 31.034
R35528 net2.n118 net2.n117 15.431
R35529 net2 net2.n135 11.103
R35530 net2.n38 net2.n37 9.3
R35531 net2.n104 net2.n103 9.3
R35532 net2.n96 net2.n95 9.3
R35533 net2.n29 net2.n28 9.3
R35534 net2.n133 net2.n132 9.3
R35535 net2.n122 net2.n121 9.3
R35536 net2.n120 net2.n119 9.3
R35537 net2.n129 net2.n128 9.3
R35538 net2.n128 net2.n127 9.3
R35539 net2.n131 net2.n130 9.3
R35540 net2.n135 net2.n134 9.3
R35541 net2.n16 net2.n15 8.282
R35542 net2.n79 net2.n78 8.282
R35543 net2.n29 net2.n25 5.647
R35544 net2.n96 net2.n92 5.647
R35545 net2.n128 net2.n124 5.647
R35546 net2.n76 net2.n75 4.65
R35547 net2.n80 net2.n79 4.5
R35548 net2.n87 net2.n86 4.5
R35549 net2.n21 net2.n16 4.5
R35550 net2.n98 net2.n97 4.5
R35551 net2.n74 net2.n73 4.5
R35552 net2.n32 net2.n31 4.5
R35553 net2.n110 net2.n108 4.5
R35554 net2.n43 net2.n42 4.5
R35555 net2.n27 net2.n26 4.137
R35556 net2.n94 net2.n93 4.137
R35557 net2.n126 net2.n125 4.137
R35558 net2.n42 net2.n40 3.764
R35559 net2.n97 net2.n90 3.764
R35560 net2 net2.n115 3.424
R35561 net2.n31 net2.n30 3.388
R35562 net2.n108 net2.n107 3.388
R35563 net2.n31 net2.n29 3.011
R35564 net2.n16 net2.n13 3.011
R35565 net2.n108 net2.n106 3.011
R35566 net2.n42 net2.n41 2.635
R35567 net2.n86 net2.n85 2.635
R35568 net2.n97 net2.n96 2.635
R35569 net2.n120 net2.n118 1.57
R35570 net2.n111 net2.n110 1.5
R35571 net2.n44 net2.n43 1.5
R35572 net2.n114 net2.n113 0.853
R35573 net2.n25 net2.n24 0.752
R35574 net2.n92 net2.n91 0.752
R35575 net2.n124 net2.n123 0.752
R35576 net2.n46 net2.n45 0.704
R35577 net2.n131 net2.n129 0.144
R35578 net2.n129 net2.n122 0.04
R35579 net2.n18 net2.n17 0.035
R35580 net2.n82 net2.n81 0.035
R35581 net2.n1 net2.n0 0.035
R35582 net2.n63 net2.n62 0.035
R35583 net2.n135 net2.n133 0.035
R35584 net2.n11 net2.n10 0.034
R35585 net2.n72 net2.n71 0.034
R35586 net2.n101 net2.n100 0.032
R35587 net2.n70 net2.n69 0.032
R35588 net2.n47 net2.n46 0.031
R35589 net2.n58 net2.n57 0.031
R35590 net2.n35 net2.n34 0.03
R35591 net2.n104 net2.n102 0.03
R35592 net2.n9 net2.n8 0.03
R35593 net2.n68 net2.n67 0.03
R35594 net2.n38 net2.n36 0.028
R35595 net2.n20 net2.n19 0.028
R35596 net2.n84 net2.n83 0.028
R35597 net2.n6 net2.n5 0.028
R35598 net2.n3 net2.n2 0.028
R35599 net2.n65 net2.n64 0.028
R35600 net2.n111 net2.n72 0.028
R35601 net2.n45 net2.n44 0.027
R35602 net2.n51 net2.n50 0.027
R35603 net2.n54 net2.n53 0.027
R35604 net2.n44 net2.n11 0.026
R35605 net2.n80 net2.n76 0.022
R35606 net2.n61 net2.n60 0.022
R35607 net2.n113 net2.n111 0.022
R35608 net2.n76 net2.n74 0.02
R35609 net2.n60 net2.n59 0.02
R35610 net2.n114 net2.n58 0.019
R35611 net2.n115 net2.n114 0.019
R35612 net2.n43 net2.n12 0.018
R35613 net2.n39 net2.n38 0.018
R35614 net2.n36 net2.n35 0.018
R35615 net2.n98 net2.n89 0.018
R35616 net2.n10 net2.n9 0.018
R35617 net2.n32 net2.n23 0.017
R35618 net2.n102 net2.n101 0.017
R35619 net2.n105 net2.n104 0.017
R35620 net2.n110 net2.n109 0.017
R35621 net2.n8 net2.n7 0.017
R35622 net2.n69 net2.n68 0.017
R35623 net2.n71 net2.n70 0.017
R35624 net2.n33 net2.n32 0.015
R35625 net2.n22 net2.n21 0.015
R35626 net2.n110 net2.n105 0.015
R35627 net2.n5 net2.n4 0.015
R35628 net2.n43 net2.n39 0.013
R35629 net2.n88 net2.n87 0.013
R35630 net2.n99 net2.n98 0.013
R35631 net2.n67 net2.n66 0.013
R35632 net2.n52 net2.n51 0.012
R35633 net2.n53 net2.n52 0.012
R35634 net2.n113 net2.n112 0.012
R35635 net2.n23 net2.n22 0.011
R35636 net2.n89 net2.n88 0.011
R35637 net2.n49 net2.n48 0.011
R35638 net2.n56 net2.n55 0.011
R35639 net2.n133 net2.n131 0.01
R35640 net2.n81 net2.n80 0.009
R35641 net2.n62 net2.n61 0.009
R35642 net2.n19 net2.n18 0.007
R35643 net2.n83 net2.n82 0.007
R35644 net2.n2 net2.n1 0.007
R35645 net2.n64 net2.n63 0.007
R35646 net2.n48 net2.n47 0.006
R35647 net2.n50 net2.n49 0.006
R35648 net2.n55 net2.n54 0.006
R35649 net2.n57 net2.n56 0.006
R35650 net2.n122 net2.n120 0.005
R35651 net2.n34 net2.n33 0.003
R35652 net2.n87 net2.n84 0.003
R35653 net2.n100 net2.n99 0.003
R35654 net2.n66 net2.n65 0.003
R35655 net2.n21 net2.n20 0.001
R35656 net2.n7 net2.n6 0.001
R35657 net2.n4 net2.n3 0.001
C0 a_15549_1034# net5 0.01fF
C1 a_23049_n8352# net4 0.06fF
C2 a_47405_2164# p_bais 0.02fF
C3 a_47558_n6837# net5_ota 0.04fF
C4 VDD Nbais 2.52fF
C5 VBN p_bais 3.78fF
C6 VBN net1 2.17fF
C7 p_bais net4 2.55fF
C8 UBP net6_ota 0.06fF
C9 net7 net3 5.26fF
C10 VBP net5 8.04fF
C11 a_37427_n9995# VDD 0.60fF
C12 net3 VOP 2.37fF
C13 net4 net1 3.00fF
C14 net6_ota net6 0.03fF
C15 net1_ota VON 0.09fF
C16 a_44684_n6035# net6_ota 0.01fF
C17 VON DNB 1.52fF
C18 VOP net5_ota 0.16fF
C19 a_34413_n132# VOP 0.05fF
C20 a_30462_n9995# net6 0.06fF
C21 a_25506_n10355# VOP 0.01fF
C22 VDD UP 5.78fF
C23 VBN Nbais 1.33fF
C24 VBP p_bais 3.15fF
C25 VDD VON 5.39fF
C26 p_bais net5 1.09fF
C27 VBN net2 0.53fF
C28 VBP net1 0.33fF
C29 Nbais net4 1.85fF
C30 net7 net6_ota 4.02fF
C31 net4 net2 1.05fF
C32 net3_ota VON 0.52fF
C33 net5 net1 0.42fF
C34 net6_ota VOP 1.10fF
C35 VOP DN 0.80fF
C36 a_30462_n9995# net7 0.20fF
C37 a_26106_n10355# net5 0.02fF
C38 a_15549_1034# Nbais 0.01fF
C39 a_49408_2164# net1_ota 0.07fF
C40 a_37408_3034# VDD 0.72fF
C41 VBN UP 3.05fF
C42 VDD UBP 4.92fF
C43 VBP Nbais 3.31fF
C44 Nbais net5 0.40fF
C45 VBN VON 4.60fF
C46 VDD net6 6.28fF
C47 VBP net2 0.02fF
C48 net3 net6_ota 0.51fF
C49 p_bais net1 1.01fF
C50 a_44684_n6035# VDD 0.31fF
C51 net5 net2 0.27fF
C52 net6_ota net5_ota 0.97fF
C53 net1_ota VOP 0.11fF
C54 VOP DNB 1.25fF
C55 a_25506_n10355# DN 0.02fF
C56 a_23049_n8352# Nbais 0.03fF
C57 a_49408_2164# VDD 0.38fF
C58 a_49408_2164# net3_ota 0.04fF
C59 a_30443_3034# net7 0.06fF
C60 VBP UP 0.14fF
C61 VBN UBP 1.82fF
C62 p_bais Nbais 1.38fF
C63 VDD net7 36.84fF
C64 Nbais net1 0.08fF
C65 VDD VOP 4.24fF
C66 p_bais net2 0.35fF
C67 UP net5 0.01fF
C68 VBP VON 4.51fF
C69 VBN net6 1.14fF
C70 a_44684_n6035# a_45884_n6035# 0.01fF
C71 net3_ota VOP 0.03fF
C72 net1 net2 1.83fF
C73 net5 VON 1.96fF
C74 a_33213_n132# VON 0.07fF
C75 VBN net7 1.12fF
C76 VDD net3 7.06fF
C77 p_bais UP 0.41fF
C78 p_bais VON 7.23fF
C79 VBP net6 7.47fF
C80 Nbais net2 0.19fF
C81 VBN VOP 3.01fF
C82 VDD net5_ota 0.56fF
C83 a_34413_n132# VDD 0.77fF
C84 DN DNB 4.30fF
C85 a_33213_n132# net6 0.03fF
C86 a_22549_1034# VBN 0.03fF
C87 a_26106_n10355# VON 0.02fF
C88 a_22549_1034# net4 0.05fF
C89 a_49058_n6837# VOP 0.03fF
C90 VDD net6_ota 5.08fF
C91 VBP net7 3.03fF
C92 VBN net3 0.87fF
C93 p_bais UBP 0.34fF
C94 VBN net5_ota 0.28fF
C95 VDD DN 0.67fF
C96 p_bais net6 4.97fF
C97 VBP VOP 1.98fF
C98 a_45884_n6035# net5_ota 0.02fF
C99 net5 VOP 1.32fF
C100 a_30462_n9995# VDD 0.57fF
C101 a_33213_n132# VOP 0.04fF
C102 a_22549_1034# net5 0.05fF
C103 a_47748_n2804# VDD 0.09fF
C104 VBN net6_ota 4.12fF
C105 VDD net1_ota 4.21fF
C106 VBP net3 1.63fF
C107 p_bais net7 8.64fF
C108 a_45884_n6035# net6_ota 0.02fF
C109 net3 net5 0.18fF
C110 p_bais VOP 6.01fF
C111 UP VON 0.18fF
C112 net1_ota net3_ota 4.89fF
C113 VDD DNB 0.41fF
C114 a_37427_n9995# net6 0.18fF
C115 a_33213_n132# a_34413_n132# 0.03fF
C116 a_26106_n10355# VOP 0.01fF
C117 a_48948_n2804# VDD 0.09fF
C118 a_25506_n10355# net5 0.02fF
C119 a_47405_2164# net1_ota 0.07fF
C120 a_30443_3034# VDD 0.75fF
C121 p_bais net3 7.27fF
C122 VBP net6_ota 0.50fF
C123 VDD net3_ota 3.35fF
C124 UP UBP 7.52fF
C125 UBP VON 0.02fF
C126 UP net6 0.05fF
C127 a_37427_n9995# net7 0.07fF
C128 VON net6 4.02fF
C129 net5 DN 0.06fF
C130 a_30462_n9995# VBP 0.01fF
C131 a_15049_n8352# Nbais 0.01fF
C132 a_47405_2164# VDD 0.38fF
C133 a_25506_n10355# a_26106_n10355# 0.02fF
C134 a_47405_2164# net3_ota 0.05fF
C135 VDD VBN 6.05fF
C136 a_45884_n6035# VDD 0.30fF
C137 p_bais net6_ota 1.18fF
C138 VBP net1_ota 0.11fF
C139 UP net7 0.04fF
C140 UBP net6 0.04fF
C141 UP VOP 0.02fF
C142 net7 VON 2.19fF
C143 w_4269_n7633# VDD 5.00fF
C144 net5 DNB 0.03fF
C145 VON VOP 13.08fF
C146 a_37408_3034# net7 0.17fF
C147 VDD VBP 9.33fF
C148 UP net3 0.49fF
C149 UBP net7 0.04fF
C150 VBP net3_ota 0.35fF
C151 p_bais net1_ota 1.02fF
C152 VBN net4 7.17fF
C153 net7 net6 23.07fF
C154 Nbais DN 1.04fF
C155 UBP VOP 0.12fF
C156 net3 VON 1.14fF
C157 net6 VOP 5.35fF
C158 VON net5_ota 0.13fF
C159 a_34413_n132# VON 0.03fF
C160 a_33213_n132# VDD 0.78fF
C161 a_26106_n10355# DNB 0.02fF
C162 a_15549_1034# VBN 0.02fF
C163 a_15549_1034# net4 0.07fF
C164 a_30443_3034# p_bais 0.06fF
C165 VBN VBP 3.12fF
C166 VDD p_bais 14.51fF
C167 VBP net4 0.38fF
C168 VBN net5 2.74fF
C169 UBP net3 0.79fF
C170 p_bais net3_ota 0.84fF
C171 net3 net6 2.26fF
C172 net4 net5 4.02fF
C173 net7 VOP 3.10fF
C174 net6_ota VON 1.50fF
C175 w_4269_n7633# VBP 2.47fF
C176 VON DN 0.09fF
C177 a_44684_n6035# net5_ota 0.01fF
C178 a_34413_n132# net6 0.04fF
.ends

