*** VCO Circuit implementation 

.subckt vco VDD GND vp vn vctrl ibias_vco 

** current mirrror cct**
M4 net1 ibias_vco VDD VDD sky130_fd_pr__pfet_01v8 L=0.5u W=1000u nf=50 m=1
M5 ibias_vco ibias_vco VDD VDD sky130_fd_pr__pfet_01v8 L=0.5u W=200u nf=10 m=1

** cross coupled cct**
M11 vp vn net1 net1 sky130_fd_pr__pfet_01v8 L=0.15u W=250u nf=5 m=1
M1 vn vp net1 net1 sky130_fd_pr__pfet_01v8 L=0.15u W=250u nf=5 m=1

M2 vp vn GND GND sky130_fd_pr__nfet_01v8 L=0.15u W=100u nf=5 m=1
M7 vn vp GND GND sky130_fd_pr__nfet_01v8 L=0.15u W=100u nf=5 m=1

** Varactor cct**
M6 vctrl vn vctrl gnd sky130_fd_pr__nfet_01v8_lvt L=8u W=17u nf=1 m=1
M3 vctrl vp vctrl gnd sky130_fd_pr__nfet_01v8_lvt L=8u W=17u nf=1 m=1

.ends