*** biasing Circuit implementation 

.subckt ind_model ind1 ind2
**************************************
*************ASTIC-hexa***************
**************************************
R0 net1 ind2 4.734 m=1
L1 ind1 net1 3.924n m=1

** R1 net2 ind2 2.367 m=1

C3 ind1 net3 11.14f m=10
R2 net3 GND 4.65 m=1

C2 ind2 net4 11.14f m=10
R3 net4 GND 4.65 m=1

**************************************
*************Original schematic*******
**************************************
** L1 vp net4 4n m=1
** R1 vp vn 1182 m=1
** R2 net4 vn 3 m=1
** C1 vp vn 5f m=10
** C3 vp GND 5f m=5
** C2 vn GND 5f m=5

** inductor model cct
**************************************
***** after modification *************
**************************************
** L1 vp net4 2.2n m=1
** R1 vp vn 678 m=1
** R2 net4 vn 1.7 m=1
** *C1 vp vn 5f m=10
** C3 vp GND 5f m=5
** C2 vn GND 5f m=5

**************************************
*************ASTIC********************
**************************************
** L1 vp net4 4.077n m=1
** R2 net4 vn 4.8 m=1
** 
** C3 vp netc3 11.8f m=10
** RC3 netc3 GND 4.65 m=1
** 
** C2 vn netc2 11.8f m=10
** RC2 netc2 GND 4.65 m=1

**************************************
*************Original*****************
**************************************
** L1 vp net4 4n m=1
** R1 vp vn 1182 m=1
** R2 net4 vn 3 m=1
** C1 vp vn 5f m=10
** C3 vp GND 5f m=5
** C2 vn GND 5f m=5

.ends