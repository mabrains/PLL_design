* NGSPICE file created from DIVIDER.eXMt - technology: sky130A

.subckt DIVIDER P0 P1 P2 P7 P6 P5 P4 P3 fin modo modi fout0 modi0 fout1 modi1 modi2
+ fout2 modi3 fout3 fout4 modi4 fout5 modi5 fout6 modi6 fout VDD GND
XM0 a_n3749_8439# fout2.t3 a_n4036_12366# GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=1.16e+12p ps=9.16e+06u W=2 L=0.15
XM1 a_n13930_2482# fout5.t3 a_n14130_2482# GND.t42 sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=3.48e+12p ps=2.516e+07u W=6 L=0.15
XM2 fout6.t2 a_n14423_5865.t4 a_n14633_2483# GND.t57 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.516e+07u W=6 L=0.15
XM3 VDD.t122 fin.t0 a_n24539_11543.t0 VDD.t121 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM4 GND.t97 fout6.t3 a_n15556_2475# GND.t96 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u W=2 L=0.15
XM5 a_n15024_8436# a_n15419_8436# VDD.t149 VDD.t148 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u W=4 L=0.15
XM6 a_n18023_11547# a_n18753_11548.t4 fout1.t1 GND sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=0p ps=0u W=6 L=0.15
XM7 a_n5255_5996# a_n6002_2899.t2 a_n5699_5899# VDD.t144 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=1.16e+12p ps=8.58e+06u W=4 L=0.15
XM8 a_n11277_8440# fout2.t4 VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u W=4 L=0.15
XM9 a_n11129_2476# fout4.t3 a_n11555_5898# GND.t121 sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=5.8e+11p ps=4.58e+06u W=2 L=0.15
XM10 GND a_n20158_11542.t3 a_n21540_12270.t1 GND sky130_fd_pr__nfet_01v8 ad=6.96e+13p pd=5.2176e+08u as=0p ps=0u W=2 L=0.15
XM11 GND a_n14372_11547.t3 a_n15755_12275.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM12 a_n17810_11459# a_n17562_12353.t2 a_n16468_12355# GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=1.16e+12p ps=9.16e+06u W=2 L=0.15
XM13 a_n10992_8440# fout1.t3 a_n11283_12359# GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=1.16e+12p ps=9.16e+06u W=2 L=0.15
XM14 a_n10596_8440# a_n10992_8440# VDD.t42 VDD.t41 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u W=4 L=0.15
XM15 a_n9889_12279.t0 a_n8507_11550.t3 VDD.t233 VDD.t232 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM16 a_n20386_2489# a_n22077_2481# GND.t85 GND.t84 sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=0p ps=0u W=6 L=0.15
XM17 a_n15419_8436# a_n17562_12353.t3 a_n15705_8436# VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=2.32e+12p ps=1.716e+07u W=4 L=0.15
XM18 VDD.t193 a_n18722_2907.t3 a_n18744_6000.t0 VDD.t192 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM19 VDD.t22 modi1.t2 a_n14372_11547.t0 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM20 a_n18744_6000.t1 a_n18722_2907.t4 GND.t44 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM21 modi0.t1 fout0.t3 a_n15024_8436# VDD.t85 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM22 a_n7001_2908.t1 modi4.t2 a_n6652_2485# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.516e+07u W=6 L=0.15
XM23 VDD.t64 a_n5699_5899# a_n5936_5996# VDD.t63 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.716e+07u W=4 L=0.15
XM24 GND modi1.t3 a_n12600_11551# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.516e+07u W=6 L=0.15
XM25 a_n14423_5865.t2 fout5.t4 VDD.t142 VDD.t141 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM26 GND a_n2702_11550.t3 a_n4084_12278.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM27 a_n21491_8431# a_n21540_12270.t2 VDD.t84 VDD.t83 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u W=4 L=0.15
XM28 a_n15419_8436# fout0.t4 a_n15707_12363# GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=1.16e+12p ps=9.16e+06u W=2 L=0.15
XM29 GND fout1.t4 a_n14284_11547# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.516e+07u W=6 L=0.15
XM30 a_n22643_8431# fin.t1 a_n22934_12350# GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=1.16e+12p ps=9.16e+06u W=2 L=0.15
XM31 a_n9554_8440# a_n11697_12356.t2 a_n9840_8440# VDD.t145 sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=2.32e+12p ps=1.716e+07u W=4 L=0.15
XM32 VDD.t50 a_n23172_5903# a_n23409_6000# VDD.t49 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.716e+07u W=4 L=0.15
XM33 a_n2913_2485# a_n4604_2477# GND.t48 GND.t47 sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=0p ps=0u W=6 L=0.15
XM34 GND modi2.t2 a_n6795_11551# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.516e+07u W=6 L=0.15
XM35 a_n23348_12347.t0 fin.t2 VDD.t120 VDD.t119 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM36 a_n12857_2907.t2 modi5.t2 VDD.t46 VDD.t45 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM37 a_n4516_2477# a_n6002_2899.t3 a_n4604_2477# GND.t87 sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=5.8e+11p ps=4.58e+06u W=2 L=0.15
XM38 a_n24497_6006.t1 a_n24474_2912.t3 GND.t110 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM39 GND a_n6140_11462# a_n6353_11550# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.516e+07u W=6 L=0.15
XM40 VDD.t235 a_n11944_11462# fout2.t2 VDD.t234 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM41 VDD.t66 a_n24497_6006.t2 a_n22728_6000# VDD.t65 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.716e+07u W=4 L=0.15
XM42 GND.t92 a_n7023_6002.t2 a_n5273_2477# GND.t91 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u W=2 L=0.15
XM43 a_n21540_12270.t0 a_n20158_11542.t4 VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM44 a_n3835_2477# fout3.t3 a_n4261_5899# GND.t102 sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=5.8e+11p ps=4.58e+06u W=2 L=0.15
XM45 GND.t30 fout.t3 a_n21308_2481# GND.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u W=2 L=0.15
XM46 VDD.t87 fout0.t5 a_n18753_11548.t1 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM47 GND.t41 a_n5699_5899# a_n5954_2477# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u W=2 L=0.15
XM48 a_n9841_12367# a_n9889_12279.t2 GND GND sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u W=2 L=0.15
XM49 VDD.t237 a_n17419_5897# a_n17657_5994# VDD.t236 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.716e+07u W=4 L=0.15
XM50 VDD.t140 fout5.t5 a_n9674_5995# VDD.t139 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.716e+07u W=4 L=0.15
XM51 a_n9554_8440# fout1.t5 a_n9841_12367# GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u W=2 L=0.15
XM52 a_n8558_5866.t0 modi4.t3 VDD.t107 VDD.t106 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM53 VDD.t132 fout6.t4 a_n15538_5994# VDD.t131 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.716e+07u W=4 L=0.15
XM54 VDD.t166 a_n12888_11551.t4 fout2.t0 VDD.t165 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM55 VDD.t95 modi2.t3 a_n7083_11551.t2 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM56 a_n12880_6001.t1 a_n12857_2907.t3 GND.t120 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM57 a_n6353_11550# a_n7083_11551.t4 fout3.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM58 a_n20175_5871.t1 P7.t0 VDD.t105 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM59 a_n6002_2899.t0 fout3.t4 GND.t104 GND.t103 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM60 fout5.t2 a_n10460_2476# VDD.t191 VDD.t190 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM61 a_n16237_2475# a_n17722_2897.t2 a_n16325_2475# GND.t78 sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=5.8e+11p ps=4.58e+06u W=2 L=0.15
XM62 a_n19682_2488# fout6.t5 a_n19882_2488# GND.t98 sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=3.48e+12p ps=2.516e+07u W=6 L=0.15
XM63 a_n20815_12350# a_n21205_8431# GND GND sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u W=2 L=0.15
XM64 a_n20175_5871.t3 modi6.t2 VDD.t175 VDD.t174 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM65 fout5.t0 a_n8558_5866.t4 a_n8769_2484# GND.t101 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.516e+07u W=6 L=0.15
XM66 a_n15556_2475# fout5.t6 a_n15981_5897# GND.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u W=2 L=0.15
XM67 a_n8419_11550# modi2.t4 a_n8507_11550.t1 GND sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=0p ps=0u W=6 L=0.15
XM68 a_n18665_11548# P1.t0 a_n18753_11548.t3 GND sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=0p ps=0u W=6 L=0.15
XM69 a_n17143_8436# fout1.t6 VDD.t185 VDD.t184 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u W=4 L=0.15
XM70 a_n2209_2484# fout3.t5 a_n2409_2484# GND.t105 sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=3.48e+12p ps=2.516e+07u W=6 L=0.15
XM71 GND fout1.t7 a_n11697_12356.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM72 VDD.t72 a_n24539_11543.t4 fout0.t1 VDD.t71 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM73 a_n16462_8436# a_n16857_8436# VDD.t214 VDD.t213 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u W=4 L=0.15
XM74 a_n18722_2907.t0 modi6.t3 VDD.t89 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM75 GND fout0.t6 a_n20070_11542# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.516e+07u W=6 L=0.15
XM76 a_n17149_12355# fout1.t8 GND GND sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u W=2 L=0.15
XM77 VDD.t187 a_n12857_2907.t4 a_n12880_6001.t0 VDD.t186 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM78 GND fout3.t6 a_n2614_11550# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.516e+07u W=6 L=0.15
XM79 VDD.t157 a_n7083_11551.t5 fout3.t2 VDD.t156 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM80 GND fout2.t5 a_n5892_12356.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM81 fout6.t0 a_n16325_2475# VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM82 a_n7001_2908.t2 fout4.t4 VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM83 a_n16857_8436# a_n17562_12353.t4 a_n17143_8436# VDD.t108 sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u W=4 L=0.15
XM84 a_n17562_12353.t0 fout0.t7 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM85 VDD.t18 fout2.t6 a_n8507_11550.t0 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM86 a_n11112_5995# a_n11858_2898.t2 a_n11555_5898# VDD.t162 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=1.16e+12p ps=8.58e+06u W=4 L=0.15
XM87 a_n8266_2483# modi4.t4 GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=0p ps=0u W=6 L=0.15
XM88 VDD.t206 fout1.t9 a_n12888_11551.t2 VDD.t205 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM89 fout.t0 a_n20175_5871.t4 VDD.t110 VDD.t109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM90 a_n12857_2907.t0 fout5.t7 VDD.t138 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM91 a_n22253_12350# a_n22643_8431# GND GND sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u W=2 L=0.15
XM92 a_n4797_12358# a_n5187_8439# GND GND sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u W=2 L=0.15
XM93 a_n23475_2903.t1 fout6.t6 GND.t94 GND.t93 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM94 a_n2702_5867.t0 fout3.t7 VDD.t177 VDD.t176 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM95 a_n15707_12363# a_n15755_12275.t2 GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM96 a_n22928_8431# fout0.t8 VDD.t28 VDD.t27 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u W=4 L=0.15
XM97 a_n21989_2481# a_n23475_2903.t2 a_n22077_2481# GND.t88 sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=5.8e+11p ps=4.58e+06u W=2 L=0.15
XM98 VDD.t8 a_n10117_5898# a_n10355_5995# VDD.t7 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.716e+07u W=4 L=0.15
XM99 VDD.t70 a_n11555_5898# a_n11793_5995# VDD.t69 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.716e+07u W=4 L=0.15
XM100 a_n5954_2477# a_n6002_2899.t4 modi3.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM101 a_n21308_2481# fout6.t7 a_n21734_5903# GND.t128 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u W=2 L=0.15
XM102 GND.t28 a_n23172_5903# a_n23427_2481# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u W=2 L=0.15
XM103 VDD.t80 a_n12880_6001.t2 a_n11112_5995# VDD.t79 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM104 a_n10602_12359# a_n10992_8440# GND GND sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u W=2 L=0.15
XM105 VDD.t130 fout6.t8 a_n23475_2903.t0 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM106 a_n9164_12359# a_n9554_8440# GND GND sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u W=2 L=0.15
XM107 fout4.t2 a_n2702_5867.t4 VDD.t204 VDD.t203 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM108 VDD.t179 fout3.t8 a_n6002_2899.t1 VDD.t178 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM109 a_n4036_12366# a_n4084_12278.t2 GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM110 a_n17810_11459# fout0.t9 a_n16462_8436# VDD.t198 sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u W=4 L=0.15
XM111 a_n18722_2907.t2 modi6.t4 a_n18372_2483# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.516e+07u W=6 L=0.15
XM112 a_n4498_5996# fout3.t9 a_n4604_2477# VDD.t180 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=1.16e+12p ps=8.58e+06u W=4 L=0.15
XM113 GND fout0.t10 a_n17562_12353.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM114 VDD.t101 modi0.t2 a_n20158_11542.t1 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM115 a_n24474_2912.t1 modi.t0 VDD.t74 VDD.t73 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM116 a_n18465_11548# fout0.t11 a_n18665_11548# GND sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=0p ps=0u W=6 L=0.15
XM117 modi2.t1 a_n5892_12356.t2 a_n3360_12358# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u W=2 L=0.15
XM118 a_n3817_5996# a_n6002_2899.t5 a_n4261_5899# VDD.t217 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=1.16e+12p ps=8.58e+06u W=4 L=0.15
XM119 modo.t1 a_n23348_12347.t2 a_n20815_12350# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM120 a_n10992_8440# a_n11697_12356.t3 a_n11277_8440# VDD.t173 sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u W=4 L=0.15
XM121 a_n12157_11550# a_n12888_11551.t5 fout2.t1 GND sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=0p ps=0u W=6 L=0.15
XM122 a_n9840_8440# a_n9889_12279.t3 VDD.t48 VDD.t47 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM123 a_n21972_6000# fout6.t9 a_n22077_2481# VDD.t128 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=1.16e+12p ps=8.58e+06u W=4 L=0.15
XM124 a_n14633_2483# a_n16325_2475# GND.t23 GND.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM125 a_n24451_11543# P0.t0 a_n24539_11543.t2 GND sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=0p ps=0u W=6 L=0.15
XM126 a_n11944_11462# fout1.t10 a_n10596_8440# VDD.t207 sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u W=4 L=0.15
XM127 a_n17674_2475# a_n17722_2897.t3 modi5.t0 GND sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u W=2 L=0.15
XM128 a_n3360_12358# a_n3749_8439# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM129 a_n11697_12356.t0 fout1.t11 VDD.t209 VDD.t208 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM130 a_n18722_2907.t1 fout6.t10 VDD.t127 VDD.t126 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM131 a_n14423_5865.t3 P6.t0 a_n13930_2482# GND.t135 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM132 a_n24125_2489# fout.t4 GND.t31 GND sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=0p ps=0u W=6 L=0.15
XM133 VDD.t197 fout0.t12 a_n20158_11542.t2 VDD.t196 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM134 a_n21291_6000# a_n23475_2903.t3 a_n21734_5903# VDD.t215 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=1.16e+12p ps=8.58e+06u W=4 L=0.15
XM135 VDD.t151 modo.t2 a_n24539_11543.t1 VDD.t150 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM136 a_n5273_2477# fout3.t10 a_n5699_5899# GND.t114 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u W=2 L=0.15
XM137 GND.t154 a_n17419_5897# a_n17674_2475# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM138 VDD.t155 a_n18753_11548.t5 fout1.t2 VDD.t154 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM139 a_n4035_8439# a_n4084_12278.t3 VDD.t170 VDD.t169 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u W=4 L=0.15
XM140 a_n16219_5994# fout5.t8 a_n16325_2475# VDD.t136 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=1.16e+12p ps=8.58e+06u W=4 L=0.15
XM141 GND.t69 fout5.t9 a_n9691_2476# GND.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u W=2 L=0.15
XM142 GND a_n23595_11454# a_n23808_11542# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.516e+07u W=6 L=0.15
XM143 a_n5473_8439# fout3.t11 VDD.t182 VDD.t181 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u W=4 L=0.15
XM144 GND a_n11944_11462# a_n12157_11550# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM145 a_n21205_8431# a_n23348_12347.t3 a_n21491_8431# VDD.t201 sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u W=4 L=0.15
XM146 a_n14284_11547# modi1.t4 a_n14372_11547.t2 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM147 VDD.t239 P0.t1 a_n24539_11543.t3 VDD.t238 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM148 a_n4792_8439# a_n5187_8439# VDD.t195 VDD.t194 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u W=4 L=0.15
XM149 a_n3354_8439# a_n3749_8439# VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u W=4 L=0.15
XM150 a_n15538_5994# a_n17722_2897.t4 a_n15981_5897# VDD.t222 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u W=4 L=0.15
XM151 VDD.t36 a_n21734_5903# a_n21972_6000# VDD.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM152 modo.t0 fin.t3 a_n20810_8431# VDD.t118 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.716e+07u W=4 L=0.15
XM153 a_n6652_2485# fout4.t5 GND.t18 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM154 a_n17722_2897.t1 fout5.t10 GND.t71 GND.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM155 fout.t2 a_n22077_2481# VDD.t116 VDD.t115 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM156 VDD.t76 P3.t0 a_n7083_11551.t1 VDD.t75 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM157 a_n6140_11462# a_n5892_12356.t3 a_n4797_12358# GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u W=2 L=0.15
XM158 a_n3749_8439# a_n5892_12356.t4 a_n4035_8439# VDD.t55 sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u W=4 L=0.15
XM159 a_n21492_12358# a_n21540_12270.t3 GND GND sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u W=2 L=0.15
XM160 VDD.t114 a_n6140_11462# fout3.t0 VDD.t113 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM161 a_n5892_12356.t0 fout2.t7 VDD.t16 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM162 a_n14423_5865.t1 P6.t1 VDD.t78 VDD.t77 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM163 fout6.t1 a_n14423_5865.t5 VDD.t93 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM164 a_n7001_2908.t0 modi4.t5 VDD.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM165 a_n16857_8436# fout0.t13 a_n17149_12355# GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u W=2 L=0.15
XM166 a_n15030_12355# a_n15419_8436# GND GND sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u W=2 L=0.15
XM167 a_n23427_2481# a_n23475_2903.t4 modi6.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM168 GND modi0.t3 a_n18465_11548# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM169 a_n11944_11462# a_n11697_12356.t4 a_n10602_12359# GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u W=2 L=0.15
XM170 GND.t46 a_n24497_6006.t3 a_n22746_2481# GND.t45 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u W=2 L=0.15
XM171 fout4.t0 a_n4604_2477# VDD.t68 VDD.t67 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM172 a_n12857_2907.t1 modi5.t3 a_n12508_2484# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.516e+07u W=6 L=0.15
XM173 a_n18372_2483# fout6.t11 GND.t95 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM174 a_n22746_2481# fout6.t12 a_n23172_5903# GND.t153 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u W=2 L=0.15
XM175 VDD.t103 modi0.t4 a_n18753_11548.t2 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM176 a_n20070_11542# modi0.t5 a_n20158_11542.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM177 GND.t107 a_n15981_5897# a_n16237_2475# GND.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM178 a_n24251_11543# fin.t4 a_n24451_11543# GND sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=0p ps=0u W=6 L=0.15
XM179 a_n6995_11551# P3.t1 a_n7083_11551.t3 GND sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=0p ps=0u W=6 L=0.15
XM180 a_n15705_8436# a_n15755_12275.t3 VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM181 VDD.t172 a_n24474_2912.t4 a_n24497_6006.t0 VDD.t171 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM182 a_n5187_8439# fout2.t8 a_n5478_12358# GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=1.16e+12p ps=9.16e+06u W=2 L=0.15
XM183 VDD.t57 fout3.t12 a_n2702_11550.t0 VDD.t56 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM184 a_n8558_5866.t2 fout4.t6 VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM185 VDD.t44 P1.t1 a_n18753_11548.t0 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM186 a_n5936_5996# fout3.t13 modi3.t0 VDD.t58 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM187 modi0.t0 a_n17562_12353.t5 a_n15030_12355# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM188 a_n11810_2476# a_n11858_2898.t3 modi4.t0 GND sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u W=2 L=0.15
XM189 a_n23595_11454# a_n23348_12347.t4 a_n22253_12350# GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u W=2 L=0.15
XM190 VDD.t54 a_n17810_11459# fout1.t0 VDD.t53 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM191 a_n10372_2476# a_n11858_2898.t4 a_n10460_2476# GND.t115 sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=5.8e+11p ps=4.58e+06u W=2 L=0.15
XM192 a_n2614_11550# modi3.t2 a_n2702_11550.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM193 a_n8769_2484# a_n10460_2476# GND.t125 GND.t124 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM194 GND.t51 a_n12880_6001.t3 a_n11129_2476# GND.t50 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM195 a_n20175_5871.t0 P7.t1 a_n19682_2488# GND.t155 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM196 VDD.t14 fout2.t9 a_n7083_11551.t0 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM197 a_n23409_6000# fout6.t13 modi6.t1 VDD.t125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM198 a_n20175_5871.t2 fout6.t14 VDD.t124 VDD.t123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM199 GND.t7 a_n10117_5898# a_n10372_2476# GND.t6 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM200 GND.t49 a_n11555_5898# a_n11810_2476# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM201 a_n22247_8431# a_n22643_8431# VDD.t40 VDD.t39 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u W=4 L=0.15
XM202 a_n12800_11551# P2.t0 a_n12888_11551.t0 GND sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=0p ps=0u W=6 L=0.15
XM203 a_n4084_12278.t0 a_n2702_11550.t4 VDD.t189 VDD.t188 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM204 a_n9691_2476# fout4.t7 a_n10117_5898# GND.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u W=2 L=0.15
XM205 a_n19882_2488# modi6.t5 GND.t134 GND.t133 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM206 a_n22728_6000# a_n23475_2903.t5 a_n23172_5903# VDD.t216 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u W=4 L=0.15
XM207 a_n2702_5867.t1 P4.t0 a_n2209_2484# GND.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM208 fout5.t1 a_n8558_5866.t5 VDD.t164 VDD.t163 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM209 VDD.t225 fout4.t8 a_n11858_2898.t0 VDD.t224 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM210 GND a_n17810_11459# a_n18023_11547# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM211 modi1.t1 a_n11697_12356.t5 a_n9164_12359# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM212 a_n17657_5994# fout5.t11 modi5.t1 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM213 a_n22643_8431# a_n23348_12347.t5 a_n22928_8431# VDD.t202 sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u W=4 L=0.15
XM214 a_n2409_2484# modi3.t3 GND.t146 GND.t145 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM215 a_n9674_5995# a_n11858_2898.t5 a_n10117_5898# VDD.t183 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u W=4 L=0.15
XM216 GND a_n8507_11550.t4 a_n9889_12279.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM217 a_n11858_2898.t1 fout4.t9 GND.t143 GND.t142 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM218 a_n5478_12358# fout3.t14 GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM219 a_n23595_11454# fin.t5 a_n22247_8431# VDD.t117 sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u W=4 L=0.15
XM220 VDD.t231 a_n23595_11454# fout0.t2 VDD.t230 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM221 VDD.t159 modi2.t5 a_n8507_11550.t2 VDD.t158 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM222 GND.t21 a_n21734_5903# a_n21989_2481# GND.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM223 a_n8558_5866.t3 P5.t0 VDD.t221 VDD.t220 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM224 a_n9159_8440# a_n9554_8440# VDD.t60 VDD.t59 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u W=4 L=0.15
XM225 a_n8066_2483# fout4.t10 a_n8266_2483# GND.t144 sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=0p ps=0u W=6 L=0.15
XM226 VDD.t168 a_n15981_5897# a_n16219_5994# VDD.t167 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM227 a_n16993_2475# fout5.t12 a_n17419_5897# GND.t66 sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=5.8e+11p ps=4.58e+06u W=2 L=0.15
XM228 VDD.t112 a_n4261_5899# a_n4498_5996# VDD.t111 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM229 GND modo.t3 a_n24251_11543# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM230 a_n16468_12355# a_n16857_8436# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM231 VDD.t200 modi1.t5 a_n12888_11551.t3 VDD.t199 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM232 a_n2702_5867.t2 P4.t1 VDD.t147 VDD.t146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM233 a_n11283_12359# fout2.t10 GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM234 GND fout2.t11 a_n8419_11550# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM235 a_n12508_2484# fout5.t13 GND.t67 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM236 a_n14130_2482# modi5.t4 GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM237 fout.t1 a_n20175_5871.t5 a_n20386_2489# GND.t79 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM238 VDD.t153 a_n7023_6002.t3 a_n5255_5996# VDD.t152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM239 VDD.t227 fout4.t11 a_n3817_5996# VDD.t226 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM240 VDD.t211 fout1.t12 a_n14372_11547.t1 VDD.t210 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM241 VDD.t97 P2.t1 a_n12888_11551.t1 VDD.t96 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM242 a_n16976_5994# a_n17722_2897.t5 a_n17419_5897# VDD.t223 sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=1.16e+12p ps=8.58e+06u W=4 L=0.15
XM243 VDD.t134 fout5.t14 a_n17722_2897.t0 VDD.t133 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM244 a_n2702_5867.t3 modi3.t4 VDD.t219 VDD.t218 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM245 a_n20810_8431# a_n21205_8431# VDD.t82 VDD.t81 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM246 VDD.t229 modi3.t5 a_n2702_11550.t2 VDD.t228 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM247 a_n21205_8431# fin.t6 a_n21492_12358# GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u W=2 L=0.15
XM248 a_n15755_12275.t0 a_n14372_11547.t4 VDD.t91 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM249 VDD.t52 fout.t5 a_n21291_6000# VDD.t51 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM250 modi1.t0 fout1.t13 a_n9159_8440# VDD.t212 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM251 a_n7023_6002.t1 a_n7001_2908.t3 GND.t40 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM252 a_n22934_12350# fout0.t14 GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM253 a_n12600_11551# fout1.t14 a_n12800_11551# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM254 GND.t81 a_n4261_5899# a_n4516_2477# GND.t80 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM255 a_n23808_11542# a_n24539_11543.t5 fout0.t0 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM256 a_n5187_8439# a_n5892_12356.t5 a_n5473_8439# VDD.t143 sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u W=4 L=0.15
XM257 fout4.t1 a_n2702_5867.t5 a_n2913_2485# GND.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM258 GND fin.t7 a_n23348_12347.t1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM259 GND.t73 fout4.t12 a_n3835_2477# GND.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM260 a_n6140_11462# fout2.t12 a_n4792_8439# VDD.t12 sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u W=4 L=0.15
XM261 modi2.t0 fout2.t13 a_n3354_8439# VDD.t11 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM262 VDD.t161 a_n18744_6000.t2 a_n16976_5994# VDD.t160 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM263 a_n24474_2912.t2 modi.t1 a_n24125_2489# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM264 a_n6795_11551# fout2.t14 a_n6995_11551# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM265 a_n14423_5865.t0 modi5.t5 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM266 a_n8558_5866.t1 P5.t1 a_n8066_2483# GND.t111 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=6 L=0.15
XM267 GND.t148 a_n18744_6000.t3 a_n16993_2475# GND.t147 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u W=2 L=0.15
XM268 a_n10355_5995# fout4.t13 a_n10460_2476# VDD.t98 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u W=4 L=0.15
XM269 a_n24474_2912.t0 fout.t6 VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM270 a_n11793_5995# fout4.t14 modi4.t1 VDD.t99 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
XM271 VDD.t62 a_n7001_2908.t4 a_n7023_6002.t0 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u W=4 L=0.15
R0 fout2.n109 fout2.t14 1038.92
R1 fout2.n139 fout2.t11 1037.29
R2 fout2.n140 fout2.t6 797.225
R3 fout2.n125 fout2.t9 795.548
R4 fout2.n509 fout2.t4 732.329
R5 fout2.n37 fout2.t13 731.671
R6 fout2.n12 fout2.t12 731.671
R7 fout2.n0 fout2.t7 730.667
R8 fout2.n86 fout2.t8 400.616
R9 fout2.n57 fout2.t3 400.598
R10 fout2.n524 fout2.t10 397.317
R11 fout2.n0 fout2.t5 395.829
R12 fout2.n349 fout2.n348 13.176
R13 fout2.n161 fout2.t2 11.718
R14 fout2.n161 fout2.t0 10.996
R15 fout2.n169 fout2.n167 9.3
R16 fout2.n471 fout2.n470 9.3
R17 fout2.n217 fout2.n216 9.3
R18 fout2.n219 fout2.n218 9.3
R19 fout2.n276 fout2.n275 9.3
R20 fout2.n273 fout2.n272 9.3
R21 fout2.n231 fout2.n230 9.3
R22 fout2.n229 fout2.n228 9.3
R23 fout2.n355 fout2.n354 9.3
R24 fout2.n254 fout2.n253 9.3
R25 fout2.n262 fout2.n261 9.3
R26 fout2.n265 fout2.n264 9.3
R27 fout2.n385 fout2.n384 9.3
R28 fout2.n382 fout2.n381 9.3
R29 fout2.n466 fout2.n465 9.3
R30 fout2.n464 fout2.n463 9.3
R31 fout2.n457 fout2.n456 8.097
R32 fout2.n264 fout2.n263 5.457
R33 fout2.n384 fout2.n383 5.08
R34 fout2.n455 fout2.n454 4.65
R35 fout2.n394 fout2.n393 4.65
R36 fout2.n476 fout2.n469 4.5
R37 fout2.n450 fout2.n449 4.5
R38 fout2.n443 fout2.n442 4.5
R39 fout2.n374 fout2.n373 4.5
R40 fout2.n364 fout2.n363 4.5
R41 fout2.n351 fout2.n350 4.5
R42 fout2.n327 fout2.n326 4.5
R43 fout2.n259 fout2.n251 4.5
R44 fout2.n282 fout2.n281 4.5
R45 fout2.n227 fout2.n226 4.5
R46 fout2.n239 fout2.n238 4.5
R47 fout2.n246 fout2.n245 4.5
R48 fout2.n290 fout2.n289 4.5
R49 fout2.n270 fout2.n269 4.5
R50 fout2.n436 fout2.n435 4.5
R51 fout2.n215 fout2.n214 4.5
R52 fout2.n485 fout2.n482 4.5
R53 fout2.n172 fout2.n171 4.5
R54 fout2.n238 fout2.n236 4.314
R55 fout2.n289 fout2.n286 3.944
R56 fout2.n449 fout2.n448 3.937
R57 fout2.n435 fout2.n434 3.567
R58 fout2.n395 fout2.n388 3.033
R59 fout2.n459 fout2.n458 3.033
R60 fout2.n456 fout2.t1 2.9
R61 fout2.n288 fout2.n287 2.258
R62 fout2.n433 fout2.n432 2.258
R63 fout2.n244 fout2.n243 1.882
R64 fout2.n245 fout2.n244 1.882
R65 fout2.n441 fout2.n440 1.882
R66 fout2.n497 fout2.n161 1.516
R67 fout2.n435 fout2.n433 1.505
R68 fout2.n442 fout2.n441 1.505
R69 fout2.n477 fout2.n476 1.5
R70 fout2.n328 fout2.n327 1.5
R71 fout2.n365 fout2.n364 1.5
R72 fout2.n396 fout2.n395 1.5
R73 fout2.n375 fout2.n374 1.5
R74 fout2.n486 fout2.n485 1.5
R75 fout2.n173 fout2.n172 1.5
R76 fout2.n46 fout2.n45 1.435
R77 fout2.n75 fout2.n74 1.435
R78 fout2.n153 fout2.n139 1.388
R79 fout2.n111 fout2.n109 1.355
R80 fout2.n126 fout2.n125 1.355
R81 fout2.n141 fout2.n140 1.354
R82 fout2.n526 fout2.n524 1.354
R83 fout2.n510 fout2.n509 1.354
R84 fout2.n38 fout2.n37 1.354
R85 fout2.n13 fout2.n12 1.354
R86 fout2.n112 fout2.n111 1.142
R87 fout2.n39 fout2.n38 1.142
R88 fout2.n14 fout2.n13 1.142
R89 fout2.n527 fout2.n526 1.142
R90 fout2.n40 fout2.n39 1.138
R91 fout2.n69 fout2.n14 1.138
R92 fout2.n113 fout2.n112 1.138
R93 fout2.n528 fout2.n527 1.138
R94 fout2.n511 fout2.n510 1.137
R95 fout2.n537 fout2.n536 1.137
R96 fout2.n502 fout2.n501 1.137
R97 fout2.n532 fout2.n531 1.137
R98 fout2.n517 fout2.n516 1.137
R99 fout2.n23 fout2.n22 1.137
R100 fout2.n52 fout2.n51 1.137
R101 fout2.n18 fout2.n17 1.137
R102 fout2.n29 fout2.n28 1.137
R103 fout2.n47 fout2.n46 1.137
R104 fout2.n66 fout2.n65 1.137
R105 fout2.n81 fout2.n80 1.137
R106 fout2.n62 fout2.n61 1.137
R107 fout2.n4 fout2.n3 1.137
R108 fout2.n76 fout2.n75 1.137
R109 fout2.n127 fout2.n126 1.137
R110 fout2.n95 fout2.n94 1.137
R111 fout2.n118 fout2.n117 1.137
R112 fout2.n91 fout2.n90 1.137
R113 fout2.n102 fout2.n101 1.137
R114 fout2.n97 fout2.n96 1.136
R115 fout2.n539 fout2.n538 1.136
R116 fout2.n129 fout2.n128 1.136
R117 fout2.n84 fout2.n83 1.136
R118 fout2.n68 fout2.n67 1.136
R119 fout2.n55 fout2.n54 1.136
R120 fout2.n25 fout2.n24 1.136
R121 fout2.n513 fout2.n512 1.136
R122 fout2.n214 fout2.n213 1.129
R123 fout2.n289 fout2.n288 1.129
R124 fout2.n281 fout2.n280 1.129
R125 fout2.n291 fout2.n290 1.042
R126 fout2.n308 fout2.n307 0.853
R127 fout2.n398 fout2.n397 0.853
R128 fout2.n492 fout2.n491 0.853
R129 fout2.n185 fout2.n184 0.853
R130 fout2.n541 fout2.n160 0.827
R131 fout2.n171 fout2.n170 0.752
R132 fout2.n363 fout2.n362 0.752
R133 fout2.n373 fout2.n372 0.752
R134 fout2.n449 fout2.n447 0.752
R135 fout2.n469 fout2.n468 0.752
R136 fout2.n482 fout2.n481 0.752
R137 fout2.n175 fout2.n174 0.717
R138 fout2.n497 fout2.n496 0.689
R139 fout2.n498 fout2.n497 0.68
R140 fout2.n354 fout2.n353 0.536
R141 fout2.n253 fout2.n252 0.536
R142 fout2.n275 fout2.n274 0.475
R143 fout2.n393 fout2.n392 0.475
R144 fout2.n541 fout2.n540 0.47
R145 fout2.n154 fout2.n153 0.44
R146 fout2.n458 fout2.n457 0.382
R147 fout2.n225 fout2.n224 0.382
R148 fout2.n226 fout2.n225 0.376
R149 fout2.n238 fout2.n237 0.376
R150 fout2.n269 fout2.n268 0.376
R151 fout2.n251 fout2.n250 0.376
R152 fout2.n326 fout2.n325 0.376
R153 fout2.n350 fout2.n349 0.376
R154 fout2.n213 fout2.n212 0.349
R155 fout2.n468 fout2.n467 0.349
R156 fout2 fout2.n130 0.213
R157 fout2.n88 fout2.n87 0.152
R158 fout2.n57 fout2.n56 0.123
R159 fout2.n86 fout2.n85 0.123
R160 fout2.n58 fout2.n57 0.091
R161 fout2 fout2.n541 0.086
R162 fout2.n524 fout2.n523 0.083
R163 fout2.n509 fout2.n508 0.083
R164 fout2.n37 fout2.n36 0.083
R165 fout2.n12 fout2.n11 0.083
R166 fout2.n139 fout2.n138 0.076
R167 fout2.n109 fout2.n108 0.075
R168 fout2.n125 fout2.n124 0.075
R169 fout2.n87 fout2.n86 0.07
R170 fout2.n135 fout2.n134 0.059
R171 fout2.n266 fout2.n265 0.047
R172 fout2.n256 fout2.n255 0.047
R173 fout2.n345 fout2.n344 0.047
R174 fout2.n358 fout2.n357 0.047
R175 fout2.n386 fout2.n385 0.047
R176 fout2.n473 fout2.n472 0.047
R177 fout2.n452 fout2.n451 0.043
R178 fout2.n421 fout2.n420 0.043
R179 fout2.n235 fout2.n234 0.041
R180 fout2.n202 fout2.n201 0.041
R181 fout2.n461 fout2.n460 0.035
R182 fout2.n329 fout2.n328 0.035
R183 fout2.n334 fout2.n333 0.035
R184 fout2.n427 fout2.n426 0.035
R185 fout2.n222 fout2.n221 0.034
R186 fout2.n343 fout2.n342 0.034
R187 fout2.n347 fout2.n346 0.034
R188 fout2.n464 fout2.n462 0.034
R189 fout2.n182 fout2.n181 0.034
R190 fout2.n180 fout2.n179 0.034
R191 fout2.n298 fout2.n297 0.034
R192 fout2.n305 fout2.n304 0.034
R193 fout2.n365 fout2.n341 0.034
R194 fout2.n367 fout2.n366 0.034
R195 fout2.n380 fout2.n379 0.034
R196 fout2.n429 fout2.n428 0.034
R197 fout2.n149 fout2.n148 0.032
R198 fout2.n148 fout2.n147 0.032
R199 fout2.n536 fout2.n534 0.032
R200 fout2.n22 fout2.n20 0.032
R201 fout2.n61 fout2.n60 0.032
R202 fout2.n94 fout2.n92 0.032
R203 fout2.n220 fout2.n219 0.032
R204 fout2.n395 fout2.n394 0.032
R205 fout2.n459 fout2.n455 0.032
R206 fout2.n303 fout2.n302 0.032
R207 fout2.n477 fout2.n429 0.032
R208 fout2.n153 fout2.n152 0.032
R209 fout2.n187 fout2.n186 0.031
R210 fout2.n198 fout2.n197 0.031
R211 fout2.n310 fout2.n309 0.031
R212 fout2.n321 fout2.n320 0.031
R213 fout2.n400 fout2.n399 0.031
R214 fout2.n411 fout2.n410 0.031
R215 fout2.n494 fout2.n493 0.031
R216 fout2.n143 fout2.n142 0.03
R217 fout2.n229 fout2.n227 0.03
R218 fout2.n273 fout2.n271 0.03
R219 fout2.n258 fout2.n257 0.03
R220 fout2.n360 fout2.n359 0.03
R221 fout2.n474 fout2.n473 0.03
R222 fout2.n183 fout2.n182 0.03
R223 fout2.n177 fout2.n176 0.03
R224 fout2.n301 fout2.n300 0.03
R225 fout2.n339 fout2.n338 0.03
R226 fout2.n368 fout2.n367 0.03
R227 fout2.n424 fout2.n423 0.03
R228 fout2.n491 fout2.n490 0.03
R229 fout2.n152 fout2.n151 0.028
R230 fout2.n150 fout2.n149 0.028
R231 fout2.n147 fout2.n146 0.028
R232 fout2.n145 fout2.n144 0.028
R233 fout2.n523 fout2.n522 0.028
R234 fout2.n521 fout2.n520 0.028
R235 fout2.n506 fout2.n505 0.028
R236 fout2.n508 fout2.n507 0.028
R237 fout2.n516 fout2.n515 0.028
R238 fout2.n531 fout2.n530 0.028
R239 fout2.n536 fout2.n535 0.028
R240 fout2.n501 fout2.n499 0.028
R241 fout2.n45 fout2.n44 0.028
R242 fout2.n43 fout2.n42 0.028
R243 fout2.n34 fout2.n33 0.028
R244 fout2.n36 fout2.n35 0.028
R245 fout2.n51 fout2.n50 0.028
R246 fout2.n17 fout2.n16 0.028
R247 fout2.n22 fout2.n21 0.028
R248 fout2.n28 fout2.n26 0.028
R249 fout2.n74 fout2.n73 0.028
R250 fout2.n72 fout2.n71 0.028
R251 fout2.n9 fout2.n8 0.028
R252 fout2.n11 fout2.n10 0.028
R253 fout2.n80 fout2.n79 0.028
R254 fout2.n61 fout2.n59 0.028
R255 fout2.n65 fout2.n64 0.028
R256 fout2.n3 fout2.n1 0.028
R257 fout2.n101 fout2.n100 0.028
R258 fout2.n90 fout2.n89 0.028
R259 fout2.n94 fout2.n93 0.028
R260 fout2.n117 fout2.n115 0.028
R261 fout2.n172 fout2.n169 0.028
R262 fout2.n210 fout2.n209 0.028
R263 fout2.n233 fout2.n232 0.028
R264 fout2.n248 fout2.n247 0.028
R265 fout2.n290 fout2.n249 0.028
R266 fout2.n279 fout2.n278 0.028
R267 fout2.n395 fout2.n387 0.028
R268 fout2.n439 fout2.n438 0.028
R269 fout2.n453 fout2.n452 0.028
R270 fout2.n476 fout2.n466 0.028
R271 fout2.n173 fout2.n165 0.028
R272 fout2.n200 fout2.n199 0.028
R273 fout2.n207 fout2.n206 0.028
R274 fout2.n291 fout2.n208 0.028
R275 fout2.n296 fout2.n295 0.028
R276 fout2.n306 fout2.n305 0.028
R277 fout2.n323 fout2.n322 0.028
R278 fout2.n336 fout2.n335 0.028
R279 fout2.n397 fout2.n396 0.028
R280 fout2.n416 fout2.n415 0.028
R281 fout2.n422 fout2.n421 0.028
R282 fout2.n487 fout2.n486 0.028
R283 fout2.n191 fout2.n190 0.027
R284 fout2.n194 fout2.n193 0.027
R285 fout2.n314 fout2.n313 0.027
R286 fout2.n317 fout2.n316 0.027
R287 fout2.n404 fout2.n403 0.027
R288 fout2.n407 fout2.n406 0.027
R289 fout2.n138 fout2.n137 0.026
R290 fout2.n136 fout2.n135 0.026
R291 fout2.n134 fout2.n133 0.026
R292 fout2.n132 fout2.n131 0.026
R293 fout2.n217 fout2.n215 0.026
R294 fout2.n270 fout2.n267 0.026
R295 fout2.n390 fout2.n389 0.026
R296 fout2.n437 fout2.n436 0.026
R297 fout2.n293 fout2.n292 0.026
R298 fout2.n307 fout2.n299 0.026
R299 fout2.n378 fout2.n377 0.026
R300 fout2.n414 fout2.n413 0.026
R301 fout2.n419 fout2.n418 0.026
R302 fout2.n489 fout2.n488 0.026
R303 fout2.n108 fout2.n107 0.025
R304 fout2.n106 fout2.n105 0.025
R305 fout2.n122 fout2.n121 0.025
R306 fout2.n124 fout2.n123 0.025
R307 fout2.n174 fout2.n173 0.024
R308 fout2.n277 fout2.n276 0.024
R309 fout2.n394 fout2.n391 0.024
R310 fout2.n164 fout2.n163 0.024
R311 fout2.n204 fout2.n203 0.024
R312 fout2.n299 fout2.n298 0.024
R313 fout2.n332 fout2.n331 0.024
R314 fout2.n375 fout2.n369 0.024
R315 fout2.n157 fout2.n156 0.023
R316 fout2.n241 fout2.n240 0.022
R317 fout2.n267 fout2.n266 0.022
R318 fout2.n355 fout2.n352 0.022
R319 fout2.n391 fout2.n390 0.022
R320 fout2.n446 fout2.n445 0.022
R321 fout2.n163 fout2.n162 0.022
R322 fout2.n307 fout2.n306 0.022
R323 fout2.n331 fout2.n330 0.022
R324 fout2.n396 fout2.n380 0.022
R325 fout2.n379 fout2.n378 0.022
R326 fout2.n284 fout2.n283 0.02
R327 fout2.n282 fout2.n279 0.02
R328 fout2.n278 fout2.n277 0.02
R329 fout2.n387 fout2.n386 0.02
R330 fout2.n371 fout2.n370 0.02
R331 fout2.n184 fout2.n183 0.02
R332 fout2.n297 fout2.n296 0.02
R333 fout2.n397 fout2.n368 0.02
R334 fout2.n490 fout2.n489 0.02
R335 fout2.n486 fout2.n480 0.02
R336 fout2.n185 fout2.n175 0.019
R337 fout2.n186 fout2.n185 0.019
R338 fout2.n308 fout2.n198 0.019
R339 fout2.n309 fout2.n308 0.019
R340 fout2.n398 fout2.n321 0.019
R341 fout2.n399 fout2.n398 0.019
R342 fout2.n492 fout2.n411 0.019
R343 fout2.n493 fout2.n492 0.019
R344 fout2.n455 fout2.n453 0.018
R345 fout2.n205 fout2.n204 0.018
R346 fout2.n491 fout2.n477 0.018
R347 fout2.n144 fout2.n143 0.017
R348 fout2.n142 fout2.n141 0.017
R349 fout2.n526 fout2.n525 0.017
R350 fout2.n516 fout2.n514 0.017
R351 fout2.n501 fout2.n500 0.017
R352 fout2.n510 fout2.n504 0.017
R353 fout2.n46 fout2.n41 0.017
R354 fout2.n51 fout2.n49 0.017
R355 fout2.n28 fout2.n27 0.017
R356 fout2.n38 fout2.n32 0.017
R357 fout2.n75 fout2.n70 0.017
R358 fout2.n80 fout2.n78 0.017
R359 fout2.n3 fout2.n2 0.017
R360 fout2.n13 fout2.n7 0.017
R361 fout2.n111 fout2.n110 0.017
R362 fout2.n101 fout2.n99 0.017
R363 fout2.n117 fout2.n116 0.017
R364 fout2.n126 fout2.n120 0.017
R365 fout2.n232 fout2.n231 0.017
R366 fout2.n260 fout2.n259 0.017
R367 fout2.n257 fout2.n256 0.017
R368 fout2.n484 fout2.n483 0.017
R369 fout2.n292 fout2.n291 0.017
R370 fout2.n295 fout2.n294 0.017
R371 fout2.n304 fout2.n303 0.017
R372 fout2.n302 fout2.n301 0.017
R373 fout2.n377 fout2.n376 0.017
R374 fout2.n418 fout2.n417 0.017
R375 fout2.n423 fout2.n422 0.017
R376 fout2.n480 fout2.n479 0.017
R377 fout2.n532 fout2.n529 0.016
R378 fout2.n537 fout2.n533 0.016
R379 fout2.n23 fout2.n19 0.016
R380 fout2.n66 fout2.n63 0.016
R381 fout2.n151 fout2.n150 0.015
R382 fout2.n146 fout2.n145 0.015
R383 fout2.n522 fout2.n521 0.015
R384 fout2.n507 fout2.n506 0.015
R385 fout2.n44 fout2.n43 0.015
R386 fout2.n35 fout2.n34 0.015
R387 fout2.n73 fout2.n72 0.015
R388 fout2.n10 fout2.n9 0.015
R389 fout2.n211 fout2.n210 0.015
R390 fout2.n221 fout2.n220 0.015
R391 fout2.n249 fout2.n248 0.015
R392 fout2.n359 fout2.n358 0.015
R393 fout2.n364 fout2.n361 0.015
R394 fout2.n438 fout2.n437 0.015
R395 fout2.n443 fout2.n439 0.015
R396 fout2.n475 fout2.n474 0.015
R397 fout2.n181 fout2.n180 0.015
R398 fout2.n179 fout2.n178 0.015
R399 fout2.n208 fout2.n207 0.015
R400 fout2.n338 fout2.n337 0.015
R401 fout2.n341 fout2.n340 0.015
R402 fout2.n366 fout2.n365 0.015
R403 fout2.n415 fout2.n414 0.015
R404 fout2.n417 fout2.n416 0.015
R405 fout2.n137 fout2.n136 0.013
R406 fout2.n133 fout2.n132 0.013
R407 fout2.n107 fout2.n106 0.013
R408 fout2.n123 fout2.n122 0.013
R409 fout2.n223 fout2.n222 0.013
R410 fout2.n247 fout2.n246 0.013
R411 fout2.n262 fout2.n260 0.013
R412 fout2.n460 fout2.n459 0.013
R413 fout2.n462 fout2.n461 0.013
R414 fout2.n206 fout2.n205 0.013
R415 fout2.n426 fout2.n425 0.013
R416 fout2.n428 fout2.n427 0.013
R417 fout2.n496 fout2.n495 0.013
R418 fout2.n538 fout2.n532 0.012
R419 fout2.n538 fout2.n537 0.012
R420 fout2.n24 fout2.n18 0.012
R421 fout2.n24 fout2.n23 0.012
R422 fout2.n67 fout2.n62 0.012
R423 fout2.n67 fout2.n66 0.012
R424 fout2.n96 fout2.n91 0.012
R425 fout2.n96 fout2.n95 0.012
R426 fout2.n192 fout2.n191 0.012
R427 fout2.n193 fout2.n192 0.012
R428 fout2.n315 fout2.n314 0.012
R429 fout2.n316 fout2.n315 0.012
R430 fout2.n405 fout2.n404 0.012
R431 fout2.n406 fout2.n405 0.012
R432 fout2.n519 fout2.n518 0.011
R433 fout2.n512 fout2.n503 0.011
R434 fout2.n54 fout2.n53 0.011
R435 fout2.n31 fout2.n30 0.011
R436 fout2.n83 fout2.n82 0.011
R437 fout2.n6 fout2.n5 0.011
R438 fout2.n104 fout2.n103 0.011
R439 fout2.n128 fout2.n119 0.011
R440 fout2.n285 fout2.n284 0.011
R441 fout2.n189 fout2.n188 0.011
R442 fout2.n196 fout2.n195 0.011
R443 fout2.n312 fout2.n311 0.011
R444 fout2.n319 fout2.n318 0.011
R445 fout2.n402 fout2.n401 0.011
R446 fout2.n409 fout2.n408 0.011
R447 fout2.n52 fout2.n48 0.01
R448 fout2.n81 fout2.n77 0.01
R449 fout2.n102 fout2.n98 0.01
R450 fout2.n118 fout2.n114 0.01
R451 fout2.n155 fout2.n154 0.01
R452 fout2.n156 fout2.n155 0.01
R453 fout2.n159 fout2.n158 0.009
R454 fout2.n169 fout2.n168 0.009
R455 fout2.n242 fout2.n241 0.009
R456 fout2.n246 fout2.n242 0.009
R457 fout2.n344 fout2.n343 0.009
R458 fout2.n445 fout2.n444 0.009
R459 fout2.n165 fout2.n164 0.009
R460 fout2.n330 fout2.n329 0.009
R461 fout2.n239 fout2.n235 0.007
R462 fout2.n327 fout2.n324 0.007
R463 fout2.n346 fout2.n345 0.007
R464 fout2.n352 fout2.n351 0.007
R465 fout2.n444 fout2.n443 0.007
R466 fout2.n472 fout2.n471 0.007
R467 fout2.n203 fout2.n202 0.007
R468 fout2.n328 fout2.n323 0.007
R469 fout2.n333 fout2.n332 0.007
R470 fout2.n335 fout2.n334 0.007
R471 fout2.n488 fout2.n487 0.007
R472 fout2.n479 fout2.n478 0.007
R473 fout2.n518 fout2.n517 0.006
R474 fout2.n503 fout2.n502 0.006
R475 fout2.n512 fout2.n511 0.006
R476 fout2.n54 fout2.n47 0.006
R477 fout2.n53 fout2.n52 0.006
R478 fout2.n30 fout2.n29 0.006
R479 fout2.n83 fout2.n76 0.006
R480 fout2.n82 fout2.n81 0.006
R481 fout2.n5 fout2.n4 0.006
R482 fout2.n103 fout2.n102 0.006
R483 fout2.n119 fout2.n118 0.006
R484 fout2.n128 fout2.n127 0.006
R485 fout2.n188 fout2.n187 0.006
R486 fout2.n190 fout2.n189 0.006
R487 fout2.n195 fout2.n194 0.006
R488 fout2.n197 fout2.n196 0.006
R489 fout2.n311 fout2.n310 0.006
R490 fout2.n313 fout2.n312 0.006
R491 fout2.n318 fout2.n317 0.006
R492 fout2.n320 fout2.n319 0.006
R493 fout2.n401 fout2.n400 0.006
R494 fout2.n403 fout2.n402 0.006
R495 fout2.n408 fout2.n407 0.006
R496 fout2.n410 fout2.n409 0.006
R497 fout2.n495 fout2.n494 0.006
R498 fout2.n158 fout2.n157 0.005
R499 fout2.n160 fout2.n159 0.005
R500 fout2.n215 fout2.n211 0.005
R501 fout2.n219 fout2.n217 0.005
R502 fout2.n290 fout2.n285 0.005
R503 fout2.n283 fout2.n282 0.005
R504 fout2.n255 fout2.n254 0.005
R505 fout2.n356 fout2.n355 0.005
R506 fout2.n431 fout2.n430 0.005
R507 fout2.n451 fout2.n450 0.005
R508 fout2.n376 fout2.n375 0.005
R509 fout2.n420 fout2.n419 0.005
R510 fout2.n97 fout2.n88 0.004
R511 fout2.n540 fout2.n539 0.004
R512 fout2.n25 fout2.n15 0.003
R513 fout2.n56 fout2.n55 0.003
R514 fout2.n68 fout2.n58 0.003
R515 fout2.n85 fout2.n84 0.003
R516 fout2.n130 fout2.n129 0.003
R517 fout2.n513 fout2.n498 0.003
R518 fout2.n172 fout2.n166 0.003
R519 fout2.n364 fout2.n360 0.003
R520 fout2.n385 fout2.n382 0.003
R521 fout2.n374 fout2.n371 0.003
R522 fout2.n450 fout2.n446 0.003
R523 fout2.n466 fout2.n464 0.003
R524 fout2.n476 fout2.n475 0.003
R525 fout2.n485 fout2.n484 0.003
R526 fout2.n294 fout2.n293 0.003
R527 fout2.n425 fout2.n424 0.003
R528 fout2.n527 fout2.n519 0.003
R529 fout2.n112 fout2.n104 0.003
R530 fout2.n14 fout2.n6 0.003
R531 fout2.n39 fout2.n31 0.003
R532 fout2.n113 fout2.n97 0.002
R533 fout2.n539 fout2.n528 0.002
R534 fout2.n129 fout2.n113 0.002
R535 fout2.n84 fout2.n69 0.002
R536 fout2.n55 fout2.n40 0.002
R537 fout2.n69 fout2.n68 0.002
R538 fout2.n40 fout2.n25 0.002
R539 fout2.n528 fout2.n513 0.002
R540 fout2.n227 fout2.n223 0.001
R541 fout2.n231 fout2.n229 0.001
R542 fout2.n234 fout2.n233 0.001
R543 fout2.n240 fout2.n239 0.001
R544 fout2.n276 fout2.n273 0.001
R545 fout2.n271 fout2.n270 0.001
R546 fout2.n265 fout2.n262 0.001
R547 fout2.n259 fout2.n258 0.001
R548 fout2.n351 fout2.n347 0.001
R549 fout2.n357 fout2.n356 0.001
R550 fout2.n436 fout2.n431 0.001
R551 fout2.n178 fout2.n177 0.001
R552 fout2.n201 fout2.n200 0.001
R553 fout2.n337 fout2.n336 0.001
R554 fout2.n340 fout2.n339 0.001
R555 fout2.n413 fout2.n412 0.001
R556 fout2.n87 fout2.n0 0.001
R557 GND.t91 GND.n1080 73112.5
R558 GND.t70 GND.t96 3181.77
R559 GND.t93 GND.t29 3178.99
R560 GND.t103 GND.t72 3178.99
R561 GND.t142 GND.t68 3169.21
R562 GND.t88 GND.t20 3007.96
R563 GND.t29 GND.t128 3007.96
R564 GND.t78 GND.t106 3007.96
R565 GND.t96 GND.t43 3007.96
R566 GND.t115 GND.t6 3007.96
R567 GND.t68 GND.t19 3007.96
R568 GND.t87 GND.t80 3007.96
R569 GND.t72 GND.t102 3007.96
R570 GND.n29 GND.t88 2521.24
R571 GND.n965 GND.t115 2521.24
R572 GND.n620 GND.t78 2511.5
R573 GND.n1080 GND.t87 2511.5
R574 GND.t124 GND.t142 2199.81
R575 GND.t22 GND.t70 2197.82
R576 GND.t84 GND.t93 2189.94
R577 GND.t47 GND.t103 2189.94
R578 GND.n1237 GND.n1236 1893.67
R579 GND.n543 GND.n420 1881.76
R580 GND.n888 GND.n765 1881.76
R581 GND.n1163 GND.n1145 1475.95
R582 GND.n1175 GND.n1174 1475.95
R583 GND.n1185 GND.n1184 1475.95
R584 GND.n1196 GND.n1131 1475.95
R585 GND.n1198 GND.n1124 1475.95
R586 GND.n1210 GND.n1209 1475.95
R587 GND.n1222 GND.n1221 1475.95
R588 GND.n1236 GND.n1110 1475.95
R589 GND.n1238 GND.n1237 1475.95
R590 GND.n1248 GND.n1247 1475.95
R591 GND.n1261 GND.n1096 1475.95
R592 GND.n481 GND.n480 1466.67
R593 GND.n492 GND.n455 1466.67
R594 GND.n494 GND.n448 1466.67
R595 GND.n506 GND.n505 1466.67
R596 GND.n516 GND.n515 1466.67
R597 GND.n527 GND.n434 1466.67
R598 GND.n529 GND.n426 1466.67
R599 GND.n543 GND.n542 1466.67
R600 GND.n554 GND.n420 1466.67
R601 GND.n556 GND.n414 1466.67
R602 GND.n570 GND.n569 1466.67
R603 GND.n826 GND.n825 1466.67
R604 GND.n837 GND.n800 1466.67
R605 GND.n839 GND.n793 1466.67
R606 GND.n851 GND.n850 1466.67
R607 GND.n861 GND.n860 1466.67
R608 GND.n872 GND.n779 1466.67
R609 GND.n874 GND.n771 1466.67
R610 GND.n888 GND.n887 1466.67
R611 GND.n899 GND.n765 1466.67
R612 GND.n901 GND.n759 1466.67
R613 GND.n915 GND.n914 1466.67
R614 GND.n1410 GND.n1399 1008.92
R615 GND.n1897 GND.n1892 1002.53
R616 GND.n1648 GND.n1643 1002.53
R617 GND.n1161 GND.n1152 1002.53
R618 GND.n473 GND.n468 996.226
R619 GND.n818 GND.n813 996.226
R620 GND.t79 GND.t84 917.985
R621 GND.t57 GND.t22 917.985
R622 GND.t101 GND.t124 917.985
R623 GND.t54 GND.t47 917.985
R624 GND.n2067 GND.t135 886.33
R625 GND.n1818 GND.t111 886.33
R626 GND.n2104 GND.t155 882.813
R627 GND.n1377 GND.t86 882.813
R628 GND.t133 GND.t79 854.676
R629 GND.t145 GND.t54 854.676
R630 GND.t2 GND.t57 851.159
R631 GND.t4 GND.t101 851.159
R632 GND.n620 GND.n391 760.672
R633 GND.n965 GND.n736 760.672
R634 GND.n29 GND.n26 760.624
R635 GND.n1300 GND.n1084 759.292
R636 GND.t98 GND.t133 703.437
R637 GND.t42 GND.t2 703.437
R638 GND.t144 GND.t4 703.437
R639 GND.t105 GND.t145 703.437
R640 GND.t155 GND.t98 703.436
R641 GND.t135 GND.t42 703.436
R642 GND.t111 GND.t144 703.436
R643 GND.t86 GND.t105 703.436
R644 GND.n472 GND.n471 585
R645 GND.n473 GND.n472 585
R646 GND.n463 GND.n462 585
R647 GND.n462 GND.n461 585
R648 GND.n484 GND.n483 585
R649 GND.n483 GND.n482 585
R650 GND.n454 GND.n452 585
R651 GND.n493 GND.n454 585
R652 GND.n503 GND.n502 585
R653 GND.n504 GND.n503 585
R654 GND.n442 GND.n441 585
R655 GND.n441 GND.n440 585
R656 GND.n519 GND.n518 585
R657 GND.n518 GND.n517 585
R658 GND.n433 GND.n431 585
R659 GND.n528 GND.n433 585
R660 GND.n540 GND.n539 585
R661 GND.n541 GND.n540 585
R662 GND.n419 GND.n418 585
R663 GND.n555 GND.n419 585
R664 GND.n567 GND.n566 585
R665 GND.n568 GND.n567 585
R666 GND.n409 GND.n407 585
R667 GND.n407 GND.n406 585
R668 GND.n611 GND.n610 585
R669 GND.n579 GND.n578 585
R670 GND.n583 GND.n581 585
R671 GND.n591 GND.n586 585
R672 GND.n390 GND.n388 585
R673 GND.n402 GND.n399 585
R674 GND.n401 GND.n400 585
R675 GND.n587 GND.n389 585
R676 GND.n585 GND.n584 585
R677 GND.n598 GND.n580 585
R678 GND.n609 GND.n608 585
R679 GND.n618 GND.n617 585
R680 GND.n619 GND.n618 585
R681 GND.n565 GND.n413 585
R682 GND.n569 GND.n413 585
R683 GND.n558 GND.n557 585
R684 GND.n557 GND.n556 585
R685 GND.n470 GND.n469 585
R686 GND.n469 GND.n468 585
R687 GND.n460 GND.n459 585
R688 GND.n481 GND.n460 585
R689 GND.n491 GND.n490 585
R690 GND.n492 GND.n491 585
R691 GND.n450 GND.n449 585
R692 GND.n449 GND.n448 585
R693 GND.n508 GND.n507 585
R694 GND.n507 GND.n506 585
R695 GND.n439 GND.n438 585
R696 GND.n516 GND.n439 585
R697 GND.n526 GND.n525 585
R698 GND.n527 GND.n526 585
R699 GND.n428 GND.n427 585
R700 GND.n427 GND.n426 585
R701 GND.n404 GND.n403 585
R702 GND.n467 GND.n466 585
R703 GND.n1896 GND.n1895 585
R704 GND.n1897 GND.n1896 585
R705 GND.n1888 GND.n1886 585
R706 GND.n1886 GND.n1885 585
R707 GND.n2058 GND.n2057 585
R708 GND.n1906 GND.n1905 585
R709 GND.n2046 GND.n2045 585
R710 GND.n2036 GND.n2035 585
R711 GND.n2030 GND.n2029 585
R712 GND.n2020 GND.n2019 585
R713 GND.n2014 GND.n2013 585
R714 GND.n1996 GND.n1995 585
R715 GND.n1932 GND.n1929 585
R716 GND.n1984 GND.n1935 585
R717 GND.n1940 GND.n1938 585
R718 GND.n1970 GND.n1943 585
R719 GND.n1948 GND.n1946 585
R720 GND.n1956 GND.n1951 585
R721 GND.n1854 GND.n1852 585
R722 GND.n1880 GND.n1877 585
R723 GND.n1879 GND.n1878 585
R724 GND.n1952 GND.n1853 585
R725 GND.n1950 GND.n1949 585
R726 GND.n1963 GND.n1945 585
R727 GND.n1942 GND.n1941 585
R728 GND.n1977 GND.n1937 585
R729 GND.n1934 GND.n1933 585
R730 GND.n1994 GND.n1993 585
R731 GND.n1894 GND.n1893 585
R732 GND.n1893 GND.n1892 585
R733 GND.n2059 GND.n1887 585
R734 GND.n1904 GND.n1903 585
R735 GND.n2048 GND.n2047 585
R736 GND.n2038 GND.n2037 585
R737 GND.n2032 GND.n2031 585
R738 GND.n2022 GND.n2021 585
R739 GND.n2016 GND.n2015 585
R740 GND.n1882 GND.n1881 585
R741 GND.n1891 GND.n1890 585
R742 GND.n817 GND.n816 585
R743 GND.n818 GND.n817 585
R744 GND.n808 GND.n807 585
R745 GND.n807 GND.n806 585
R746 GND.n829 GND.n828 585
R747 GND.n828 GND.n827 585
R748 GND.n799 GND.n797 585
R749 GND.n838 GND.n799 585
R750 GND.n848 GND.n847 585
R751 GND.n849 GND.n848 585
R752 GND.n787 GND.n786 585
R753 GND.n786 GND.n785 585
R754 GND.n864 GND.n863 585
R755 GND.n863 GND.n862 585
R756 GND.n778 GND.n776 585
R757 GND.n873 GND.n778 585
R758 GND.n885 GND.n884 585
R759 GND.n886 GND.n885 585
R760 GND.n764 GND.n763 585
R761 GND.n900 GND.n764 585
R762 GND.n912 GND.n911 585
R763 GND.n913 GND.n912 585
R764 GND.n754 GND.n752 585
R765 GND.n752 GND.n751 585
R766 GND.n956 GND.n955 585
R767 GND.n924 GND.n923 585
R768 GND.n928 GND.n926 585
R769 GND.n936 GND.n931 585
R770 GND.n735 GND.n733 585
R771 GND.n747 GND.n744 585
R772 GND.n746 GND.n745 585
R773 GND.n932 GND.n734 585
R774 GND.n930 GND.n929 585
R775 GND.n943 GND.n925 585
R776 GND.n954 GND.n953 585
R777 GND.n963 GND.n962 585
R778 GND.n964 GND.n963 585
R779 GND.n910 GND.n758 585
R780 GND.n914 GND.n758 585
R781 GND.n903 GND.n902 585
R782 GND.n902 GND.n901 585
R783 GND.n815 GND.n814 585
R784 GND.n814 GND.n813 585
R785 GND.n805 GND.n804 585
R786 GND.n826 GND.n805 585
R787 GND.n836 GND.n835 585
R788 GND.n837 GND.n836 585
R789 GND.n795 GND.n794 585
R790 GND.n794 GND.n793 585
R791 GND.n853 GND.n852 585
R792 GND.n852 GND.n851 585
R793 GND.n784 GND.n783 585
R794 GND.n861 GND.n784 585
R795 GND.n871 GND.n870 585
R796 GND.n872 GND.n871 585
R797 GND.n773 GND.n772 585
R798 GND.n772 GND.n771 585
R799 GND.n749 GND.n748 585
R800 GND.n812 GND.n811 585
R801 GND.n1647 GND.n1646 585
R802 GND.n1648 GND.n1647 585
R803 GND.n1639 GND.n1637 585
R804 GND.n1637 GND.n1636 585
R805 GND.n1809 GND.n1808 585
R806 GND.n1657 GND.n1656 585
R807 GND.n1797 GND.n1796 585
R808 GND.n1787 GND.n1786 585
R809 GND.n1781 GND.n1780 585
R810 GND.n1771 GND.n1770 585
R811 GND.n1765 GND.n1764 585
R812 GND.n1747 GND.n1746 585
R813 GND.n1683 GND.n1680 585
R814 GND.n1735 GND.n1686 585
R815 GND.n1691 GND.n1689 585
R816 GND.n1721 GND.n1694 585
R817 GND.n1699 GND.n1697 585
R818 GND.n1707 GND.n1702 585
R819 GND.n1605 GND.n1603 585
R820 GND.n1631 GND.n1628 585
R821 GND.n1630 GND.n1629 585
R822 GND.n1703 GND.n1604 585
R823 GND.n1701 GND.n1700 585
R824 GND.n1714 GND.n1696 585
R825 GND.n1693 GND.n1692 585
R826 GND.n1728 GND.n1688 585
R827 GND.n1685 GND.n1684 585
R828 GND.n1745 GND.n1744 585
R829 GND.n1645 GND.n1644 585
R830 GND.n1644 GND.n1643 585
R831 GND.n1810 GND.n1638 585
R832 GND.n1655 GND.n1654 585
R833 GND.n1799 GND.n1798 585
R834 GND.n1789 GND.n1788 585
R835 GND.n1783 GND.n1782 585
R836 GND.n1773 GND.n1772 585
R837 GND.n1767 GND.n1766 585
R838 GND.n1633 GND.n1632 585
R839 GND.n1642 GND.n1641 585
R840 GND.n1158 GND.n1153 585
R841 GND.n1153 GND.n1152 585
R842 GND.n1151 GND.n1149 585
R843 GND.n1162 GND.n1151 585
R844 GND.n1172 GND.n1171 585
R845 GND.n1173 GND.n1172 585
R846 GND.n1139 GND.n1138 585
R847 GND.n1138 GND.n1137 585
R848 GND.n1188 GND.n1187 585
R849 GND.n1187 GND.n1186 585
R850 GND.n1130 GND.n1128 585
R851 GND.n1197 GND.n1130 585
R852 GND.n1207 GND.n1206 585
R853 GND.n1208 GND.n1207 585
R854 GND.n1119 GND.n1118 585
R855 GND.n1118 GND.n1117 585
R856 GND.n1225 GND.n1224 585
R857 GND.n1224 GND.n1223 585
R858 GND.n1105 GND.n1104 585
R859 GND.n1104 GND.n1103 585
R860 GND.n1251 GND.n1250 585
R861 GND.n1250 GND.n1249 585
R862 GND.n1099 GND.n1094 585
R863 GND.n1262 GND.n1094 585
R864 GND.n1090 GND.n1088 585
R865 GND.n1292 GND.n1291 585
R866 GND.n1273 GND.n1272 585
R867 GND.n1276 GND.n1275 585
R868 GND.n1309 GND.n1078 585
R869 GND.n1306 GND.n1305 585
R870 GND.n1308 GND.n1301 585
R871 GND.n1277 GND.n1079 585
R872 GND.n1300 GND.n1079 585
R873 GND.n1274 GND.n1086 585
R874 GND.n1300 GND.n1086 585
R875 GND.n1290 GND.n1082 585
R876 GND.n1300 GND.n1082 585
R877 GND.n1299 GND.n1298 585
R878 GND.n1300 GND.n1299 585
R879 GND.n1264 GND.n1095 585
R880 GND.n1264 GND.n1263 585
R881 GND.n1252 GND.n1097 585
R882 GND.n1097 GND.n1096 585
R883 GND.n1246 GND.n1245 585
R884 GND.n1247 GND.n1246 585
R885 GND.n1160 GND.n1159 585
R886 GND.n1161 GND.n1160 585
R887 GND.n1147 GND.n1146 585
R888 GND.n1146 GND.n1145 585
R889 GND.n1177 GND.n1176 585
R890 GND.n1176 GND.n1175 585
R891 GND.n1136 GND.n1135 585
R892 GND.n1185 GND.n1136 585
R893 GND.n1195 GND.n1194 585
R894 GND.n1196 GND.n1195 585
R895 GND.n1126 GND.n1125 585
R896 GND.n1125 GND.n1124 585
R897 GND.n1212 GND.n1211 585
R898 GND.n1211 GND.n1210 585
R899 GND.n1116 GND.n1115 585
R900 GND.n1222 GND.n1116 585
R901 GND.n1304 GND.n1303 585
R902 GND.n1157 GND.n1156 585
R903 GND.n1406 GND.n1400 585
R904 GND.n1400 GND.n1399 585
R905 GND.n1407 GND.n1397 585
R906 GND.n1411 GND.n1397 585
R907 GND.n1393 GND.n1391 585
R908 GND.n1553 GND.n1552 585
R909 GND.n1424 GND.n1423 585
R910 GND.n1429 GND.n1428 585
R911 GND.n1434 GND.n1433 585
R912 GND.n1439 GND.n1438 585
R913 GND.n1444 GND.n1443 585
R914 GND.n1451 GND.n1450 585
R915 GND.n1456 GND.n1455 585
R916 GND.n1460 GND.n1459 585
R917 GND.n1464 GND.n1463 585
R918 GND.n1468 GND.n1467 585
R919 GND.n1472 GND.n1471 585
R920 GND.n1476 GND.n1475 585
R921 GND.n1570 GND.n1361 585
R922 GND.n1567 GND.n1566 585
R923 GND.n1569 GND.n1562 585
R924 GND.n1477 GND.n1362 585
R925 GND.n1561 GND.n1362 585
R926 GND.n1474 GND.n1379 585
R927 GND.n1561 GND.n1379 585
R928 GND.n1470 GND.n1375 585
R929 GND.n1561 GND.n1375 585
R930 GND.n1466 GND.n1381 585
R931 GND.n1561 GND.n1381 585
R932 GND.n1462 GND.n1373 585
R933 GND.n1561 GND.n1373 585
R934 GND.n1458 GND.n1383 585
R935 GND.n1561 GND.n1383 585
R936 GND.n1454 GND.n1371 585
R937 GND.n1561 GND.n1371 585
R938 GND.n1409 GND.n1408 585
R939 GND.n1410 GND.n1409 585
R940 GND.n1415 GND.n1414 585
R941 GND.n1554 GND.n1392 585
R942 GND.n1422 GND.n1421 585
R943 GND.n1426 GND.n1425 585
R944 GND.n1431 GND.n1430 585
R945 GND.n1436 GND.n1435 585
R946 GND.n1441 GND.n1440 585
R947 GND.n1565 GND.n1564 585
R948 GND.n1405 GND.n1404 585
R949 GND.n2113 GND.n2112 483.388
R950 GND.n1403 GND.n1399 483.388
R951 GND.n1898 GND.n1897 480.395
R952 GND.n1649 GND.n1648 480.395
R953 GND.n1155 GND.n1152 480.395
R954 GND.n38 GND.n37 477.439
R955 GND.n474 GND.n473 477.439
R956 GND.n819 GND.n818 477.439
R957 GND.n2119 GND.n2118 448.407
R958 GND.n1411 GND.n1410 448.407
R959 GND.n1892 GND.n1885 445.569
R960 GND.n1643 GND.n1636 445.569
R961 GND.n1162 GND.n1161 445.569
R962 GND.n44 GND.n43 442.767
R963 GND.n468 GND.n461 442.767
R964 GND.n813 GND.n806 442.767
R965 GND.n1223 GND.n1110 417.721
R966 GND.n1238 GND.n1103 417.721
R967 GND.n145 GND.n144 415.094
R968 GND.n169 GND.n168 415.094
R969 GND.n542 GND.n541 415.094
R970 GND.n555 GND.n554 415.094
R971 GND.n887 GND.n886 415.094
R972 GND.n900 GND.n899 415.094
R973 GND.n1173 GND.n1145 389.873
R974 GND.n58 GND.n57 387.421
R975 GND.n482 GND.n481 387.421
R976 GND.n827 GND.n826 387.421
R977 GND.n1221 GND.n1117 362.025
R978 GND.n1249 GND.n1248 362.025
R979 GND.n129 GND.n128 359.748
R980 GND.n183 GND.n182 359.748
R981 GND.n529 GND.n528 359.748
R982 GND.n568 GND.n414 359.748
R983 GND.n874 GND.n873 359.748
R984 GND.n913 GND.n759 359.748
R985 GND.n1175 GND.n1137 334.177
R986 GND.n72 GND.n71 332.075
R987 GND.n493 GND.n492 332.075
R988 GND.n838 GND.n837 332.075
R989 GND.n1209 GND.n1208 306.329
R990 GND.n1262 GND.n1261 306.329
R991 GND.n115 GND.n114 304.402
R992 GND.n517 GND.n434 304.402
R993 GND.n570 GND.n406 304.402
R994 GND.n862 GND.n779 304.402
R995 GND.n915 GND.n751 304.402
R996 GND.n142 GND.n141 292.5
R997 GND.n164 GND.n163 292.5
R998 GND.n547 GND.n421 292.5
R999 GND.n421 GND.n420 292.5
R1000 GND.n545 GND.n544 292.5
R1001 GND.n544 GND.n543 292.5
R1002 GND.n2004 GND.n2003 292.5
R1003 GND.n2006 GND.n2005 292.5
R1004 GND.n892 GND.n766 292.5
R1005 GND.n766 GND.n765 292.5
R1006 GND.n890 GND.n889 292.5
R1007 GND.n889 GND.n888 292.5
R1008 GND.n1755 GND.n1754 292.5
R1009 GND.n1757 GND.n1756 292.5
R1010 GND.n1113 GND.n1109 292.5
R1011 GND.n1237 GND.n1109 292.5
R1012 GND.n1235 GND.n1234 292.5
R1013 GND.n1236 GND.n1235 292.5
R1014 GND.n1520 GND.n1519 292.5
R1015 GND.n1446 GND.n1445 292.5
R1016 GND.n2067 GND.n1866 291.574
R1017 GND.n2067 GND.n1864 291.574
R1018 GND.n1818 GND.n1617 291.574
R1019 GND.n1818 GND.n1615 291.574
R1020 GND.n1561 GND.n1369 291.565
R1021 GND.n1561 GND.n1386 290.636
R1022 GND.n2067 GND.n1869 289.739
R1023 GND.n2067 GND.n1861 289.739
R1024 GND.n1818 GND.n1620 289.739
R1025 GND.n1818 GND.n1612 289.739
R1026 GND.n1561 GND.n1367 289.713
R1027 GND.n1561 GND.n1388 288.796
R1028 GND.n620 GND.n394 287.969
R1029 GND.n965 GND.n739 287.969
R1030 GND.n2067 GND.n1872 287.927
R1031 GND.n2067 GND.n1858 287.927
R1032 GND.n1818 GND.n1623 287.927
R1033 GND.n1818 GND.n1609 287.927
R1034 GND.n1561 GND.n1365 287.884
R1035 GND.n1561 GND.n1390 286.978
R1036 GND.n620 GND.n397 286.196
R1037 GND.n965 GND.n742 286.196
R1038 GND.n2067 GND.n1875 286.138
R1039 GND.n2067 GND.n1855 286.138
R1040 GND.n1818 GND.n1626 286.138
R1041 GND.n1818 GND.n1606 286.138
R1042 GND.n1561 GND.n1363 286.078
R1043 GND.n1186 GND.n1185 278.481
R1044 GND.n620 GND.n398 276.819
R1045 GND.n965 GND.n743 276.819
R1046 GND.n86 GND.n85 276.729
R1047 GND.n504 GND.n448 276.729
R1048 GND.n849 GND.n793 276.729
R1049 GND.n2067 GND.n1876 276.679
R1050 GND.n1818 GND.n1627 276.679
R1051 GND.n1307 GND.n1300 276.679
R1052 GND.n1568 GND.n1561 276.537
R1053 GND.n2067 GND.n2066 250.632
R1054 GND.n1198 GND.n1197 250.632
R1055 GND.n101 GND.n100 249.056
R1056 GND.n515 GND.n440 249.056
R1057 GND.n860 GND.n785 249.056
R1058 GND.n1412 GND.n1377 224.203
R1059 GND.n1818 GND.n1817 222.784
R1060 GND.n1197 GND.n1196 222.784
R1061 GND.n100 GND.n99 221.383
R1062 GND.n506 GND.n440 221.383
R1063 GND.n851 GND.n785 221.383
R1064 GND.n1186 GND.n1131 194.936
R1065 GND.n87 GND.n86 193.71
R1066 GND.n505 GND.n504 193.71
R1067 GND.n850 GND.n849 193.71
R1068 GND.n368 GND.n367 185
R1069 GND.n382 GND.n381 185
R1070 GND.n348 GND.n347 185
R1071 GND.n362 GND.n361 185
R1072 GND.n630 GND.n629 185
R1073 GND.n644 GND.n643 185
R1074 GND.n650 GND.n649 185
R1075 GND.n664 GND.n663 185
R1076 GND.n672 GND.n671 185
R1077 GND.n686 GND.n685 185
R1078 GND.n713 GND.n712 185
R1079 GND.n727 GND.n726 185
R1080 GND.n693 GND.n692 185
R1081 GND.n707 GND.n706 185
R1082 GND.n975 GND.n974 185
R1083 GND.n989 GND.n988 185
R1084 GND.n995 GND.n994 185
R1085 GND.n1009 GND.n1008 185
R1086 GND.n1017 GND.n1016 185
R1087 GND.n1031 GND.n1030 185
R1088 GND.n1058 GND.n1057 185
R1089 GND.n1072 GND.n1071 185
R1090 GND.n1038 GND.n1037 185
R1091 GND.n1052 GND.n1051 185
R1092 GND.n1319 GND.n1318 185
R1093 GND.n1333 GND.n1332 185
R1094 GND.n1339 GND.n1338 185
R1095 GND.n1353 GND.n1352 185
R1096 GND.n1580 GND.n1579 185
R1097 GND.n1594 GND.n1593 185
R1098 GND.n1829 GND.n1828 185
R1099 GND.n1843 GND.n1842 185
R1100 GND.n2078 GND.n2077 185
R1101 GND.n2092 GND.n2091 185
R1102 GND.n1208 GND.n1124 167.088
R1103 GND.n1263 GND.n1262 167.088
R1104 GND.n114 GND.n113 166.037
R1105 GND.n28 GND.n27 166.037
R1106 GND.n517 GND.n516 166.037
R1107 GND.n619 GND.n406 166.037
R1108 GND.n862 GND.n861 166.037
R1109 GND.n964 GND.n751 166.037
R1110 GND.n1184 GND.n1137 139.24
R1111 GND.n73 GND.n72 138.364
R1112 GND.n494 GND.n493 138.364
R1113 GND.n839 GND.n838 138.364
R1114 GND.n2005 GND.n2004 126.377
R1115 GND.n1756 GND.n1755 126.377
R1116 GND.n1235 GND.n1109 126.377
R1117 GND.n544 GND.n421 125.196
R1118 GND.n889 GND.n766 125.196
R1119 GND.n264 GND.t28 124.695
R1120 GND.n284 GND.t94 124.695
R1121 GND.n304 GND.t30 124.695
R1122 GND.n326 GND.t44 124.695
R1123 GND.n351 GND.t154 124.695
R1124 GND.n633 GND.t71 124.695
R1125 GND.n653 GND.t97 124.695
R1126 GND.n675 GND.t120 124.695
R1127 GND.n696 GND.t49 124.695
R1128 GND.n978 GND.t143 124.695
R1129 GND.n998 GND.t69 124.695
R1130 GND.n1020 GND.t40 124.695
R1131 GND.n1041 GND.t41 124.695
R1132 GND.n1322 GND.t104 124.695
R1133 GND.n1342 GND.t73 124.695
R1134 GND.n2348 GND.t110 124.695
R1135 GND.n1583 GND.t81 124.695
R1136 GND.n1832 GND.t7 124.695
R1137 GND.n2081 GND.t107 124.695
R1138 GND.n2326 GND.t21 124.695
R1139 GND.n2 GND.t46 124.688
R1140 GND.n716 GND.t51 124.688
R1141 GND.n1061 GND.t92 124.688
R1142 GND.n371 GND.t148 124.686
R1143 GND.n1561 GND.n1370 120.066
R1144 GND.n383 GND.n382 118.319
R1145 GND.n363 GND.n362 118.319
R1146 GND.n645 GND.n644 118.319
R1147 GND.n665 GND.n664 118.319
R1148 GND.n687 GND.n686 118.319
R1149 GND.n728 GND.n727 118.319
R1150 GND.n708 GND.n707 118.319
R1151 GND.n990 GND.n989 118.319
R1152 GND.n1010 GND.n1009 118.319
R1153 GND.n1032 GND.n1031 118.319
R1154 GND.n1073 GND.n1072 118.319
R1155 GND.n1053 GND.n1052 118.319
R1156 GND.n1334 GND.n1333 118.319
R1157 GND.n1354 GND.n1353 118.319
R1158 GND.n1595 GND.n1594 118.319
R1159 GND.n1844 GND.n1843 118.319
R1160 GND.n2093 GND.n2092 118.319
R1161 GND.n1210 GND.n1117 111.392
R1162 GND.n1249 GND.n1096 111.392
R1163 GND.n128 GND.n127 110.691
R1164 GND.n182 GND.n181 110.691
R1165 GND.n528 GND.n527 110.691
R1166 GND.n569 GND.n568 110.691
R1167 GND.n873 GND.n872 110.691
R1168 GND.n914 GND.n913 110.691
R1169 GND.n376 GND.n375 109.655
R1170 GND.n356 GND.n355 109.655
R1171 GND.n638 GND.n637 109.655
R1172 GND.n658 GND.n657 109.655
R1173 GND.n680 GND.n679 109.655
R1174 GND.n721 GND.n720 109.655
R1175 GND.n701 GND.n700 109.655
R1176 GND.n983 GND.n982 109.655
R1177 GND.n1003 GND.n1002 109.655
R1178 GND.n1025 GND.n1024 109.655
R1179 GND.n1066 GND.n1065 109.655
R1180 GND.n1046 GND.n1045 109.655
R1181 GND.n1327 GND.n1326 109.655
R1182 GND.n1347 GND.n1346 109.655
R1183 GND.n1588 GND.n1587 109.655
R1184 GND.n1837 GND.n1836 109.655
R1185 GND.n2086 GND.n2085 109.655
R1186 GND.n1414 GND.n1413 99.438
R1187 GND.n1560 GND.n1392 99.438
R1188 GND.n1421 GND.n1364 99.438
R1189 GND.n1425 GND.n1389 99.438
R1190 GND.n1430 GND.n1366 99.438
R1191 GND.n1435 GND.n1387 99.438
R1192 GND.n1440 GND.n1368 99.438
R1193 GND.n1445 GND.n1385 99.438
R1194 GND.n1519 GND.n1518 99.438
R1195 GND.n1511 GND.n1371 99.438
R1196 GND.n1505 GND.n1383 99.438
R1197 GND.n1499 GND.n1373 99.438
R1198 GND.n1493 GND.n1381 99.438
R1199 GND.n1487 GND.n1375 99.438
R1200 GND.n1481 GND.n1379 99.438
R1201 GND.n1572 GND.n1362 99.438
R1202 GND.n2065 GND.n1887 98.5
R1203 GND.n2049 GND.n2048 98.5
R1204 GND.n2033 GND.n2032 98.5
R1205 GND.n2017 GND.n2016 98.5
R1206 GND.n1993 GND.n1992 98.5
R1207 GND.n1978 GND.n1977 98.5
R1208 GND.n1964 GND.n1963 98.5
R1209 GND.n2069 GND.n1853 98.5
R1210 GND.n1816 GND.n1638 98.5
R1211 GND.n1800 GND.n1799 98.5
R1212 GND.n1784 GND.n1783 98.5
R1213 GND.n1768 GND.n1767 98.5
R1214 GND.n1744 GND.n1743 98.5
R1215 GND.n1729 GND.n1728 98.5
R1216 GND.n1715 GND.n1714 98.5
R1217 GND.n1820 GND.n1604 98.5
R1218 GND.n1164 GND.n1146 98.5
R1219 GND.n1176 GND.n1144 98.5
R1220 GND.n1183 GND.n1136 98.5
R1221 GND.n1195 GND.n1132 98.5
R1222 GND.n1199 GND.n1125 98.5
R1223 GND.n1211 GND.n1123 98.5
R1224 GND.n1220 GND.n1116 98.5
R1225 GND.n1235 GND.n1111 98.5
R1226 GND.n1239 GND.n1109 98.5
R1227 GND.n1246 GND.n1102 98.5
R1228 GND.n1260 GND.n1097 98.5
R1229 GND.n1265 GND.n1264 98.5
R1230 GND.n1299 GND.n1089 98.5
R1231 GND.n1269 GND.n1082 98.5
R1232 GND.n1281 GND.n1086 98.5
R1233 GND.n1311 GND.n1079 98.5
R1234 GND.n146 GND.n142 97.579
R1235 GND.n170 GND.n164 97.579
R1236 GND.n479 GND.n460 97.579
R1237 GND.n491 GND.n456 97.579
R1238 GND.n495 GND.n449 97.579
R1239 GND.n507 GND.n447 97.579
R1240 GND.n514 GND.n439 97.579
R1241 GND.n526 GND.n435 97.579
R1242 GND.n530 GND.n427 97.579
R1243 GND.n544 GND.n425 97.579
R1244 GND.n553 GND.n421 97.579
R1245 GND.n557 GND.n415 97.579
R1246 GND.n571 GND.n413 97.579
R1247 GND.n618 GND.n408 97.579
R1248 GND.n599 GND.n598 97.579
R1249 GND.n622 GND.n389 97.579
R1250 GND.n824 GND.n805 97.579
R1251 GND.n836 GND.n801 97.579
R1252 GND.n840 GND.n794 97.579
R1253 GND.n852 GND.n792 97.579
R1254 GND.n859 GND.n784 97.579
R1255 GND.n871 GND.n780 97.579
R1256 GND.n875 GND.n772 97.579
R1257 GND.n889 GND.n770 97.579
R1258 GND.n898 GND.n766 97.579
R1259 GND.n902 GND.n760 97.579
R1260 GND.n916 GND.n758 97.579
R1261 GND.n963 GND.n753 97.579
R1262 GND.n944 GND.n943 97.579
R1263 GND.n967 GND.n734 97.579
R1264 GND.n1 GND.n0 92.5
R1265 GND.n263 GND.n262 92.5
R1266 GND.n283 GND.n282 92.5
R1267 GND.n303 GND.n302 92.5
R1268 GND.n325 GND.n324 92.5
R1269 GND.n375 GND.n374 92.5
R1270 GND.n355 GND.n354 92.5
R1271 GND.n637 GND.n636 92.5
R1272 GND.n657 GND.n656 92.5
R1273 GND.n679 GND.n678 92.5
R1274 GND.n720 GND.n719 92.5
R1275 GND.n700 GND.n699 92.5
R1276 GND.n982 GND.n981 92.5
R1277 GND.n1002 GND.n1001 92.5
R1278 GND.n1024 GND.n1023 92.5
R1279 GND.n1065 GND.n1064 92.5
R1280 GND.n1045 GND.n1044 92.5
R1281 GND.n1326 GND.n1325 92.5
R1282 GND.n1346 GND.n1345 92.5
R1283 GND.n2347 GND.n2346 92.5
R1284 GND.n1587 GND.n1586 92.5
R1285 GND.n1836 GND.n1835 92.5
R1286 GND.n2085 GND.n2084 92.5
R1287 GND.n2325 GND.n2324 92.5
R1288 GND.n1174 GND.n1173 83.544
R1289 GND.n1933 GND.n1868 83.174
R1290 GND.n1941 GND.n1871 83.174
R1291 GND.n1949 GND.n1874 83.174
R1292 GND.n1904 GND.n1856 83.174
R1293 GND.n2037 GND.n1859 83.174
R1294 GND.n2021 GND.n1862 83.174
R1295 GND.n1684 GND.n1619 83.174
R1296 GND.n1692 GND.n1622 83.174
R1297 GND.n1700 GND.n1625 83.174
R1298 GND.n1655 GND.n1607 83.174
R1299 GND.n1788 GND.n1610 83.174
R1300 GND.n1772 GND.n1613 83.174
R1301 GND.n59 GND.n58 83.018
R1302 GND.n482 GND.n455 83.018
R1303 GND.n827 GND.n800 83.018
R1304 GND.n609 GND.n393 82.506
R1305 GND.n584 GND.n396 82.506
R1306 GND.n954 GND.n738 82.506
R1307 GND.n929 GND.n741 82.506
R1308 GND.n2228 GND.n2227 72.49
R1309 GND.n2209 GND.n2208 72.49
R1310 GND.n2004 GND.n1884 71.975
R1311 GND.n2005 GND.n1865 71.975
R1312 GND.n1755 GND.n1635 71.975
R1313 GND.n1756 GND.n1616 71.975
R1314 GND.n375 GND.t148 70.344
R1315 GND.n355 GND.t154 70.344
R1316 GND.n637 GND.t71 70.344
R1317 GND.n657 GND.t97 70.344
R1318 GND.n679 GND.t120 70.344
R1319 GND.n720 GND.t51 70.344
R1320 GND.n700 GND.t49 70.344
R1321 GND.n982 GND.t143 70.344
R1322 GND.n1002 GND.t69 70.344
R1323 GND.n1024 GND.t40 70.344
R1324 GND.n1065 GND.t92 70.344
R1325 GND.n1045 GND.t41 70.344
R1326 GND.n1326 GND.t104 70.344
R1327 GND.n1346 GND.t73 70.344
R1328 GND.n1587 GND.t81 70.344
R1329 GND.n1836 GND.t7 70.344
R1330 GND.n2085 GND.t107 70.344
R1331 GND.n1409 GND.n1400 67.542
R1332 GND.n1896 GND.n1893 66.905
R1333 GND.n1647 GND.n1644 66.905
R1334 GND.n1160 GND.n1153 66.905
R1335 GND.n472 GND.n469 66.28
R1336 GND.n817 GND.n814 66.28
R1337 GND.n1223 GND.n1222 55.696
R1338 GND.n1247 GND.n1103 55.696
R1339 GND.n1263 GND.n1080 55.696
R1340 GND.n144 GND.n143 55.345
R1341 GND.n168 GND.n167 55.345
R1342 GND.n541 GND.n426 55.345
R1343 GND.n556 GND.n555 55.345
R1344 GND.n620 GND.n619 55.345
R1345 GND.n886 GND.n771 55.345
R1346 GND.n901 GND.n900 55.345
R1347 GND.n965 GND.n964 55.345
R1348 GND.n1519 GND.n1370 52.37
R1349 GND.n1445 GND.n1370 52.37
R1350 GND.n26 GND.t153 34.332
R1351 GND.n391 GND.t66 34.33
R1352 GND.n736 GND.t121 34.33
R1353 GND.n1084 GND.t114 33.911
R1354 GND.n1084 GND.t91 33.911
R1355 GND.n391 GND.t147 33.607
R1356 GND.n736 GND.t50 33.607
R1357 GND.n26 GND.t45 33.605
R1358 GND.n2102 GND.n2101 31.928
R1359 GND.n1568 GND.n1567 31.928
R1360 GND.n1569 GND.n1568 31.928
R1361 GND.n1878 GND.n1876 31.644
R1362 GND.n1877 GND.n1876 31.644
R1363 GND.n1629 GND.n1627 31.644
R1364 GND.n1628 GND.n1627 31.644
R1365 GND.n1307 GND.n1306 31.644
R1366 GND.n1308 GND.n1307 31.644
R1367 GND.n24 GND.n23 31.364
R1368 GND.n400 GND.n398 31.364
R1369 GND.n399 GND.n398 31.364
R1370 GND.n745 GND.n743 31.364
R1371 GND.n744 GND.n743 31.364
R1372 GND.n11 GND.n10 31.034
R1373 GND.n273 GND.n272 31.034
R1374 GND.n293 GND.n292 31.034
R1375 GND.n313 GND.n312 31.034
R1376 GND.n335 GND.n334 31.034
R1377 GND.n376 GND.n367 31.034
R1378 GND.n356 GND.n347 31.034
R1379 GND.n638 GND.n629 31.034
R1380 GND.n658 GND.n649 31.034
R1381 GND.n680 GND.n671 31.034
R1382 GND.n721 GND.n712 31.034
R1383 GND.n701 GND.n692 31.034
R1384 GND.n983 GND.n974 31.034
R1385 GND.n1003 GND.n994 31.034
R1386 GND.n1025 GND.n1016 31.034
R1387 GND.n1066 GND.n1057 31.034
R1388 GND.n1046 GND.n1037 31.034
R1389 GND.n1327 GND.n1318 31.034
R1390 GND.n1347 GND.n1338 31.034
R1391 GND.n2357 GND.n2356 31.034
R1392 GND.n1588 GND.n1579 31.034
R1393 GND.n1837 GND.n1828 31.034
R1394 GND.n2086 GND.n2077 31.034
R1395 GND.n2335 GND.n2334 31.034
R1396 GND.n2111 GND.n2110 30.019
R1397 GND.n2117 GND.n2116 30.019
R1398 GND.n2316 GND.n2315 30.019
R1399 GND.n2103 GND.n2102 30.019
R1400 GND.n1404 GND.n1400 30.019
R1401 GND.n1409 GND.n1397 30.019
R1402 GND.n1570 GND.n1569 30.019
R1403 GND.n1567 GND.n1564 30.019
R1404 GND.n1896 GND.n1891 29.735
R1405 GND.n1893 GND.n1886 29.735
R1406 GND.n1878 GND.n1854 29.735
R1407 GND.n1882 GND.n1877 29.735
R1408 GND.n1647 GND.n1642 29.735
R1409 GND.n1644 GND.n1637 29.735
R1410 GND.n1629 GND.n1605 29.735
R1411 GND.n1633 GND.n1628 29.735
R1412 GND.n1156 GND.n1153 29.735
R1413 GND.n1160 GND.n1151 29.735
R1414 GND.n1309 GND.n1308 29.735
R1415 GND.n1306 GND.n1303 29.735
R1416 GND.n36 GND.n35 29.457
R1417 GND.n42 GND.n41 29.457
R1418 GND.n255 GND.n254 29.457
R1419 GND.n25 GND.n24 29.457
R1420 GND.n472 GND.n467 29.457
R1421 GND.n469 GND.n462 29.457
R1422 GND.n400 GND.n390 29.457
R1423 GND.n404 GND.n399 29.457
R1424 GND.n817 GND.n812 29.457
R1425 GND.n814 GND.n807 29.457
R1426 GND.n745 GND.n735 29.457
R1427 GND.n749 GND.n744 29.457
R1428 GND.n2210 GND.n2207 28.142
R1429 GND.n2232 GND.n2231 28.142
R1430 GND.n1443 GND.n1385 28.142
R1431 GND.n2120 GND.n2119 28.025
R1432 GND.n1412 GND.n1411 28.025
R1433 GND.n2013 GND.n2012 27.877
R1434 GND.n1997 GND.n1996 27.877
R1435 GND.n1764 GND.n1763 27.877
R1436 GND.n1748 GND.n1747 27.877
R1437 GND.n1224 GND.n1111 27.877
R1438 GND.n1239 GND.n1104 27.877
R1439 GND.n2066 GND.n1885 27.848
R1440 GND.n1817 GND.n1636 27.848
R1441 GND.n1163 GND.n1162 27.848
R1442 GND.n45 GND.n44 27.672
R1443 GND.n29 GND.n28 27.672
R1444 GND.n480 GND.n461 27.672
R1445 GND.n825 GND.n806 27.672
R1446 GND.n146 GND.n140 27.616
R1447 GND.n170 GND.n166 27.616
R1448 GND.n540 GND.n425 27.616
R1449 GND.n553 GND.n419 27.616
R1450 GND.n885 GND.n770 27.616
R1451 GND.n898 GND.n764 27.616
R1452 GND.n1450 GND.n1384 26.45
R1453 GND.n1475 GND.n1362 26.266
R1454 GND.n1172 GND.n1146 26.018
R1455 GND.n1275 GND.n1079 26.018
R1456 GND.n56 GND.n55 25.775
R1457 GND.n483 GND.n460 25.775
R1458 GND.n828 GND.n805 25.775
R1459 GND.n1438 GND.n1368 24.39
R1460 GND.n1220 GND.n1118 24.16
R1461 GND.n1250 GND.n1102 24.16
R1462 GND.n130 GND.n126 23.934
R1463 GND.n184 GND.n180 23.934
R1464 GND.n530 GND.n433 23.934
R1465 GND.n567 GND.n415 23.934
R1466 GND.n875 GND.n778 23.934
R1467 GND.n912 GND.n760 23.934
R1468 GND.n2195 GND.n2194 23.062
R1469 GND.n2243 GND.n2242 23.062
R1470 GND.n1455 GND.n1372 23.062
R1471 GND.n2020 GND.n1863 22.853
R1472 GND.n1932 GND.n1867 22.853
R1473 GND.n1771 GND.n1614 22.853
R1474 GND.n1683 GND.n1618 22.853
R1475 GND.n2144 GND.n2143 22.514
R1476 GND.n2292 GND.n2291 22.514
R1477 GND.n1471 GND.n1379 22.514
R1478 GND.n1905 GND.n1904 22.301
R1479 GND.n1949 GND.n1948 22.301
R1480 GND.n1656 GND.n1655 22.301
R1481 GND.n1700 GND.n1699 22.301
R1482 GND.n1176 GND.n1138 22.301
R1483 GND.n1272 GND.n1086 22.301
R1484 GND.n70 GND.n69 22.093
R1485 GND.n231 GND.n230 22.093
R1486 GND.n491 GND.n454 22.093
R1487 GND.n584 GND.n583 22.093
R1488 GND.n836 GND.n799 22.093
R1489 GND.n929 GND.n928 22.093
R1490 GND.n2184 GND.n2182 20.638
R1491 GND.n2257 GND.n2255 20.638
R1492 GND.n1433 GND.n1387 20.638
R1493 GND.n2029 GND.n2028 20.443
R1494 GND.n1985 GND.n1984 20.443
R1495 GND.n1780 GND.n1779 20.443
R1496 GND.n1736 GND.n1735 20.443
R1497 GND.n1207 GND.n1123 20.443
R1498 GND.n1260 GND.n1094 20.443
R1499 GND.n116 GND.n112 20.252
R1500 GND.n196 GND.n194 20.252
R1501 GND.n518 GND.n435 20.252
R1502 GND.n571 GND.n407 20.252
R1503 GND.n863 GND.n780 20.252
R1504 GND.n916 GND.n752 20.252
R1505 GND.n1459 GND.n1382 19.634
R1506 GND.n1467 GND.n1375 18.761
R1507 GND.n1187 GND.n1136 18.584
R1508 GND.n1291 GND.n1082 18.584
R1509 GND.n84 GND.n83 18.411
R1510 GND.n503 GND.n449 18.411
R1511 GND.n848 GND.n794 18.411
R1512 GND.n1428 GND.n1366 16.885
R1513 GND.n1199 GND.n1130 16.726
R1514 GND.n102 GND.n98 16.57
R1515 GND.n514 GND.n441 16.57
R1516 GND.n859 GND.n786 16.57
R1517 GND.n2170 GND.n2169 16.162
R1518 GND.n2268 GND.n2267 16.162
R1519 GND.n1463 GND.n1374 16.162
R1520 GND.n2036 GND.n1860 16.014
R1521 GND.n1940 GND.n1870 16.014
R1522 GND.n1787 GND.n1611 16.014
R1523 GND.n1691 GND.n1621 16.014
R1524 GND.n1088 GND.n1081 16.014
R1525 GND.n207 GND.n206 15.869
R1526 GND.n610 GND.n392 15.869
R1527 GND.n955 GND.n737 15.869
R1528 GND.n374 GND.n371 15.433
R1529 GND.n2 GND.n1 15.433
R1530 GND.n719 GND.n716 15.433
R1531 GND.n1064 GND.n1061 15.433
R1532 GND.n264 GND.n263 15.431
R1533 GND.n284 GND.n283 15.431
R1534 GND.n304 GND.n303 15.431
R1535 GND.n326 GND.n325 15.431
R1536 GND.n354 GND.n351 15.431
R1537 GND.n636 GND.n633 15.431
R1538 GND.n656 GND.n653 15.431
R1539 GND.n678 GND.n675 15.431
R1540 GND.n699 GND.n696 15.431
R1541 GND.n981 GND.n978 15.431
R1542 GND.n1001 GND.n998 15.431
R1543 GND.n1023 GND.n1020 15.431
R1544 GND.n1044 GND.n1041 15.431
R1545 GND.n1325 GND.n1322 15.431
R1546 GND.n1345 GND.n1342 15.431
R1547 GND.n2348 GND.n2347 15.431
R1548 GND.n1586 GND.n1583 15.431
R1549 GND.n1835 GND.n1832 15.431
R1550 GND.n2084 GND.n2081 15.431
R1551 GND.n2326 GND.n2325 15.431
R1552 GND.n2169 GND.n2168 15.009
R1553 GND.n2267 GND.n2266 15.009
R1554 GND.n1463 GND.n1381 15.009
R1555 GND.n2037 GND.n2036 14.867
R1556 GND.n1941 GND.n1940 14.867
R1557 GND.n1788 GND.n1787 14.867
R1558 GND.n1692 GND.n1691 14.867
R1559 GND.n1195 GND.n1130 14.867
R1560 GND.n1299 GND.n1088 14.867
R1561 GND.n98 GND.n97 14.728
R1562 GND.n206 GND.n205 14.728
R1563 GND.n507 GND.n441 14.728
R1564 GND.n610 GND.n609 14.728
R1565 GND.n852 GND.n786 14.728
R1566 GND.n955 GND.n954 14.728
R1567 GND.n374 GND.n373 13.552
R1568 GND.n381 GND.n380 13.552
R1569 GND.n354 GND.n353 13.552
R1570 GND.n361 GND.n360 13.552
R1571 GND.n636 GND.n635 13.552
R1572 GND.n643 GND.n642 13.552
R1573 GND.n656 GND.n655 13.552
R1574 GND.n663 GND.n662 13.552
R1575 GND.n678 GND.n677 13.552
R1576 GND.n685 GND.n684 13.552
R1577 GND.n719 GND.n718 13.552
R1578 GND.n726 GND.n725 13.552
R1579 GND.n699 GND.n698 13.552
R1580 GND.n706 GND.n705 13.552
R1581 GND.n981 GND.n980 13.552
R1582 GND.n988 GND.n987 13.552
R1583 GND.n1001 GND.n1000 13.552
R1584 GND.n1008 GND.n1007 13.552
R1585 GND.n1023 GND.n1022 13.552
R1586 GND.n1030 GND.n1029 13.552
R1587 GND.n1064 GND.n1063 13.552
R1588 GND.n1071 GND.n1070 13.552
R1589 GND.n1044 GND.n1043 13.552
R1590 GND.n1051 GND.n1050 13.552
R1591 GND.n1325 GND.n1324 13.552
R1592 GND.n1332 GND.n1331 13.552
R1593 GND.n1345 GND.n1344 13.552
R1594 GND.n1352 GND.n1351 13.552
R1595 GND.n1586 GND.n1585 13.552
R1596 GND.n1593 GND.n1592 13.552
R1597 GND.n1835 GND.n1834 13.552
R1598 GND.n1842 GND.n1841 13.552
R1599 GND.n2084 GND.n2083 13.552
R1600 GND.n2091 GND.n2090 13.552
R1601 GND.n2159 GND.n2157 13.133
R1602 GND.n2282 GND.n2280 13.133
R1603 GND.n1423 GND.n1389 13.133
R1604 GND.n2045 GND.n2044 13.009
R1605 GND.n1971 GND.n1970 13.009
R1606 GND.n1796 GND.n1795 13.009
R1607 GND.n1722 GND.n1721 13.009
R1608 GND.n1187 GND.n1132 13.009
R1609 GND.n88 GND.n84 12.887
R1610 GND.n221 GND.n219 12.887
R1611 GND.n503 GND.n447 12.887
R1612 GND.n578 GND.n577 12.887
R1613 GND.n848 GND.n792 12.887
R1614 GND.n923 GND.n922 12.887
R1615 GND.n2131 GND.n2130 12.845
R1616 GND.n2305 GND.n2304 12.845
R1617 GND.n2132 GND.n2131 12.845
R1618 GND.n2304 GND.n2303 12.845
R1619 GND.n1391 GND.n1363 12.845
R1620 GND.n1414 GND.n1363 12.845
R1621 GND.n1887 GND.n1855 12.727
R1622 GND.n1956 GND.n1875 12.727
R1623 GND.n2057 GND.n1855 12.727
R1624 GND.n1875 GND.n1853 12.727
R1625 GND.n1638 GND.n1606 12.727
R1626 GND.n1707 GND.n1626 12.727
R1627 GND.n1808 GND.n1606 12.727
R1628 GND.n1626 GND.n1604 12.727
R1629 GND.n1467 GND.n1380 12.649
R1630 GND.n244 GND.n243 12.61
R1631 GND.n243 GND.n242 12.61
R1632 GND.n591 GND.n397 12.61
R1633 GND.n397 GND.n389 12.61
R1634 GND.n936 GND.n742 12.61
R1635 GND.n742 GND.n734 12.61
R1636 GND.n1291 GND.n1087 12.532
R1637 GND.n1459 GND.n1373 11.257
R1638 GND.n1207 GND.n1125 11.15
R1639 GND.n1264 GND.n1094 11.15
R1640 GND.n112 GND.n111 11.046
R1641 GND.n194 GND.n193 11.046
R1642 GND.n518 GND.n439 11.046
R1643 GND.n618 GND.n407 11.046
R1644 GND.n863 GND.n784 11.046
R1645 GND.n963 GND.n752 11.046
R1646 GND.n1552 GND.n1390 11.045
R1647 GND.n1392 GND.n1390 11.045
R1648 GND.n1300 GND.n1080 9.734
R1649 GND.n2114 GND.n2113 9.413
R1650 GND.n1403 GND.n1402 9.413
R1651 GND.n1899 GND.n1898 9.411
R1652 GND.n1650 GND.n1649 9.411
R1653 GND.n1155 GND.n1154 9.411
R1654 GND.n39 GND.n38 9.41
R1655 GND.n475 GND.n474 9.41
R1656 GND.n820 GND.n819 9.41
R1657 GND.n1552 GND.n1364 9.38
R1658 GND.n2106 GND.n2105 9.33
R1659 GND.n1563 GND.n1358 9.33
R1660 GND.n1883 GND.n1849 9.329
R1661 GND.n1634 GND.n1600 9.329
R1662 GND.n1302 GND.n1075 9.329
R1663 GND.n31 GND.n30 9.329
R1664 GND.n405 GND.n385 9.329
R1665 GND.n750 GND.n730 9.329
R1666 GND.n252 GND.n251 9.3
R1667 GND.n239 GND.n238 9.3
R1668 GND.n227 GND.n226 9.3
R1669 GND.n214 GND.n213 9.3
R1670 GND.n202 GND.n201 9.3
R1671 GND.n190 GND.n189 9.3
R1672 GND.n176 GND.n175 9.3
R1673 GND.n160 GND.n159 9.3
R1674 GND.n150 GND.n149 9.3
R1675 GND.n134 GND.n133 9.3
R1676 GND.n120 GND.n119 9.3
R1677 GND.n106 GND.n105 9.3
R1678 GND.n92 GND.n91 9.3
R1679 GND.n78 GND.n77 9.3
R1680 GND.n64 GND.n63 9.3
R1681 GND.n50 GND.n49 9.3
R1682 GND.n52 GND.n51 9.3
R1683 GND.n48 GND.n47 9.3
R1684 GND.n47 GND.n46 9.3
R1685 GND.n46 GND.n45 9.3
R1686 GND.n66 GND.n65 9.3
R1687 GND.n62 GND.n61 9.3
R1688 GND.n61 GND.n60 9.3
R1689 GND.n60 GND.n59 9.3
R1690 GND.n80 GND.n79 9.3
R1691 GND.n76 GND.n75 9.3
R1692 GND.n75 GND.n74 9.3
R1693 GND.n74 GND.n73 9.3
R1694 GND.n94 GND.n93 9.3
R1695 GND.n90 GND.n89 9.3
R1696 GND.n89 GND.n88 9.3
R1697 GND.n88 GND.n87 9.3
R1698 GND.n108 GND.n107 9.3
R1699 GND.n104 GND.n103 9.3
R1700 GND.n103 GND.n102 9.3
R1701 GND.n102 GND.n101 9.3
R1702 GND.n122 GND.n121 9.3
R1703 GND.n118 GND.n117 9.3
R1704 GND.n117 GND.n116 9.3
R1705 GND.n116 GND.n115 9.3
R1706 GND.n136 GND.n135 9.3
R1707 GND.n132 GND.n131 9.3
R1708 GND.n131 GND.n130 9.3
R1709 GND.n130 GND.n129 9.3
R1710 GND.n152 GND.n151 9.3
R1711 GND.n148 GND.n147 9.3
R1712 GND.n147 GND.n146 9.3
R1713 GND.n146 GND.n145 9.3
R1714 GND.n158 GND.n157 9.3
R1715 GND.n172 GND.n171 9.3
R1716 GND.n171 GND.n170 9.3
R1717 GND.n170 GND.n169 9.3
R1718 GND.n174 GND.n173 9.3
R1719 GND.n186 GND.n185 9.3
R1720 GND.n185 GND.n184 9.3
R1721 GND.n184 GND.n183 9.3
R1722 GND.n188 GND.n187 9.3
R1723 GND.n198 GND.n197 9.3
R1724 GND.n197 GND.n196 9.3
R1725 GND.n196 GND.n195 9.3
R1726 GND.n200 GND.n199 9.3
R1727 GND.n210 GND.n209 9.3
R1728 GND.n209 GND.n208 9.3
R1729 GND.n212 GND.n211 9.3
R1730 GND.n223 GND.n222 9.3
R1731 GND.n222 GND.n221 9.3
R1732 GND.n225 GND.n224 9.3
R1733 GND.n235 GND.n234 9.3
R1734 GND.n234 GND.n233 9.3
R1735 GND.n237 GND.n236 9.3
R1736 GND.n248 GND.n247 9.3
R1737 GND.n247 GND.n246 9.3
R1738 GND.n250 GND.n249 9.3
R1739 GND.n259 GND.n258 9.3
R1740 GND.n258 GND.n257 9.3
R1741 GND.n17 GND.n16 9.3
R1742 GND.n6 GND.n5 9.3
R1743 GND.n4 GND.n3 9.3
R1744 GND.n13 GND.n12 9.3
R1745 GND.n12 GND.n11 9.3
R1746 GND.n15 GND.n14 9.3
R1747 GND.n19 GND.n18 9.3
R1748 GND.n279 GND.n278 9.3
R1749 GND.n268 GND.n267 9.3
R1750 GND.n266 GND.n265 9.3
R1751 GND.n275 GND.n274 9.3
R1752 GND.n274 GND.n273 9.3
R1753 GND.n277 GND.n276 9.3
R1754 GND.n281 GND.n280 9.3
R1755 GND.n299 GND.n298 9.3
R1756 GND.n288 GND.n287 9.3
R1757 GND.n286 GND.n285 9.3
R1758 GND.n295 GND.n294 9.3
R1759 GND.n294 GND.n293 9.3
R1760 GND.n297 GND.n296 9.3
R1761 GND.n301 GND.n300 9.3
R1762 GND.n319 GND.n318 9.3
R1763 GND.n308 GND.n307 9.3
R1764 GND.n306 GND.n305 9.3
R1765 GND.n315 GND.n314 9.3
R1766 GND.n314 GND.n313 9.3
R1767 GND.n317 GND.n316 9.3
R1768 GND.n321 GND.n320 9.3
R1769 GND.n2313 GND.n2312 9.3
R1770 GND.n2300 GND.n2299 9.3
R1771 GND.n2288 GND.n2287 9.3
R1772 GND.n2275 GND.n2274 9.3
R1773 GND.n2263 GND.n2262 9.3
R1774 GND.n2250 GND.n2249 9.3
R1775 GND.n2238 GND.n2237 9.3
R1776 GND.n2224 GND.n2223 9.3
R1777 GND.n2214 GND.n2213 9.3
R1778 GND.n2200 GND.n2199 9.3
R1779 GND.n2188 GND.n2187 9.3
R1780 GND.n2175 GND.n2174 9.3
R1781 GND.n2163 GND.n2162 9.3
R1782 GND.n2150 GND.n2149 9.3
R1783 GND.n2138 GND.n2137 9.3
R1784 GND.n2125 GND.n2124 9.3
R1785 GND.n2216 GND.n2215 9.3
R1786 GND.n2202 GND.n2201 9.3
R1787 GND.n2190 GND.n2189 9.3
R1788 GND.n2177 GND.n2176 9.3
R1789 GND.n2165 GND.n2164 9.3
R1790 GND.n2152 GND.n2151 9.3
R1791 GND.n2140 GND.n2139 9.3
R1792 GND.n2127 GND.n2126 9.3
R1793 GND.n2123 GND.n2122 9.3
R1794 GND.n2122 GND.n2121 9.3
R1795 GND.n2121 GND.n2120 9.3
R1796 GND.n2136 GND.n2135 9.3
R1797 GND.n2135 GND.n2134 9.3
R1798 GND.n2148 GND.n2147 9.3
R1799 GND.n2147 GND.n2146 9.3
R1800 GND.n2161 GND.n2160 9.3
R1801 GND.n2160 GND.n2159 9.3
R1802 GND.n2173 GND.n2172 9.3
R1803 GND.n2172 GND.n2171 9.3
R1804 GND.n2186 GND.n2185 9.3
R1805 GND.n2185 GND.n2184 9.3
R1806 GND.n2198 GND.n2197 9.3
R1807 GND.n2197 GND.n2196 9.3
R1808 GND.n2212 GND.n2211 9.3
R1809 GND.n2211 GND.n2210 9.3
R1810 GND.n2222 GND.n2221 9.3
R1811 GND.n2234 GND.n2233 9.3
R1812 GND.n2233 GND.n2232 9.3
R1813 GND.n2236 GND.n2235 9.3
R1814 GND.n2246 GND.n2245 9.3
R1815 GND.n2245 GND.n2244 9.3
R1816 GND.n2248 GND.n2247 9.3
R1817 GND.n2259 GND.n2258 9.3
R1818 GND.n2258 GND.n2257 9.3
R1819 GND.n2261 GND.n2260 9.3
R1820 GND.n2271 GND.n2270 9.3
R1821 GND.n2270 GND.n2269 9.3
R1822 GND.n2273 GND.n2272 9.3
R1823 GND.n2284 GND.n2283 9.3
R1824 GND.n2283 GND.n2282 9.3
R1825 GND.n2286 GND.n2285 9.3
R1826 GND.n2296 GND.n2295 9.3
R1827 GND.n2295 GND.n2294 9.3
R1828 GND.n2298 GND.n2297 9.3
R1829 GND.n2309 GND.n2308 9.3
R1830 GND.n2308 GND.n2307 9.3
R1831 GND.n2311 GND.n2310 9.3
R1832 GND.n2320 GND.n2319 9.3
R1833 GND.n2319 GND.n2318 9.3
R1834 GND.n341 GND.n340 9.3
R1835 GND.n330 GND.n329 9.3
R1836 GND.n328 GND.n327 9.3
R1837 GND.n337 GND.n336 9.3
R1838 GND.n336 GND.n335 9.3
R1839 GND.n339 GND.n338 9.3
R1840 GND.n343 GND.n342 9.3
R1841 GND.n387 GND.n386 9.3
R1842 GND.n594 GND.n582 9.3
R1843 GND.n601 GND.n576 9.3
R1844 GND.n606 GND.n605 9.3
R1845 GND.n614 GND.n410 9.3
R1846 GND.n412 GND.n411 9.3
R1847 GND.n561 GND.n560 9.3
R1848 GND.n550 GND.n422 9.3
R1849 GND.n536 GND.n429 9.3
R1850 GND.n532 GND.n430 9.3
R1851 GND.n522 GND.n436 9.3
R1852 GND.n511 GND.n444 9.3
R1853 GND.n446 GND.n445 9.3
R1854 GND.n497 GND.n451 9.3
R1855 GND.n487 GND.n457 9.3
R1856 GND.n476 GND.n465 9.3
R1857 GND.n535 GND.n424 9.3
R1858 GND.n534 GND.n533 9.3
R1859 GND.n524 GND.n523 9.3
R1860 GND.n443 GND.n437 9.3
R1861 GND.n510 GND.n509 9.3
R1862 GND.n499 GND.n498 9.3
R1863 GND.n489 GND.n488 9.3
R1864 GND.n464 GND.n458 9.3
R1865 GND.n478 GND.n477 9.3
R1866 GND.n479 GND.n478 9.3
R1867 GND.n480 GND.n479 9.3
R1868 GND.n486 GND.n485 9.3
R1869 GND.n485 GND.n456 9.3
R1870 GND.n456 GND.n455 9.3
R1871 GND.n496 GND.n453 9.3
R1872 GND.n496 GND.n495 9.3
R1873 GND.n495 GND.n494 9.3
R1874 GND.n501 GND.n500 9.3
R1875 GND.n501 GND.n447 9.3
R1876 GND.n505 GND.n447 9.3
R1877 GND.n513 GND.n512 9.3
R1878 GND.n514 GND.n513 9.3
R1879 GND.n515 GND.n514 9.3
R1880 GND.n521 GND.n520 9.3
R1881 GND.n520 GND.n435 9.3
R1882 GND.n435 GND.n434 9.3
R1883 GND.n531 GND.n432 9.3
R1884 GND.n531 GND.n530 9.3
R1885 GND.n530 GND.n529 9.3
R1886 GND.n538 GND.n537 9.3
R1887 GND.n538 GND.n425 9.3
R1888 GND.n542 GND.n425 9.3
R1889 GND.n549 GND.n548 9.3
R1890 GND.n552 GND.n551 9.3
R1891 GND.n553 GND.n552 9.3
R1892 GND.n554 GND.n553 9.3
R1893 GND.n559 GND.n417 9.3
R1894 GND.n562 GND.n416 9.3
R1895 GND.n416 GND.n415 9.3
R1896 GND.n415 GND.n414 9.3
R1897 GND.n564 GND.n563 9.3
R1898 GND.n573 GND.n572 9.3
R1899 GND.n572 GND.n571 9.3
R1900 GND.n571 GND.n570 9.3
R1901 GND.n616 GND.n615 9.3
R1902 GND.n613 GND.n612 9.3
R1903 GND.n612 GND.n408 9.3
R1904 GND.n607 GND.n574 9.3
R1905 GND.n604 GND.n575 9.3
R1906 GND.n577 GND.n575 9.3
R1907 GND.n603 GND.n602 9.3
R1908 GND.n600 GND.n597 9.3
R1909 GND.n600 GND.n599 9.3
R1910 GND.n596 GND.n595 9.3
R1911 GND.n593 GND.n590 9.3
R1912 GND.n593 GND.n592 9.3
R1913 GND.n589 GND.n588 9.3
R1914 GND.n624 GND.n623 9.3
R1915 GND.n623 GND.n622 9.3
R1916 GND.n366 GND.n365 9.3
R1917 GND.n370 GND.n369 9.3
R1918 GND.n373 GND.n372 9.3
R1919 GND.n378 GND.n377 9.3
R1920 GND.n377 GND.n376 9.3
R1921 GND.n380 GND.n379 9.3
R1922 GND.n384 GND.n383 9.3
R1923 GND.n346 GND.n345 9.3
R1924 GND.n350 GND.n349 9.3
R1925 GND.n353 GND.n352 9.3
R1926 GND.n358 GND.n357 9.3
R1927 GND.n357 GND.n356 9.3
R1928 GND.n360 GND.n359 9.3
R1929 GND.n364 GND.n363 9.3
R1930 GND.n628 GND.n627 9.3
R1931 GND.n632 GND.n631 9.3
R1932 GND.n635 GND.n634 9.3
R1933 GND.n640 GND.n639 9.3
R1934 GND.n639 GND.n638 9.3
R1935 GND.n642 GND.n641 9.3
R1936 GND.n646 GND.n645 9.3
R1937 GND.n648 GND.n647 9.3
R1938 GND.n652 GND.n651 9.3
R1939 GND.n655 GND.n654 9.3
R1940 GND.n660 GND.n659 9.3
R1941 GND.n659 GND.n658 9.3
R1942 GND.n662 GND.n661 9.3
R1943 GND.n666 GND.n665 9.3
R1944 GND.n1851 GND.n1850 9.3
R1945 GND.n1959 GND.n1947 9.3
R1946 GND.n1966 GND.n1944 9.3
R1947 GND.n1973 GND.n1939 9.3
R1948 GND.n1980 GND.n1936 9.3
R1949 GND.n1987 GND.n1931 9.3
R1950 GND.n1930 GND.n1928 9.3
R1951 GND.n2000 GND.n1925 9.3
R1952 GND.n2009 GND.n1920 9.3
R1953 GND.n1921 GND.n1918 9.3
R1954 GND.n2025 GND.n1914 9.3
R1955 GND.n1915 GND.n1912 9.3
R1956 GND.n2041 GND.n1909 9.3
R1957 GND.n1907 GND.n1902 9.3
R1958 GND.n2054 GND.n2053 9.3
R1959 GND.n2062 GND.n1889 9.3
R1960 GND.n2008 GND.n2007 9.3
R1961 GND.n1922 GND.n1919 9.3
R1962 GND.n2024 GND.n2023 9.3
R1963 GND.n1916 GND.n1913 9.3
R1964 GND.n2040 GND.n2039 9.3
R1965 GND.n1910 GND.n1908 9.3
R1966 GND.n2052 GND.n1901 9.3
R1967 GND.n2061 GND.n2060 9.3
R1968 GND.n2064 GND.n2063 9.3
R1969 GND.n2065 GND.n2064 9.3
R1970 GND.n2066 GND.n2065 9.3
R1971 GND.n2055 GND.n1900 9.3
R1972 GND.n2056 GND.n2055 9.3
R1973 GND.n2051 GND.n2050 9.3
R1974 GND.n2050 GND.n2049 9.3
R1975 GND.n2043 GND.n2042 9.3
R1976 GND.n2044 GND.n2043 9.3
R1977 GND.n2034 GND.n1911 9.3
R1978 GND.n2034 GND.n2033 9.3
R1979 GND.n2027 GND.n2026 9.3
R1980 GND.n2028 GND.n2027 9.3
R1981 GND.n2018 GND.n1917 9.3
R1982 GND.n2018 GND.n2017 9.3
R1983 GND.n2011 GND.n2010 9.3
R1984 GND.n2012 GND.n2011 9.3
R1985 GND.n2002 GND.n2001 9.3
R1986 GND.n1999 GND.n1998 9.3
R1987 GND.n1998 GND.n1997 9.3
R1988 GND.n1927 GND.n1926 9.3
R1989 GND.n1991 GND.n1990 9.3
R1990 GND.n1992 GND.n1991 9.3
R1991 GND.n1989 GND.n1988 9.3
R1992 GND.n1986 GND.n1983 9.3
R1993 GND.n1986 GND.n1985 9.3
R1994 GND.n1982 GND.n1981 9.3
R1995 GND.n1979 GND.n1976 9.3
R1996 GND.n1979 GND.n1978 9.3
R1997 GND.n1975 GND.n1974 9.3
R1998 GND.n1972 GND.n1969 9.3
R1999 GND.n1972 GND.n1971 9.3
R2000 GND.n1968 GND.n1967 9.3
R2001 GND.n1965 GND.n1962 9.3
R2002 GND.n1965 GND.n1964 9.3
R2003 GND.n1961 GND.n1960 9.3
R2004 GND.n1958 GND.n1955 9.3
R2005 GND.n1958 GND.n1957 9.3
R2006 GND.n1954 GND.n1953 9.3
R2007 GND.n2071 GND.n2070 9.3
R2008 GND.n2070 GND.n2069 9.3
R2009 GND.n670 GND.n669 9.3
R2010 GND.n674 GND.n673 9.3
R2011 GND.n677 GND.n676 9.3
R2012 GND.n682 GND.n681 9.3
R2013 GND.n681 GND.n680 9.3
R2014 GND.n684 GND.n683 9.3
R2015 GND.n688 GND.n687 9.3
R2016 GND.n732 GND.n731 9.3
R2017 GND.n939 GND.n927 9.3
R2018 GND.n946 GND.n921 9.3
R2019 GND.n951 GND.n950 9.3
R2020 GND.n959 GND.n755 9.3
R2021 GND.n757 GND.n756 9.3
R2022 GND.n906 GND.n905 9.3
R2023 GND.n895 GND.n767 9.3
R2024 GND.n881 GND.n774 9.3
R2025 GND.n877 GND.n775 9.3
R2026 GND.n867 GND.n781 9.3
R2027 GND.n856 GND.n789 9.3
R2028 GND.n791 GND.n790 9.3
R2029 GND.n842 GND.n796 9.3
R2030 GND.n832 GND.n802 9.3
R2031 GND.n821 GND.n810 9.3
R2032 GND.n880 GND.n769 9.3
R2033 GND.n879 GND.n878 9.3
R2034 GND.n869 GND.n868 9.3
R2035 GND.n788 GND.n782 9.3
R2036 GND.n855 GND.n854 9.3
R2037 GND.n844 GND.n843 9.3
R2038 GND.n834 GND.n833 9.3
R2039 GND.n809 GND.n803 9.3
R2040 GND.n823 GND.n822 9.3
R2041 GND.n824 GND.n823 9.3
R2042 GND.n825 GND.n824 9.3
R2043 GND.n831 GND.n830 9.3
R2044 GND.n830 GND.n801 9.3
R2045 GND.n801 GND.n800 9.3
R2046 GND.n841 GND.n798 9.3
R2047 GND.n841 GND.n840 9.3
R2048 GND.n840 GND.n839 9.3
R2049 GND.n846 GND.n845 9.3
R2050 GND.n846 GND.n792 9.3
R2051 GND.n850 GND.n792 9.3
R2052 GND.n858 GND.n857 9.3
R2053 GND.n859 GND.n858 9.3
R2054 GND.n860 GND.n859 9.3
R2055 GND.n866 GND.n865 9.3
R2056 GND.n865 GND.n780 9.3
R2057 GND.n780 GND.n779 9.3
R2058 GND.n876 GND.n777 9.3
R2059 GND.n876 GND.n875 9.3
R2060 GND.n875 GND.n874 9.3
R2061 GND.n883 GND.n882 9.3
R2062 GND.n883 GND.n770 9.3
R2063 GND.n887 GND.n770 9.3
R2064 GND.n894 GND.n893 9.3
R2065 GND.n897 GND.n896 9.3
R2066 GND.n898 GND.n897 9.3
R2067 GND.n899 GND.n898 9.3
R2068 GND.n904 GND.n762 9.3
R2069 GND.n907 GND.n761 9.3
R2070 GND.n761 GND.n760 9.3
R2071 GND.n760 GND.n759 9.3
R2072 GND.n909 GND.n908 9.3
R2073 GND.n918 GND.n917 9.3
R2074 GND.n917 GND.n916 9.3
R2075 GND.n916 GND.n915 9.3
R2076 GND.n961 GND.n960 9.3
R2077 GND.n958 GND.n957 9.3
R2078 GND.n957 GND.n753 9.3
R2079 GND.n952 GND.n919 9.3
R2080 GND.n949 GND.n920 9.3
R2081 GND.n922 GND.n920 9.3
R2082 GND.n948 GND.n947 9.3
R2083 GND.n945 GND.n942 9.3
R2084 GND.n945 GND.n944 9.3
R2085 GND.n941 GND.n940 9.3
R2086 GND.n938 GND.n935 9.3
R2087 GND.n938 GND.n937 9.3
R2088 GND.n934 GND.n933 9.3
R2089 GND.n969 GND.n968 9.3
R2090 GND.n968 GND.n967 9.3
R2091 GND.n711 GND.n710 9.3
R2092 GND.n715 GND.n714 9.3
R2093 GND.n718 GND.n717 9.3
R2094 GND.n723 GND.n722 9.3
R2095 GND.n722 GND.n721 9.3
R2096 GND.n725 GND.n724 9.3
R2097 GND.n729 GND.n728 9.3
R2098 GND.n691 GND.n690 9.3
R2099 GND.n695 GND.n694 9.3
R2100 GND.n698 GND.n697 9.3
R2101 GND.n703 GND.n702 9.3
R2102 GND.n702 GND.n701 9.3
R2103 GND.n705 GND.n704 9.3
R2104 GND.n709 GND.n708 9.3
R2105 GND.n973 GND.n972 9.3
R2106 GND.n977 GND.n976 9.3
R2107 GND.n980 GND.n979 9.3
R2108 GND.n985 GND.n984 9.3
R2109 GND.n984 GND.n983 9.3
R2110 GND.n987 GND.n986 9.3
R2111 GND.n991 GND.n990 9.3
R2112 GND.n993 GND.n992 9.3
R2113 GND.n997 GND.n996 9.3
R2114 GND.n1000 GND.n999 9.3
R2115 GND.n1005 GND.n1004 9.3
R2116 GND.n1004 GND.n1003 9.3
R2117 GND.n1007 GND.n1006 9.3
R2118 GND.n1011 GND.n1010 9.3
R2119 GND.n1602 GND.n1601 9.3
R2120 GND.n1710 GND.n1698 9.3
R2121 GND.n1717 GND.n1695 9.3
R2122 GND.n1724 GND.n1690 9.3
R2123 GND.n1731 GND.n1687 9.3
R2124 GND.n1738 GND.n1682 9.3
R2125 GND.n1681 GND.n1679 9.3
R2126 GND.n1751 GND.n1676 9.3
R2127 GND.n1760 GND.n1671 9.3
R2128 GND.n1672 GND.n1669 9.3
R2129 GND.n1776 GND.n1665 9.3
R2130 GND.n1666 GND.n1663 9.3
R2131 GND.n1792 GND.n1660 9.3
R2132 GND.n1658 GND.n1653 9.3
R2133 GND.n1805 GND.n1804 9.3
R2134 GND.n1813 GND.n1640 9.3
R2135 GND.n1759 GND.n1758 9.3
R2136 GND.n1673 GND.n1670 9.3
R2137 GND.n1775 GND.n1774 9.3
R2138 GND.n1667 GND.n1664 9.3
R2139 GND.n1791 GND.n1790 9.3
R2140 GND.n1661 GND.n1659 9.3
R2141 GND.n1803 GND.n1652 9.3
R2142 GND.n1812 GND.n1811 9.3
R2143 GND.n1815 GND.n1814 9.3
R2144 GND.n1816 GND.n1815 9.3
R2145 GND.n1817 GND.n1816 9.3
R2146 GND.n1806 GND.n1651 9.3
R2147 GND.n1807 GND.n1806 9.3
R2148 GND.n1802 GND.n1801 9.3
R2149 GND.n1801 GND.n1800 9.3
R2150 GND.n1794 GND.n1793 9.3
R2151 GND.n1795 GND.n1794 9.3
R2152 GND.n1785 GND.n1662 9.3
R2153 GND.n1785 GND.n1784 9.3
R2154 GND.n1778 GND.n1777 9.3
R2155 GND.n1779 GND.n1778 9.3
R2156 GND.n1769 GND.n1668 9.3
R2157 GND.n1769 GND.n1768 9.3
R2158 GND.n1762 GND.n1761 9.3
R2159 GND.n1763 GND.n1762 9.3
R2160 GND.n1753 GND.n1752 9.3
R2161 GND.n1750 GND.n1749 9.3
R2162 GND.n1749 GND.n1748 9.3
R2163 GND.n1678 GND.n1677 9.3
R2164 GND.n1742 GND.n1741 9.3
R2165 GND.n1743 GND.n1742 9.3
R2166 GND.n1740 GND.n1739 9.3
R2167 GND.n1737 GND.n1734 9.3
R2168 GND.n1737 GND.n1736 9.3
R2169 GND.n1733 GND.n1732 9.3
R2170 GND.n1730 GND.n1727 9.3
R2171 GND.n1730 GND.n1729 9.3
R2172 GND.n1726 GND.n1725 9.3
R2173 GND.n1723 GND.n1720 9.3
R2174 GND.n1723 GND.n1722 9.3
R2175 GND.n1719 GND.n1718 9.3
R2176 GND.n1716 GND.n1713 9.3
R2177 GND.n1716 GND.n1715 9.3
R2178 GND.n1712 GND.n1711 9.3
R2179 GND.n1709 GND.n1706 9.3
R2180 GND.n1709 GND.n1708 9.3
R2181 GND.n1705 GND.n1704 9.3
R2182 GND.n1822 GND.n1821 9.3
R2183 GND.n1821 GND.n1820 9.3
R2184 GND.n1015 GND.n1014 9.3
R2185 GND.n1019 GND.n1018 9.3
R2186 GND.n1022 GND.n1021 9.3
R2187 GND.n1027 GND.n1026 9.3
R2188 GND.n1026 GND.n1025 9.3
R2189 GND.n1029 GND.n1028 9.3
R2190 GND.n1033 GND.n1032 9.3
R2191 GND.n1077 GND.n1076 9.3
R2192 GND.n1283 GND.n1271 9.3
R2193 GND.n1288 GND.n1287 9.3
R2194 GND.n1295 GND.n1091 9.3
R2195 GND.n1093 GND.n1092 9.3
R2196 GND.n1255 GND.n1098 9.3
R2197 GND.n1242 GND.n1106 9.3
R2198 GND.n1108 GND.n1107 9.3
R2199 GND.n1228 GND.n1227 9.3
R2200 GND.n1217 GND.n1120 9.3
R2201 GND.n1122 GND.n1121 9.3
R2202 GND.n1201 GND.n1127 9.3
R2203 GND.n1191 GND.n1133 9.3
R2204 GND.n1180 GND.n1141 9.3
R2205 GND.n1143 GND.n1142 9.3
R2206 GND.n1166 GND.n1148 9.3
R2207 GND.n1229 GND.n1112 9.3
R2208 GND.n1216 GND.n1215 9.3
R2209 GND.n1214 GND.n1213 9.3
R2210 GND.n1203 GND.n1202 9.3
R2211 GND.n1193 GND.n1192 9.3
R2212 GND.n1140 GND.n1134 9.3
R2213 GND.n1179 GND.n1178 9.3
R2214 GND.n1168 GND.n1167 9.3
R2215 GND.n1165 GND.n1150 9.3
R2216 GND.n1165 GND.n1164 9.3
R2217 GND.n1164 GND.n1163 9.3
R2218 GND.n1170 GND.n1169 9.3
R2219 GND.n1170 GND.n1144 9.3
R2220 GND.n1174 GND.n1144 9.3
R2221 GND.n1182 GND.n1181 9.3
R2222 GND.n1183 GND.n1182 9.3
R2223 GND.n1184 GND.n1183 9.3
R2224 GND.n1190 GND.n1189 9.3
R2225 GND.n1189 GND.n1132 9.3
R2226 GND.n1132 GND.n1131 9.3
R2227 GND.n1200 GND.n1129 9.3
R2228 GND.n1200 GND.n1199 9.3
R2229 GND.n1199 GND.n1198 9.3
R2230 GND.n1205 GND.n1204 9.3
R2231 GND.n1205 GND.n1123 9.3
R2232 GND.n1209 GND.n1123 9.3
R2233 GND.n1219 GND.n1218 9.3
R2234 GND.n1220 GND.n1219 9.3
R2235 GND.n1221 GND.n1220 9.3
R2236 GND.n1226 GND.n1114 9.3
R2237 GND.n1226 GND.n1111 9.3
R2238 GND.n1111 GND.n1110 9.3
R2239 GND.n1231 GND.n1230 9.3
R2240 GND.n1241 GND.n1240 9.3
R2241 GND.n1240 GND.n1239 9.3
R2242 GND.n1239 GND.n1238 9.3
R2243 GND.n1244 GND.n1243 9.3
R2244 GND.n1101 GND.n1100 9.3
R2245 GND.n1102 GND.n1101 9.3
R2246 GND.n1248 GND.n1102 9.3
R2247 GND.n1254 GND.n1253 9.3
R2248 GND.n1259 GND.n1258 9.3
R2249 GND.n1260 GND.n1259 9.3
R2250 GND.n1261 GND.n1260 9.3
R2251 GND.n1257 GND.n1256 9.3
R2252 GND.n1267 GND.n1266 9.3
R2253 GND.n1266 GND.n1265 9.3
R2254 GND.n1297 GND.n1296 9.3
R2255 GND.n1294 GND.n1293 9.3
R2256 GND.n1293 GND.n1089 9.3
R2257 GND.n1289 GND.n1268 9.3
R2258 GND.n1286 GND.n1270 9.3
R2259 GND.n1270 GND.n1269 9.3
R2260 GND.n1285 GND.n1284 9.3
R2261 GND.n1282 GND.n1280 9.3
R2262 GND.n1282 GND.n1281 9.3
R2263 GND.n1279 GND.n1278 9.3
R2264 GND.n1313 GND.n1312 9.3
R2265 GND.n1312 GND.n1311 9.3
R2266 GND.n1056 GND.n1055 9.3
R2267 GND.n1060 GND.n1059 9.3
R2268 GND.n1063 GND.n1062 9.3
R2269 GND.n1068 GND.n1067 9.3
R2270 GND.n1067 GND.n1066 9.3
R2271 GND.n1070 GND.n1069 9.3
R2272 GND.n1074 GND.n1073 9.3
R2273 GND.n1036 GND.n1035 9.3
R2274 GND.n1040 GND.n1039 9.3
R2275 GND.n1043 GND.n1042 9.3
R2276 GND.n1048 GND.n1047 9.3
R2277 GND.n1047 GND.n1046 9.3
R2278 GND.n1050 GND.n1049 9.3
R2279 GND.n1054 GND.n1053 9.3
R2280 GND.n1317 GND.n1316 9.3
R2281 GND.n1321 GND.n1320 9.3
R2282 GND.n1324 GND.n1323 9.3
R2283 GND.n1329 GND.n1328 9.3
R2284 GND.n1328 GND.n1327 9.3
R2285 GND.n1331 GND.n1330 9.3
R2286 GND.n1335 GND.n1334 9.3
R2287 GND.n1337 GND.n1336 9.3
R2288 GND.n1341 GND.n1340 9.3
R2289 GND.n1344 GND.n1343 9.3
R2290 GND.n1349 GND.n1348 9.3
R2291 GND.n1348 GND.n1347 9.3
R2292 GND.n1351 GND.n1350 9.3
R2293 GND.n1355 GND.n1354 9.3
R2294 GND.n1360 GND.n1359 9.3
R2295 GND.n1483 GND.n1473 9.3
R2296 GND.n1489 GND.n1469 9.3
R2297 GND.n1495 GND.n1465 9.3
R2298 GND.n1501 GND.n1461 9.3
R2299 GND.n1507 GND.n1457 9.3
R2300 GND.n1513 GND.n1453 9.3
R2301 GND.n1452 GND.n1449 9.3
R2302 GND.n1525 GND.n1442 9.3
R2303 GND.n1530 GND.n1437 9.3
R2304 GND.n1535 GND.n1432 9.3
R2305 GND.n1540 GND.n1427 9.3
R2306 GND.n1545 GND.n1420 9.3
R2307 GND.n1550 GND.n1549 9.3
R2308 GND.n1557 GND.n1394 9.3
R2309 GND.n1396 GND.n1395 9.3
R2310 GND.n1524 GND.n1523 9.3
R2311 GND.n1529 GND.n1528 9.3
R2312 GND.n1534 GND.n1533 9.3
R2313 GND.n1539 GND.n1538 9.3
R2314 GND.n1544 GND.n1543 9.3
R2315 GND.n1548 GND.n1419 9.3
R2316 GND.n1556 GND.n1555 9.3
R2317 GND.n1417 GND.n1416 9.3
R2318 GND.n1401 GND.n1398 9.3
R2319 GND.n1413 GND.n1398 9.3
R2320 GND.n1413 GND.n1412 9.3
R2321 GND.n1559 GND.n1558 9.3
R2322 GND.n1560 GND.n1559 9.3
R2323 GND.n1561 GND.n1560 9.3
R2324 GND.n1551 GND.n1418 9.3
R2325 GND.n1551 GND.n1364 9.3
R2326 GND.n1561 GND.n1364 9.3
R2327 GND.n1547 GND.n1546 9.3
R2328 GND.n1546 GND.n1389 9.3
R2329 GND.n1561 GND.n1389 9.3
R2330 GND.n1542 GND.n1541 9.3
R2331 GND.n1541 GND.n1366 9.3
R2332 GND.n1561 GND.n1366 9.3
R2333 GND.n1537 GND.n1536 9.3
R2334 GND.n1536 GND.n1387 9.3
R2335 GND.n1561 GND.n1387 9.3
R2336 GND.n1532 GND.n1531 9.3
R2337 GND.n1531 GND.n1368 9.3
R2338 GND.n1561 GND.n1368 9.3
R2339 GND.n1527 GND.n1526 9.3
R2340 GND.n1526 GND.n1385 9.3
R2341 GND.n1561 GND.n1385 9.3
R2342 GND.n1448 GND.n1447 9.3
R2343 GND.n1517 GND.n1516 9.3
R2344 GND.n1518 GND.n1517 9.3
R2345 GND.n1515 GND.n1514 9.3
R2346 GND.n1512 GND.n1510 9.3
R2347 GND.n1512 GND.n1511 9.3
R2348 GND.n1509 GND.n1508 9.3
R2349 GND.n1506 GND.n1504 9.3
R2350 GND.n1506 GND.n1505 9.3
R2351 GND.n1503 GND.n1502 9.3
R2352 GND.n1500 GND.n1498 9.3
R2353 GND.n1500 GND.n1499 9.3
R2354 GND.n1497 GND.n1496 9.3
R2355 GND.n1494 GND.n1492 9.3
R2356 GND.n1494 GND.n1493 9.3
R2357 GND.n1491 GND.n1490 9.3
R2358 GND.n1488 GND.n1486 9.3
R2359 GND.n1488 GND.n1487 9.3
R2360 GND.n1485 GND.n1484 9.3
R2361 GND.n1482 GND.n1480 9.3
R2362 GND.n1482 GND.n1481 9.3
R2363 GND.n1479 GND.n1478 9.3
R2364 GND.n1574 GND.n1573 9.3
R2365 GND.n1573 GND.n1572 9.3
R2366 GND.n2363 GND.n2362 9.3
R2367 GND.n2352 GND.n2351 9.3
R2368 GND.n2350 GND.n2349 9.3
R2369 GND.n2359 GND.n2358 9.3
R2370 GND.n2358 GND.n2357 9.3
R2371 GND.n2361 GND.n2360 9.3
R2372 GND.n2365 GND.n2364 9.3
R2373 GND.n1578 GND.n1577 9.3
R2374 GND.n1582 GND.n1581 9.3
R2375 GND.n1585 GND.n1584 9.3
R2376 GND.n1590 GND.n1589 9.3
R2377 GND.n1589 GND.n1588 9.3
R2378 GND.n1592 GND.n1591 9.3
R2379 GND.n1596 GND.n1595 9.3
R2380 GND.n1827 GND.n1826 9.3
R2381 GND.n1831 GND.n1830 9.3
R2382 GND.n1834 GND.n1833 9.3
R2383 GND.n1839 GND.n1838 9.3
R2384 GND.n1838 GND.n1837 9.3
R2385 GND.n1841 GND.n1840 9.3
R2386 GND.n1845 GND.n1844 9.3
R2387 GND.n2076 GND.n2075 9.3
R2388 GND.n2080 GND.n2079 9.3
R2389 GND.n2083 GND.n2082 9.3
R2390 GND.n2088 GND.n2087 9.3
R2391 GND.n2087 GND.n2086 9.3
R2392 GND.n2090 GND.n2089 9.3
R2393 GND.n2094 GND.n2093 9.3
R2394 GND.n2341 GND.n2340 9.3
R2395 GND.n2330 GND.n2329 9.3
R2396 GND.n2328 GND.n2327 9.3
R2397 GND.n2337 GND.n2336 9.3
R2398 GND.n2336 GND.n2335 9.3
R2399 GND.n2339 GND.n2338 9.3
R2400 GND.n2343 GND.n2342 9.3
R2401 GND.n1183 GND.n1138 9.292
R2402 GND.n2156 GND.n2155 9.233
R2403 GND.n2280 GND.n2279 9.233
R2404 GND.n2157 GND.n2156 9.233
R2405 GND.n2279 GND.n2278 9.233
R2406 GND.n1423 GND.n1365 9.233
R2407 GND.n1421 GND.n1365 9.233
R2408 GND.n74 GND.n70 9.205
R2409 GND.n495 GND.n454 9.205
R2410 GND.n840 GND.n799 9.205
R2411 GND.n2048 GND.n1858 9.147
R2412 GND.n1970 GND.n1872 9.147
R2413 GND.n2045 GND.n1858 9.147
R2414 GND.n1963 GND.n1872 9.147
R2415 GND.n1799 GND.n1609 9.147
R2416 GND.n1721 GND.n1623 9.147
R2417 GND.n1796 GND.n1609 9.147
R2418 GND.n1714 GND.n1623 9.147
R2419 GND.n30 GND.n29 9.127
R2420 GND.n620 GND.n405 9.127
R2421 GND.n621 GND.n620 9.127
R2422 GND.n965 GND.n750 9.127
R2423 GND.n966 GND.n965 9.127
R2424 GND.n2067 GND.n1883 9.126
R2425 GND.n2068 GND.n2067 9.126
R2426 GND.n1818 GND.n1634 9.126
R2427 GND.n1819 GND.n1818 9.126
R2428 GND.n1310 GND.n1300 9.126
R2429 GND.n1302 GND.n1300 9.126
R2430 GND.n2105 GND.n2104 9.126
R2431 GND.n1571 GND.n1561 9.126
R2432 GND.n1563 GND.n1561 9.126
R2433 GND.n2145 GND.n2144 9.09
R2434 GND.n2293 GND.n2292 9.09
R2435 GND.n1471 GND.n1376 9.09
R2436 GND.n1300 GND.n1085 9.07
R2437 GND.n1561 GND.n1378 9.069
R2438 GND.n219 GND.n218 9.063
R2439 GND.n218 GND.n217 9.063
R2440 GND.n578 GND.n394 9.063
R2441 GND.n598 GND.n394 9.063
R2442 GND.n923 GND.n739 9.063
R2443 GND.n943 GND.n739 9.063
R2444 GND.n620 GND.n395 9.015
R2445 GND.n965 GND.n740 9.015
R2446 GND.n2067 GND.n1857 9.014
R2447 GND.n2067 GND.n1873 9.014
R2448 GND.n1818 GND.n1608 9.014
R2449 GND.n1818 GND.n1624 9.014
R2450 GND.n1300 GND.n1083 9.014
R2451 GND.n1561 GND.n1376 9.013
R2452 GND.n1905 GND.n1857 9.006
R2453 GND.n1948 GND.n1873 9.006
R2454 GND.n1656 GND.n1608 9.006
R2455 GND.n1699 GND.n1624 9.006
R2456 GND.n1272 GND.n1083 9.006
R2457 GND.n1300 GND.n1087 8.959
R2458 GND.n1561 GND.n1380 8.957
R2459 GND.n232 GND.n231 8.923
R2460 GND.n583 GND.n395 8.923
R2461 GND.n928 GND.n740 8.923
R2462 GND.n620 GND.n392 8.907
R2463 GND.n965 GND.n737 8.907
R2464 GND.n2067 GND.n1860 8.904
R2465 GND.n2067 GND.n1870 8.904
R2466 GND.n1818 GND.n1611 8.904
R2467 GND.n1818 GND.n1621 8.904
R2468 GND.n1300 GND.n1081 8.904
R2469 GND.n1561 GND.n1374 8.902
R2470 GND.n1561 GND.n1382 8.848
R2471 GND.n2067 GND.n1863 8.797
R2472 GND.n2067 GND.n1867 8.797
R2473 GND.n1818 GND.n1614 8.797
R2474 GND.n1818 GND.n1618 8.797
R2475 GND.n1561 GND.n1372 8.794
R2476 GND.n1561 GND.n1384 8.741
R2477 GND.n620 GND.n396 7.864
R2478 GND.n620 GND.n393 7.864
R2479 GND.n965 GND.n741 7.864
R2480 GND.n965 GND.n738 7.864
R2481 GND.n2067 GND.n1874 7.853
R2482 GND.n2067 GND.n1871 7.853
R2483 GND.n2067 GND.n1868 7.853
R2484 GND.n2067 GND.n1856 7.853
R2485 GND.n2067 GND.n1859 7.853
R2486 GND.n2067 GND.n1862 7.853
R2487 GND.n1818 GND.n1625 7.853
R2488 GND.n1818 GND.n1622 7.853
R2489 GND.n1818 GND.n1619 7.853
R2490 GND.n1818 GND.n1607 7.853
R2491 GND.n1818 GND.n1610 7.853
R2492 GND.n1818 GND.n1613 7.853
R2493 GND.n2194 GND.n2193 7.504
R2494 GND.n2242 GND.n2241 7.504
R2495 GND.n1455 GND.n1383 7.504
R2496 GND.n2021 GND.n2020 7.433
R2497 GND.n1933 GND.n1932 7.433
R2498 GND.n1772 GND.n1771 7.433
R2499 GND.n1684 GND.n1683 7.433
R2500 GND.n1211 GND.n1118 7.433
R2501 GND.n1250 GND.n1097 7.433
R2502 GND.n1428 GND.n1388 7.41
R2503 GND.n1425 GND.n1388 7.41
R2504 GND.n126 GND.n125 7.364
R2505 GND.n180 GND.n179 7.364
R2506 GND.n526 GND.n433 7.364
R2507 GND.n567 GND.n413 7.364
R2508 GND.n871 GND.n778 7.364
R2509 GND.n912 GND.n758 7.364
R2510 GND.n2067 GND.n1865 6.796
R2511 GND.n2067 GND.n1884 6.796
R2512 GND.n1818 GND.n1616 6.796
R2513 GND.n1818 GND.n1635 6.796
R2514 GND.n12 GND.n8 5.647
R2515 GND.n274 GND.n270 5.647
R2516 GND.n294 GND.n290 5.647
R2517 GND.n314 GND.n310 5.647
R2518 GND.n336 GND.n332 5.647
R2519 GND.n377 GND.n370 5.647
R2520 GND.n377 GND.n368 5.647
R2521 GND.n357 GND.n350 5.647
R2522 GND.n357 GND.n348 5.647
R2523 GND.n639 GND.n632 5.647
R2524 GND.n639 GND.n630 5.647
R2525 GND.n659 GND.n652 5.647
R2526 GND.n659 GND.n650 5.647
R2527 GND.n681 GND.n674 5.647
R2528 GND.n681 GND.n672 5.647
R2529 GND.n722 GND.n715 5.647
R2530 GND.n722 GND.n713 5.647
R2531 GND.n702 GND.n695 5.647
R2532 GND.n702 GND.n693 5.647
R2533 GND.n984 GND.n977 5.647
R2534 GND.n984 GND.n975 5.647
R2535 GND.n1004 GND.n997 5.647
R2536 GND.n1004 GND.n995 5.647
R2537 GND.n1026 GND.n1019 5.647
R2538 GND.n1026 GND.n1017 5.647
R2539 GND.n1067 GND.n1060 5.647
R2540 GND.n1067 GND.n1058 5.647
R2541 GND.n1047 GND.n1040 5.647
R2542 GND.n1047 GND.n1038 5.647
R2543 GND.n1328 GND.n1321 5.647
R2544 GND.n1328 GND.n1319 5.647
R2545 GND.n1348 GND.n1341 5.647
R2546 GND.n1348 GND.n1339 5.647
R2547 GND.n2358 GND.n2354 5.647
R2548 GND.n1589 GND.n1582 5.647
R2549 GND.n1589 GND.n1580 5.647
R2550 GND.n1838 GND.n1831 5.647
R2551 GND.n1838 GND.n1829 5.647
R2552 GND.n2087 GND.n2080 5.647
R2553 GND.n2087 GND.n2078 5.647
R2554 GND.n2336 GND.n2332 5.647
R2555 GND.n2134 GND.n2132 5.628
R2556 GND.n2307 GND.n2305 5.628
R2557 GND.n1560 GND.n1391 5.628
R2558 GND.n33 GND.n32 5.619
R2559 GND.n21 GND.n20 5.619
R2560 GND.n816 GND.n815 5.619
R2561 GND.n809 GND.n804 5.619
R2562 GND.n835 GND.n834 5.619
R2563 GND.n843 GND.n795 5.619
R2564 GND.n854 GND.n853 5.619
R2565 GND.n788 GND.n783 5.619
R2566 GND.n870 GND.n869 5.619
R2567 GND.n878 GND.n773 5.619
R2568 GND.n890 GND.n769 5.619
R2569 GND.n893 GND.n892 5.619
R2570 GND.n904 GND.n903 5.619
R2571 GND.n910 GND.n909 5.619
R2572 GND.n962 GND.n961 5.619
R2573 GND.n953 GND.n952 5.619
R2574 GND.n947 GND.n925 5.619
R2575 GND.n940 GND.n930 5.619
R2576 GND.n933 GND.n932 5.619
R2577 GND.n747 GND.n746 5.619
R2578 GND.n1159 GND.n1158 5.619
R2579 GND.n1167 GND.n1147 5.619
R2580 GND.n1178 GND.n1177 5.619
R2581 GND.n1140 GND.n1135 5.619
R2582 GND.n1194 GND.n1193 5.619
R2583 GND.n1202 GND.n1126 5.619
R2584 GND.n1213 GND.n1212 5.619
R2585 GND.n1215 GND.n1115 5.619
R2586 GND.n1234 GND.n1112 5.619
R2587 GND.n1230 GND.n1113 5.619
R2588 GND.n1245 GND.n1244 5.619
R2589 GND.n1253 GND.n1252 5.619
R2590 GND.n1256 GND.n1095 5.619
R2591 GND.n1298 GND.n1297 5.619
R2592 GND.n1290 GND.n1289 5.619
R2593 GND.n1284 GND.n1274 5.619
R2594 GND.n1278 GND.n1277 5.619
R2595 GND.n1305 GND.n1301 5.619
R2596 GND.n2181 GND.n2180 5.575
R2597 GND.n2255 GND.n2254 5.575
R2598 GND.n2182 GND.n2181 5.575
R2599 GND.n2254 GND.n2253 5.575
R2600 GND.n1433 GND.n1367 5.575
R2601 GND.n1430 GND.n1367 5.575
R2602 GND.n2057 GND.n2056 5.575
R2603 GND.n1957 GND.n1956 5.575
R2604 GND.n1808 GND.n1807 5.575
R2605 GND.n1708 GND.n1707 5.575
R2606 GND.n1172 GND.n1144 5.575
R2607 GND.n471 GND.n470 5.551
R2608 GND.n464 GND.n459 5.551
R2609 GND.n490 GND.n489 5.551
R2610 GND.n498 GND.n450 5.551
R2611 GND.n509 GND.n508 5.551
R2612 GND.n443 GND.n438 5.551
R2613 GND.n525 GND.n524 5.551
R2614 GND.n533 GND.n428 5.551
R2615 GND.n545 GND.n424 5.551
R2616 GND.n548 GND.n547 5.551
R2617 GND.n559 GND.n558 5.551
R2618 GND.n565 GND.n564 5.551
R2619 GND.n617 GND.n616 5.551
R2620 GND.n608 GND.n607 5.551
R2621 GND.n602 GND.n580 5.551
R2622 GND.n595 GND.n585 5.551
R2623 GND.n588 GND.n587 5.551
R2624 GND.n402 GND.n401 5.551
R2625 GND.n60 GND.n56 5.523
R2626 GND.n246 GND.n244 5.523
R2627 GND.n483 GND.n456 5.523
R2628 GND.n592 GND.n591 5.523
R2629 GND.n828 GND.n801 5.523
R2630 GND.n937 GND.n936 5.523
R2631 GND.n2032 GND.n1861 5.523
R2632 GND.n1984 GND.n1869 5.523
R2633 GND.n2029 GND.n1861 5.523
R2634 GND.n1977 GND.n1869 5.523
R2635 GND.n1783 GND.n1612 5.523
R2636 GND.n1735 GND.n1620 5.523
R2637 GND.n1780 GND.n1612 5.523
R2638 GND.n1728 GND.n1620 5.523
R2639 GND.n1475 GND.n1378 5.488
R2640 GND.n1275 GND.n1085 5.437
R2641 GND.n1895 GND.n1894 5.421
R2642 GND.n2060 GND.n2059 5.421
R2643 GND.n1903 GND.n1901 5.421
R2644 GND.n2047 GND.n1908 5.421
R2645 GND.n2039 GND.n2038 5.421
R2646 GND.n2031 GND.n1913 5.421
R2647 GND.n2023 GND.n2022 5.421
R2648 GND.n2015 GND.n1919 5.421
R2649 GND.n2007 GND.n2006 5.421
R2650 GND.n2003 GND.n2002 5.421
R2651 GND.n1994 GND.n1927 5.421
R2652 GND.n1988 GND.n1934 5.421
R2653 GND.n1981 GND.n1937 5.421
R2654 GND.n1974 GND.n1942 5.421
R2655 GND.n1967 GND.n1945 5.421
R2656 GND.n1960 GND.n1950 5.421
R2657 GND.n1953 GND.n1952 5.421
R2658 GND.n1880 GND.n1879 5.421
R2659 GND.n1646 GND.n1645 5.421
R2660 GND.n1811 GND.n1810 5.421
R2661 GND.n1654 GND.n1652 5.421
R2662 GND.n1798 GND.n1659 5.421
R2663 GND.n1790 GND.n1789 5.421
R2664 GND.n1782 GND.n1664 5.421
R2665 GND.n1774 GND.n1773 5.421
R2666 GND.n1766 GND.n1670 5.421
R2667 GND.n1758 GND.n1757 5.421
R2668 GND.n1754 GND.n1753 5.421
R2669 GND.n1745 GND.n1678 5.421
R2670 GND.n1739 GND.n1685 5.421
R2671 GND.n1732 GND.n1688 5.421
R2672 GND.n1725 GND.n1693 5.421
R2673 GND.n1718 GND.n1696 5.421
R2674 GND.n1711 GND.n1701 5.421
R2675 GND.n1704 GND.n1703 5.421
R2676 GND.n1631 GND.n1630 5.421
R2677 GND.n2108 GND.n2107 5.358
R2678 GND.n2099 GND.n2098 5.358
R2679 GND.n1408 GND.n1406 5.358
R2680 GND.n1416 GND.n1415 5.358
R2681 GND.n1555 GND.n1554 5.358
R2682 GND.n1422 GND.n1419 5.358
R2683 GND.n1544 GND.n1426 5.358
R2684 GND.n1539 GND.n1431 5.358
R2685 GND.n1534 GND.n1436 5.358
R2686 GND.n1529 GND.n1441 5.358
R2687 GND.n1524 GND.n1446 5.358
R2688 GND.n1520 GND.n1448 5.358
R2689 GND.n1514 GND.n1454 5.358
R2690 GND.n1508 GND.n1458 5.358
R2691 GND.n1502 GND.n1462 5.358
R2692 GND.n1496 GND.n1466 5.358
R2693 GND.n1490 GND.n1470 5.358
R2694 GND.n1484 GND.n1474 5.358
R2695 GND.n1478 GND.n1477 5.358
R2696 GND.n1566 GND.n1562 5.358
R2697 GND.n155 GND.n153 5.307
R2698 GND.n155 GND.n154 5.307
R2699 GND.n891 GND.n890 5.307
R2700 GND.n892 GND.n891 5.307
R2701 GND.n1234 GND.n1233 5.307
R2702 GND.n1233 GND.n1113 5.307
R2703 GND.n546 GND.n545 5.243
R2704 GND.n547 GND.n546 5.243
R2705 GND.n2006 GND.n1924 5.12
R2706 GND.n2003 GND.n1924 5.12
R2707 GND.n1757 GND.n1675 5.12
R2708 GND.n1754 GND.n1675 5.12
R2709 GND.n2219 GND.n2217 5.06
R2710 GND.n2219 GND.n2218 5.06
R2711 GND.n1521 GND.n1446 5.06
R2712 GND.n1521 GND.n1520 5.06
R2713 GND.n323 GND.t134 4.957
R2714 GND.n1013 GND.t5 4.957
R2715 GND.n1357 GND.t146 4.957
R2716 GND.n668 GND.t3 4.954
R2717 GND.n383 GND.n366 4.894
R2718 GND.n363 GND.n346 4.894
R2719 GND.n645 GND.n628 4.894
R2720 GND.n665 GND.n648 4.894
R2721 GND.n687 GND.n670 4.894
R2722 GND.n728 GND.n711 4.894
R2723 GND.n708 GND.n691 4.894
R2724 GND.n990 GND.n973 4.894
R2725 GND.n1010 GND.n993 4.894
R2726 GND.n1032 GND.n1015 4.894
R2727 GND.n1073 GND.n1056 4.894
R2728 GND.n1053 GND.n1036 4.894
R2729 GND.n1334 GND.n1317 4.894
R2730 GND.n1354 GND.n1337 4.894
R2731 GND.n1595 GND.n1578 4.894
R2732 GND.n1844 GND.n1827 4.894
R2733 GND.n2093 GND.n2076 4.894
R2734 GND.n323 GND.t85 4.862
R2735 GND.n1013 GND.t125 4.862
R2736 GND.n1357 GND.t48 4.862
R2737 GND.n668 GND.t23 4.859
R2738 GND.n1034 GND.t18 4.832
R2739 GND.n2366 GND.t31 4.832
R2740 GND.n344 GND.t95 4.829
R2741 GND.n689 GND.t67 4.829
R2742 GND.n156 GND.n155 4.65
R2743 GND.n2220 GND.n2219 4.65
R2744 GND.n546 GND.n423 4.65
R2745 GND.n1924 GND.n1923 4.65
R2746 GND.n891 GND.n768 4.65
R2747 GND.n1675 GND.n1674 4.65
R2748 GND.n1233 GND.n1232 4.65
R2749 GND.n1522 GND.n1521 4.65
R2750 GND.n10 GND.n9 4.137
R2751 GND.n272 GND.n271 4.137
R2752 GND.n292 GND.n291 4.137
R2753 GND.n312 GND.n311 4.137
R2754 GND.n334 GND.n333 4.137
R2755 GND.n382 GND.n367 4.137
R2756 GND.n362 GND.n347 4.137
R2757 GND.n644 GND.n629 4.137
R2758 GND.n664 GND.n649 4.137
R2759 GND.n686 GND.n671 4.137
R2760 GND.n727 GND.n712 4.137
R2761 GND.n707 GND.n692 4.137
R2762 GND.n989 GND.n974 4.137
R2763 GND.n1009 GND.n994 4.137
R2764 GND.n1031 GND.n1016 4.137
R2765 GND.n1072 GND.n1057 4.137
R2766 GND.n1052 GND.n1037 4.137
R2767 GND.n1333 GND.n1318 4.137
R2768 GND.n1353 GND.n1338 4.137
R2769 GND.n2356 GND.n2355 4.137
R2770 GND.n1594 GND.n1579 4.137
R2771 GND.n1843 GND.n1828 4.137
R2772 GND.n2092 GND.n2077 4.137
R2773 GND.n2334 GND.n2333 4.137
R2774 GND.n1450 GND.n1371 3.752
R2775 GND.n1438 GND.n1386 3.729
R2776 GND.n1435 GND.n1386 3.729
R2777 GND.n1224 GND.n1116 3.716
R2778 GND.n1246 GND.n1104 3.716
R2779 GND.n140 GND.n139 3.682
R2780 GND.n166 GND.n165 3.682
R2781 GND.n540 GND.n427 3.682
R2782 GND.n557 GND.n419 3.682
R2783 GND.n885 GND.n772 3.682
R2784 GND.n902 GND.n764 3.682
R2785 GND.n48 GND.n39 3.548
R2786 GND.n822 GND.n820 3.548
R2787 GND.n1154 GND.n1150 3.548
R2788 GND.n477 GND.n475 3.545
R2789 GND.n2063 GND.n1899 3.539
R2790 GND.n1814 GND.n1650 3.539
R2791 GND.n2123 GND.n2114 3.536
R2792 GND.n1402 GND.n1401 3.536
R2793 GND.n1561 GND.n1377 3.517
R2794 GND.n260 GND.n31 3.392
R2795 GND.n970 GND.n730 3.392
R2796 GND.n1314 GND.n1075 3.392
R2797 GND.n625 GND.n385 3.389
R2798 GND.n2072 GND.n1849 3.383
R2799 GND.n1823 GND.n1600 3.383
R2800 GND.n2321 GND.n2106 3.38
R2801 GND.n1575 GND.n1358 3.38
R2802 GND.n34 GND.n33 2.497
R2803 GND.n22 GND.n21 2.497
R2804 GND.n816 GND.n811 2.497
R2805 GND.n815 GND.n808 2.497
R2806 GND.n810 GND.n809 2.497
R2807 GND.n933 GND.n732 2.497
R2808 GND.n746 GND.n733 2.497
R2809 GND.n748 GND.n747 2.497
R2810 GND.n1158 GND.n1157 2.497
R2811 GND.n1159 GND.n1149 2.497
R2812 GND.n1167 GND.n1166 2.497
R2813 GND.n1278 GND.n1077 2.497
R2814 GND.n1301 GND.n1078 2.497
R2815 GND.n1305 GND.n1304 2.497
R2816 GND.n471 GND.n466 2.467
R2817 GND.n470 GND.n463 2.467
R2818 GND.n465 GND.n464 2.467
R2819 GND.n588 GND.n387 2.467
R2820 GND.n401 GND.n388 2.467
R2821 GND.n403 GND.n402 2.467
R2822 GND.n1895 GND.n1890 2.409
R2823 GND.n1894 GND.n1888 2.409
R2824 GND.n2060 GND.n1889 2.409
R2825 GND.n1953 GND.n1851 2.409
R2826 GND.n1879 GND.n1852 2.409
R2827 GND.n1881 GND.n1880 2.409
R2828 GND.n1646 GND.n1641 2.409
R2829 GND.n1645 GND.n1639 2.409
R2830 GND.n1811 GND.n1640 2.409
R2831 GND.n1704 GND.n1602 2.409
R2832 GND.n1630 GND.n1603 2.409
R2833 GND.n1632 GND.n1631 2.409
R2834 GND.n2109 GND.n2108 2.381
R2835 GND.n2100 GND.n2099 2.381
R2836 GND.n1406 GND.n1405 2.381
R2837 GND.n1408 GND.n1407 2.381
R2838 GND.n1416 GND.n1396 2.381
R2839 GND.n1478 GND.n1360 2.381
R2840 GND.n1562 GND.n1361 2.381
R2841 GND.n1566 GND.n1565 2.381
R2842 GND.n147 GND.n138 2.341
R2843 GND.n171 GND.n162 2.341
R2844 GND.n884 GND.n883 2.341
R2845 GND.n883 GND.n774 2.341
R2846 GND.n897 GND.n767 2.341
R2847 GND.n897 GND.n763 2.341
R2848 GND.n1226 GND.n1225 2.341
R2849 GND.n1227 GND.n1226 2.341
R2850 GND.n1240 GND.n1108 2.341
R2851 GND.n1240 GND.n1105 2.341
R2852 GND.n539 GND.n538 2.313
R2853 GND.n538 GND.n429 2.313
R2854 GND.n552 GND.n422 2.313
R2855 GND.n552 GND.n418 2.313
R2856 GND.n2210 GND.n2209 2.305
R2857 GND.n2232 GND.n2228 2.305
R2858 GND.n2012 GND.n1865 2.289
R2859 GND.n1997 GND.n1884 2.289
R2860 GND.n1763 GND.n1616 2.289
R2861 GND.n1748 GND.n1635 2.289
R2862 GND.n2014 GND.n2011 2.258
R2863 GND.n2011 GND.n1920 2.258
R2864 GND.n1998 GND.n1925 2.258
R2865 GND.n1998 GND.n1995 2.258
R2866 GND.n1765 GND.n1762 2.258
R2867 GND.n1762 GND.n1671 2.258
R2868 GND.n1749 GND.n1676 2.258
R2869 GND.n1749 GND.n1746 2.258
R2870 GND.n2211 GND.n2204 2.232
R2871 GND.n2233 GND.n2226 2.232
R2872 GND.n1526 GND.n1444 2.232
R2873 GND.n1526 GND.n1525 2.232
R2874 GND.n1517 GND.n1449 2.232
R2875 GND.n1517 GND.n1451 2.232
R2876 GND.n54 GND.n53 2.185
R2877 GND.n241 GND.n240 2.185
R2878 GND.n829 GND.n804 2.185
R2879 GND.n834 GND.n802 2.185
R2880 GND.n940 GND.n939 2.185
R2881 GND.n932 GND.n931 2.185
R2882 GND.n1171 GND.n1147 2.185
R2883 GND.n1178 GND.n1143 2.185
R2884 GND.n1284 GND.n1283 2.185
R2885 GND.n1277 GND.n1276 2.185
R2886 GND.n484 GND.n459 2.159
R2887 GND.n489 GND.n457 2.159
R2888 GND.n595 GND.n594 2.159
R2889 GND.n587 GND.n586 2.159
R2890 GND.n2059 GND.n2058 2.108
R2891 GND.n2054 GND.n1901 2.108
R2892 GND.n1960 GND.n1959 2.108
R2893 GND.n1952 GND.n1951 2.108
R2894 GND.n1810 GND.n1809 2.108
R2895 GND.n1805 GND.n1652 2.108
R2896 GND.n1711 GND.n1710 2.108
R2897 GND.n1703 GND.n1702 2.108
R2898 GND.n2129 GND.n2128 2.083
R2899 GND.n2302 GND.n2301 2.083
R2900 GND.n1415 GND.n1393 2.083
R2901 GND.n1555 GND.n1394 2.083
R2902 GND.n1484 GND.n1483 2.083
R2903 GND.n1477 GND.n1476 2.083
R2904 GND.n131 GND.n124 2.029
R2905 GND.n185 GND.n178 2.029
R2906 GND.n876 GND.n776 2.029
R2907 GND.n877 GND.n876 2.029
R2908 GND.n905 GND.n761 2.029
R2909 GND.n911 GND.n761 2.029
R2910 GND.n1219 GND.n1119 2.029
R2911 GND.n1219 GND.n1120 2.029
R2912 GND.n1106 GND.n1101 2.029
R2913 GND.n1251 GND.n1101 2.029
R2914 GND.n531 GND.n431 2.004
R2915 GND.n532 GND.n531 2.004
R2916 GND.n560 GND.n416 2.004
R2917 GND.n566 GND.n416 2.004
R2918 GND.n2019 GND.n2018 1.957
R2919 GND.n2018 GND.n1918 1.957
R2920 GND.n1991 GND.n1928 1.957
R2921 GND.n1991 GND.n1929 1.957
R2922 GND.n1770 GND.n1769 1.957
R2923 GND.n1769 GND.n1669 1.957
R2924 GND.n1742 GND.n1679 1.957
R2925 GND.n1742 GND.n1680 1.957
R2926 GND.n2197 GND.n2192 1.934
R2927 GND.n2245 GND.n2240 1.934
R2928 GND.n1531 GND.n1439 1.934
R2929 GND.n1531 GND.n1530 1.934
R2930 GND.n1513 GND.n1512 1.934
R2931 GND.n1512 GND.n1456 1.934
R2932 GND.n2121 GND.n2117 1.876
R2933 GND.n1413 GND.n1397 1.876
R2934 GND.n68 GND.n67 1.873
R2935 GND.n229 GND.n228 1.873
R2936 GND.n835 GND.n797 1.873
R2937 GND.n843 GND.n842 1.873
R2938 GND.n947 GND.n946 1.873
R2939 GND.n930 GND.n926 1.873
R2940 GND.n1177 GND.n1139 1.873
R2941 GND.n1141 GND.n1140 1.873
R2942 GND.n1289 GND.n1288 1.873
R2943 GND.n1274 GND.n1273 1.873
R2944 GND.n2206 GND.n2205 1.871
R2945 GND.n2231 GND.n2230 1.871
R2946 GND.n2207 GND.n2206 1.871
R2947 GND.n2230 GND.n2229 1.871
R2948 GND.n1443 GND.n1369 1.871
R2949 GND.n1440 GND.n1369 1.871
R2950 GND.n2065 GND.n1886 1.858
R2951 GND.n1816 GND.n1637 1.858
R2952 GND.n1164 GND.n1151 1.858
R2953 GND.n2016 GND.n1864 1.853
R2954 GND.n1996 GND.n1866 1.853
R2955 GND.n2013 GND.n1864 1.853
R2956 GND.n1993 GND.n1866 1.853
R2957 GND.n1767 GND.n1615 1.853
R2958 GND.n1747 GND.n1617 1.853
R2959 GND.n1764 GND.n1615 1.853
R2960 GND.n1744 GND.n1617 1.853
R2961 GND.n490 GND.n452 1.85
R2962 GND.n498 GND.n497 1.85
R2963 GND.n602 GND.n601 1.85
R2964 GND.n585 GND.n581 1.85
R2965 GND.n2105 GND.n2103 1.841
R2966 GND.n2317 GND.n2316 1.841
R2967 GND.n1571 GND.n1570 1.841
R2968 GND.n1564 GND.n1563 1.841
R2969 GND.n46 GND.n42 1.841
R2970 GND.n479 GND.n462 1.841
R2971 GND.n824 GND.n807 1.841
R2972 GND.n1883 GND.n1882 1.824
R2973 GND.n2068 GND.n1854 1.824
R2974 GND.n1634 GND.n1633 1.824
R2975 GND.n1819 GND.n1605 1.824
R2976 GND.n1310 GND.n1309 1.824
R2977 GND.n1303 GND.n1302 1.824
R2978 GND.n30 GND.n25 1.807
R2979 GND.n256 GND.n255 1.807
R2980 GND.n405 GND.n404 1.807
R2981 GND.n621 GND.n390 1.807
R2982 GND.n750 GND.n749 1.807
R2983 GND.n966 GND.n735 1.807
R2984 GND.n1906 GND.n1903 1.807
R2985 GND.n1908 GND.n1907 1.807
R2986 GND.n1967 GND.n1966 1.807
R2987 GND.n1950 GND.n1946 1.807
R2988 GND.n1657 GND.n1654 1.807
R2989 GND.n1659 GND.n1658 1.807
R2990 GND.n1718 GND.n1717 1.807
R2991 GND.n1701 GND.n1697 1.807
R2992 GND.n2142 GND.n2141 1.786
R2993 GND.n2290 GND.n2289 1.786
R2994 GND.n1554 GND.n1553 1.786
R2995 GND.n1550 GND.n1419 1.786
R2996 GND.n1490 GND.n1489 1.786
R2997 GND.n1474 GND.n1472 1.786
R2998 GND.n2113 GND.n2111 1.759
R2999 GND.n1404 GND.n1403 1.759
R3000 GND.n1898 GND.n1891 1.742
R3001 GND.n1649 GND.n1642 1.742
R3002 GND.n1156 GND.n1155 1.742
R3003 GND.n38 GND.n36 1.727
R3004 GND.n474 GND.n467 1.727
R3005 GND.n819 GND.n812 1.727
R3006 GND.n117 GND.n110 1.717
R3007 GND.n197 GND.n192 1.717
R3008 GND.n865 GND.n864 1.717
R3009 GND.n865 GND.n781 1.717
R3010 GND.n917 GND.n757 1.717
R3011 GND.n917 GND.n754 1.717
R3012 GND.n1206 GND.n1205 1.717
R3013 GND.n1205 GND.n1122 1.717
R3014 GND.n1259 GND.n1098 1.717
R3015 GND.n1259 GND.n1099 1.717
R3016 GND.n520 GND.n519 1.696
R3017 GND.n520 GND.n436 1.696
R3018 GND.n572 GND.n412 1.696
R3019 GND.n572 GND.n409 1.696
R3020 GND.n2030 GND.n2027 1.656
R3021 GND.n2027 GND.n1914 1.656
R3022 GND.n1987 GND.n1986 1.656
R3023 GND.n1986 GND.n1935 1.656
R3024 GND.n1781 GND.n1778 1.656
R3025 GND.n1778 GND.n1665 1.656
R3026 GND.n1738 GND.n1737 1.656
R3027 GND.n1737 GND.n1686 1.656
R3028 GND.n2185 GND.n2179 1.637
R3029 GND.n2258 GND.n2252 1.637
R3030 GND.n1536 GND.n1434 1.637
R3031 GND.n1536 GND.n1535 1.637
R3032 GND.n1507 GND.n1506 1.637
R3033 GND.n1506 GND.n1460 1.637
R3034 GND.n266 GND.n264 1.57
R3035 GND.n286 GND.n284 1.57
R3036 GND.n306 GND.n304 1.57
R3037 GND.n328 GND.n326 1.57
R3038 GND.n352 GND.n351 1.57
R3039 GND.n634 GND.n633 1.57
R3040 GND.n654 GND.n653 1.57
R3041 GND.n676 GND.n675 1.57
R3042 GND.n697 GND.n696 1.57
R3043 GND.n979 GND.n978 1.57
R3044 GND.n999 GND.n998 1.57
R3045 GND.n1021 GND.n1020 1.57
R3046 GND.n1042 GND.n1041 1.57
R3047 GND.n1323 GND.n1322 1.57
R3048 GND.n1343 GND.n1342 1.57
R3049 GND.n2350 GND.n2348 1.57
R3050 GND.n1584 GND.n1583 1.57
R3051 GND.n1833 GND.n1832 1.57
R3052 GND.n2082 GND.n2081 1.57
R3053 GND.n2328 GND.n2326 1.57
R3054 GND.n82 GND.n81 1.56
R3055 GND.n216 GND.n215 1.56
R3056 GND.n847 GND.n795 1.56
R3057 GND.n854 GND.n791 1.56
R3058 GND.n952 GND.n951 1.56
R3059 GND.n925 GND.n924 1.56
R3060 GND.n1188 GND.n1135 1.56
R3061 GND.n1193 GND.n1133 1.56
R3062 GND.n1297 GND.n1091 1.56
R3063 GND.n1292 GND.n1290 1.56
R3064 GND.n4 GND.n2 1.553
R3065 GND.n717 GND.n716 1.553
R3066 GND.n1062 GND.n1061 1.553
R3067 GND.n372 GND.n371 1.549
R3068 GND.n502 GND.n450 1.542
R3069 GND.n509 GND.n446 1.542
R3070 GND.n607 GND.n606 1.542
R3071 GND.n580 GND.n579 1.542
R3072 GND.n380 GND.n366 1.505
R3073 GND.n360 GND.n346 1.505
R3074 GND.n642 GND.n628 1.505
R3075 GND.n662 GND.n648 1.505
R3076 GND.n2047 GND.n2046 1.505
R3077 GND.n2039 GND.n1909 1.505
R3078 GND.n1974 GND.n1973 1.505
R3079 GND.n1945 GND.n1943 1.505
R3080 GND.n684 GND.n670 1.505
R3081 GND.n725 GND.n711 1.505
R3082 GND.n705 GND.n691 1.505
R3083 GND.n987 GND.n973 1.505
R3084 GND.n1007 GND.n993 1.505
R3085 GND.n1798 GND.n1797 1.505
R3086 GND.n1790 GND.n1660 1.505
R3087 GND.n1725 GND.n1724 1.505
R3088 GND.n1696 GND.n1694 1.505
R3089 GND.n1029 GND.n1015 1.505
R3090 GND.n1070 GND.n1056 1.505
R3091 GND.n1050 GND.n1036 1.505
R3092 GND.n1331 GND.n1317 1.505
R3093 GND.n1351 GND.n1337 1.505
R3094 GND.n1592 GND.n1578 1.505
R3095 GND.n1841 GND.n1827 1.505
R3096 GND.n2090 GND.n2076 1.505
R3097 GND.n2154 GND.n2153 1.488
R3098 GND.n2277 GND.n2276 1.488
R3099 GND.n1424 GND.n1422 1.488
R3100 GND.n1545 GND.n1544 1.488
R3101 GND.n1496 GND.n1495 1.488
R3102 GND.n1470 GND.n1468 1.488
R3103 GND.n103 GND.n96 1.404
R3104 GND.n209 GND.n204 1.404
R3105 GND.n858 GND.n787 1.404
R3106 GND.n858 GND.n789 1.404
R3107 GND.n957 GND.n755 1.404
R3108 GND.n957 GND.n956 1.404
R3109 GND.n1200 GND.n1128 1.404
R3110 GND.n1201 GND.n1200 1.404
R3111 GND.n1266 GND.n1093 1.404
R3112 GND.n1266 GND.n1090 1.404
R3113 GND.n513 GND.n442 1.387
R3114 GND.n513 GND.n444 1.387
R3115 GND.n612 GND.n410 1.387
R3116 GND.n612 GND.n611 1.387
R3117 GND.n2035 GND.n2034 1.355
R3118 GND.n2034 GND.n1912 1.355
R3119 GND.n1980 GND.n1979 1.355
R3120 GND.n1979 GND.n1938 1.355
R3121 GND.n1786 GND.n1785 1.355
R3122 GND.n1785 GND.n1663 1.355
R3123 GND.n1731 GND.n1730 1.355
R3124 GND.n1730 GND.n1689 1.355
R3125 GND.n2172 GND.n2167 1.339
R3126 GND.n2270 GND.n2265 1.339
R3127 GND.n1541 GND.n1429 1.339
R3128 GND.n1541 GND.n1540 1.339
R3129 GND.n1501 GND.n1500 1.339
R3130 GND.n1500 GND.n1464 1.339
R3131 GND.n2134 GND.n2133 1.334
R3132 GND.n2159 GND.n2158 1.334
R3133 GND.n2184 GND.n2183 1.334
R3134 GND.n2257 GND.n2256 1.334
R3135 GND.n2282 GND.n2281 1.334
R3136 GND.n2307 GND.n2306 1.334
R3137 GND.n2056 GND.n1856 1.323
R3138 GND.n2044 GND.n1859 1.323
R3139 GND.n2028 GND.n1862 1.323
R3140 GND.n1985 GND.n1868 1.323
R3141 GND.n1971 GND.n1871 1.323
R3142 GND.n1957 GND.n1874 1.323
R3143 GND.n1807 GND.n1607 1.323
R3144 GND.n1795 GND.n1610 1.323
R3145 GND.n1779 GND.n1613 1.323
R3146 GND.n1736 GND.n1619 1.323
R3147 GND.n1722 GND.n1622 1.323
R3148 GND.n1708 GND.n1625 1.323
R3149 GND.n221 GND.n220 1.312
R3150 GND.n246 GND.n245 1.312
R3151 GND.n577 GND.n393 1.312
R3152 GND.n592 GND.n396 1.312
R3153 GND.n922 GND.n738 1.312
R3154 GND.n937 GND.n741 1.312
R3155 GND.n96 GND.n95 1.248
R3156 GND.n204 GND.n203 1.248
R3157 GND.n853 GND.n787 1.248
R3158 GND.n789 GND.n788 1.248
R3159 GND.n961 GND.n755 1.248
R3160 GND.n956 GND.n953 1.248
R3161 GND.n1194 GND.n1128 1.248
R3162 GND.n1202 GND.n1201 1.248
R3163 GND.n1256 GND.n1093 1.248
R3164 GND.n1298 GND.n1090 1.248
R3165 GND.n508 GND.n442 1.233
R3166 GND.n444 GND.n443 1.233
R3167 GND.n616 GND.n410 1.233
R3168 GND.n611 GND.n608 1.233
R3169 GND.n2038 GND.n2035 1.204
R3170 GND.n1913 GND.n1912 1.204
R3171 GND.n1981 GND.n1980 1.204
R3172 GND.n1942 GND.n1938 1.204
R3173 GND.n1789 GND.n1786 1.204
R3174 GND.n1664 GND.n1663 1.204
R3175 GND.n1732 GND.n1731 1.204
R3176 GND.n1693 GND.n1689 1.204
R3177 GND.n2167 GND.n2166 1.19
R3178 GND.n2265 GND.n2264 1.19
R3179 GND.n1429 GND.n1426 1.19
R3180 GND.n1540 GND.n1539 1.19
R3181 GND.n1502 GND.n1501 1.19
R3182 GND.n1466 GND.n1464 1.19
R3183 GND.n89 GND.n82 1.092
R3184 GND.n222 GND.n216 1.092
R3185 GND.n847 GND.n846 1.092
R3186 GND.n846 GND.n791 1.092
R3187 GND.n951 GND.n920 1.092
R3188 GND.n924 GND.n920 1.092
R3189 GND.n1189 GND.n1188 1.092
R3190 GND.n1189 GND.n1133 1.092
R3191 GND.n1293 GND.n1091 1.092
R3192 GND.n1293 GND.n1292 1.092
R3193 GND.n502 GND.n501 1.079
R3194 GND.n501 GND.n446 1.079
R3195 GND.n606 GND.n575 1.079
R3196 GND.n579 GND.n575 1.079
R3197 GND.n2046 GND.n2043 1.054
R3198 GND.n2043 GND.n1909 1.054
R3199 GND.n1973 GND.n1972 1.054
R3200 GND.n1972 GND.n1943 1.054
R3201 GND.n1797 GND.n1794 1.054
R3202 GND.n1794 GND.n1660 1.054
R3203 GND.n1724 GND.n1723 1.054
R3204 GND.n1723 GND.n1694 1.054
R3205 GND.n2160 GND.n2154 1.041
R3206 GND.n2283 GND.n2277 1.041
R3207 GND.n1546 GND.n1424 1.041
R3208 GND.n1546 GND.n1545 1.041
R3209 GND.n1495 GND.n1494 1.041
R3210 GND.n1494 GND.n1468 1.041
R3211 GND.n110 GND.n109 0.936
R3212 GND.n192 GND.n191 0.936
R3213 GND.n864 GND.n783 0.936
R3214 GND.n869 GND.n781 0.936
R3215 GND.n909 GND.n757 0.936
R3216 GND.n962 GND.n754 0.936
R3217 GND.n1206 GND.n1126 0.936
R3218 GND.n1213 GND.n1122 0.936
R3219 GND.n1253 GND.n1098 0.936
R3220 GND.n1099 GND.n1095 0.936
R3221 GND.n519 GND.n438 0.925
R3222 GND.n524 GND.n436 0.925
R3223 GND.n564 GND.n412 0.925
R3224 GND.n617 GND.n409 0.925
R3225 GND.n2031 GND.n2030 0.903
R3226 GND.n2023 GND.n1914 0.903
R3227 GND.n1988 GND.n1987 0.903
R3228 GND.n1937 GND.n1935 0.903
R3229 GND.n1782 GND.n1781 0.903
R3230 GND.n1774 GND.n1665 0.903
R3231 GND.n1739 GND.n1738 0.903
R3232 GND.n1688 GND.n1686 0.903
R3233 GND.n2179 GND.n2178 0.893
R3234 GND.n2252 GND.n2251 0.893
R3235 GND.n1434 GND.n1431 0.893
R3236 GND.n1535 GND.n1534 0.893
R3237 GND.n1508 GND.n1507 0.893
R3238 GND.n1462 GND.n1460 0.893
R3239 GND.n75 GND.n68 0.78
R3240 GND.n234 GND.n229 0.78
R3241 GND.n841 GND.n797 0.78
R3242 GND.n842 GND.n841 0.78
R3243 GND.n946 GND.n945 0.78
R3244 GND.n945 GND.n926 0.78
R3245 GND.n1182 GND.n1139 0.78
R3246 GND.n1182 GND.n1141 0.78
R3247 GND.n1288 GND.n1270 0.78
R3248 GND.n1273 GND.n1270 0.78
R3249 GND.n496 GND.n452 0.771
R3250 GND.n497 GND.n496 0.771
R3251 GND.n601 GND.n600 0.771
R3252 GND.n600 GND.n581 0.771
R3253 GND.n8 GND.n7 0.752
R3254 GND.n270 GND.n269 0.752
R3255 GND.n290 GND.n289 0.752
R3256 GND.n310 GND.n309 0.752
R3257 GND.n332 GND.n331 0.752
R3258 GND.n373 GND.n370 0.752
R3259 GND.n381 GND.n368 0.752
R3260 GND.n353 GND.n350 0.752
R3261 GND.n361 GND.n348 0.752
R3262 GND.n635 GND.n632 0.752
R3263 GND.n643 GND.n630 0.752
R3264 GND.n655 GND.n652 0.752
R3265 GND.n663 GND.n650 0.752
R3266 GND.n2050 GND.n1906 0.752
R3267 GND.n2050 GND.n1907 0.752
R3268 GND.n1966 GND.n1965 0.752
R3269 GND.n1965 GND.n1946 0.752
R3270 GND.n677 GND.n674 0.752
R3271 GND.n685 GND.n672 0.752
R3272 GND.n718 GND.n715 0.752
R3273 GND.n726 GND.n713 0.752
R3274 GND.n698 GND.n695 0.752
R3275 GND.n706 GND.n693 0.752
R3276 GND.n980 GND.n977 0.752
R3277 GND.n988 GND.n975 0.752
R3278 GND.n1000 GND.n997 0.752
R3279 GND.n1008 GND.n995 0.752
R3280 GND.n1801 GND.n1657 0.752
R3281 GND.n1801 GND.n1658 0.752
R3282 GND.n1717 GND.n1716 0.752
R3283 GND.n1716 GND.n1697 0.752
R3284 GND.n1022 GND.n1019 0.752
R3285 GND.n1030 GND.n1017 0.752
R3286 GND.n1063 GND.n1060 0.752
R3287 GND.n1071 GND.n1058 0.752
R3288 GND.n1043 GND.n1040 0.752
R3289 GND.n1051 GND.n1038 0.752
R3290 GND.n1324 GND.n1321 0.752
R3291 GND.n1332 GND.n1319 0.752
R3292 GND.n1344 GND.n1341 0.752
R3293 GND.n1352 GND.n1339 0.752
R3294 GND.n2354 GND.n2353 0.752
R3295 GND.n1585 GND.n1582 0.752
R3296 GND.n1593 GND.n1580 0.752
R3297 GND.n1834 GND.n1831 0.752
R3298 GND.n1842 GND.n1829 0.752
R3299 GND.n2083 GND.n2080 0.752
R3300 GND.n2091 GND.n2078 0.752
R3301 GND.n2332 GND.n2331 0.752
R3302 GND.n2147 GND.n2142 0.744
R3303 GND.n2295 GND.n2290 0.744
R3304 GND.n1553 GND.n1551 0.744
R3305 GND.n1551 GND.n1550 0.744
R3306 GND.n1489 GND.n1488 0.744
R3307 GND.n1488 GND.n1472 0.744
R3308 GND.n124 GND.n123 0.624
R3309 GND.n178 GND.n177 0.624
R3310 GND.n870 GND.n776 0.624
R3311 GND.n878 GND.n877 0.624
R3312 GND.n905 GND.n904 0.624
R3313 GND.n911 GND.n910 0.624
R3314 GND.n1212 GND.n1119 0.624
R3315 GND.n1215 GND.n1120 0.624
R3316 GND.n1244 GND.n1106 0.624
R3317 GND.n1252 GND.n1251 0.624
R3318 GND.n525 GND.n431 0.616
R3319 GND.n533 GND.n532 0.616
R3320 GND.n560 GND.n559 0.616
R3321 GND.n566 GND.n565 0.616
R3322 GND.n2022 GND.n2019 0.602
R3323 GND.n1919 GND.n1918 0.602
R3324 GND.n1928 GND.n1927 0.602
R3325 GND.n1934 GND.n1929 0.602
R3326 GND.n1773 GND.n1770 0.602
R3327 GND.n1670 GND.n1669 0.602
R3328 GND.n1679 GND.n1678 0.602
R3329 GND.n1685 GND.n1680 0.602
R3330 GND.n2192 GND.n2191 0.595
R3331 GND.n2240 GND.n2239 0.595
R3332 GND.n1439 GND.n1436 0.595
R3333 GND.n1530 GND.n1529 0.595
R3334 GND.n1514 GND.n1513 0.595
R3335 GND.n1458 GND.n1456 0.595
R3336 GND.n61 GND.n54 0.468
R3337 GND.n247 GND.n241 0.468
R3338 GND.n830 GND.n829 0.468
R3339 GND.n830 GND.n802 0.468
R3340 GND.n939 GND.n938 0.468
R3341 GND.n938 GND.n931 0.468
R3342 GND.n1171 GND.n1170 0.468
R3343 GND.n1170 GND.n1143 0.468
R3344 GND.n1283 GND.n1282 0.468
R3345 GND.n1282 GND.n1276 0.468
R3346 GND.n485 GND.n484 0.462
R3347 GND.n485 GND.n457 0.462
R3348 GND.n594 GND.n593 0.462
R3349 GND.n593 GND.n586 0.462
R3350 GND.n2058 GND.n2055 0.451
R3351 GND.n2055 GND.n2054 0.451
R3352 GND.n1959 GND.n1958 0.451
R3353 GND.n1958 GND.n1951 0.451
R3354 GND.n1809 GND.n1806 0.451
R3355 GND.n1806 GND.n1805 0.451
R3356 GND.n1710 GND.n1709 0.451
R3357 GND.n1709 GND.n1702 0.451
R3358 GND.n2345 GND.n281 0.446
R3359 GND.n2135 GND.n2129 0.446
R3360 GND.n2308 GND.n2302 0.446
R3361 GND.n1559 GND.n1393 0.446
R3362 GND.n1559 GND.n1394 0.446
R3363 GND.n1483 GND.n1482 0.446
R3364 GND.n1482 GND.n1476 0.446
R3365 GND.n1847 GND.n709 0.446
R3366 GND.n1598 GND.n1054 0.446
R3367 GND.n2096 GND.n364 0.444
R3368 GND.n1518 GND.n1384 0.421
R3369 GND.n1597 GND.n1596 0.42
R3370 GND.n1846 GND.n1845 0.42
R3371 GND.n2095 GND.n2094 0.42
R3372 GND.n2344 GND.n2343 0.42
R3373 GND.n322 GND.n321 0.415
R3374 GND.n1012 GND.n1011 0.415
R3375 GND.n1356 GND.n1355 0.415
R3376 GND.n667 GND.n666 0.412
R3377 GND.n1576 GND.n1575 0.38
R3378 GND.n322 GND.n301 0.375
R3379 GND.n667 GND.n646 0.375
R3380 GND.n1012 GND.n991 0.375
R3381 GND.n1356 GND.n1335 0.375
R3382 GND.n2244 GND.n2243 0.367
R3383 GND.n2196 GND.n2195 0.367
R3384 GND.n1511 GND.n1372 0.367
R3385 GND.n344 GND.n343 0.364
R3386 GND.n1034 GND.n1033 0.364
R3387 GND.n2366 GND.n2365 0.364
R3388 GND.n1992 GND.n1867 0.364
R3389 GND.n2017 GND.n1863 0.364
R3390 GND.n1743 GND.n1618 0.364
R3391 GND.n1768 GND.n1614 0.364
R3392 GND.n689 GND.n688 0.361
R3393 GND.n2073 GND.n2072 0.331
R3394 GND.n2322 GND.n2321 0.331
R3395 GND.n1824 GND.n1823 0.328
R3396 GND.n261 GND.n19 0.318
R3397 GND.n971 GND.n729 0.318
R3398 GND.n1315 GND.n1074 0.318
R3399 GND.n1505 GND.n1382 0.313
R3400 GND.n138 GND.n137 0.312
R3401 GND.n162 GND.n161 0.312
R3402 GND.n884 GND.n773 0.312
R3403 GND.n774 GND.n769 0.312
R3404 GND.n893 GND.n767 0.312
R3405 GND.n903 GND.n763 0.312
R3406 GND.n1225 GND.n1115 0.312
R3407 GND.n1227 GND.n1112 0.312
R3408 GND.n1230 GND.n1108 0.312
R3409 GND.n1245 GND.n1105 0.312
R3410 GND.n626 GND.n384 0.309
R3411 GND.n539 GND.n428 0.308
R3412 GND.n429 GND.n424 0.308
R3413 GND.n548 GND.n422 0.308
R3414 GND.n558 GND.n418 0.308
R3415 GND.n2015 GND.n2014 0.301
R3416 GND.n2007 GND.n1920 0.301
R3417 GND.n2002 GND.n1925 0.301
R3418 GND.n1995 GND.n1994 0.301
R3419 GND.n1766 GND.n1765 0.301
R3420 GND.n1758 GND.n1671 0.301
R3421 GND.n1753 GND.n1676 0.301
R3422 GND.n1746 GND.n1745 0.301
R3423 GND.n2204 GND.n2203 0.297
R3424 GND.n2226 GND.n2225 0.297
R3425 GND.n1444 GND.n1441 0.297
R3426 GND.n1525 GND.n1524 0.297
R3427 GND.n1449 GND.n1448 0.297
R3428 GND.n1454 GND.n1451 0.297
R3429 GND.n971 GND.n970 0.262
R3430 GND.n1315 GND.n1314 0.262
R3431 GND.n261 GND.n260 0.26
R3432 GND.n626 GND.n625 0.26
R3433 GND.n2269 GND.n2268 0.257
R3434 GND.n2171 GND.n2170 0.257
R3435 GND.n1499 GND.n1374 0.257
R3436 GND.n1978 GND.n1870 0.255
R3437 GND.n2033 GND.n1860 0.255
R3438 GND.n1729 GND.n1621 0.255
R3439 GND.n1784 GND.n1611 0.255
R3440 GND.n1265 GND.n1081 0.255
R3441 GND.n208 GND.n207 0.253
R3442 GND.n408 GND.n392 0.253
R3443 GND.n753 GND.n737 0.253
R3444 GND.n1493 GND.n1380 0.202
R3445 GND.n1089 GND.n1087 0.2
R3446 GND.n2321 GND.n2320 0.156
R3447 GND.n1575 GND.n1574 0.156
R3448 GND.n2072 GND.n2071 0.156
R3449 GND.n1823 GND.n1822 0.156
R3450 GND.n625 GND.n624 0.156
R3451 GND.n260 GND.n259 0.156
R3452 GND.n970 GND.n969 0.156
R3453 GND.n1314 GND.n1313 0.156
R3454 GND.n39 GND.n34 0.156
R3455 GND.n47 GND.n40 0.156
R3456 GND.n258 GND.n253 0.156
R3457 GND.n31 GND.n22 0.156
R3458 GND.n820 GND.n811 0.156
R3459 GND.n823 GND.n808 0.156
R3460 GND.n823 GND.n810 0.156
R3461 GND.n968 GND.n732 0.156
R3462 GND.n968 GND.n733 0.156
R3463 GND.n748 GND.n730 0.156
R3464 GND.n1157 GND.n1154 0.156
R3465 GND.n1165 GND.n1149 0.156
R3466 GND.n1166 GND.n1165 0.156
R3467 GND.n1312 GND.n1077 0.156
R3468 GND.n1312 GND.n1078 0.156
R3469 GND.n1304 GND.n1075 0.156
R3470 GND.n475 GND.n466 0.154
R3471 GND.n478 GND.n463 0.154
R3472 GND.n478 GND.n465 0.154
R3473 GND.n623 GND.n387 0.154
R3474 GND.n623 GND.n388 0.154
R3475 GND.n403 GND.n385 0.154
R3476 GND.n1899 GND.n1890 0.15
R3477 GND.n2064 GND.n1888 0.15
R3478 GND.n2064 GND.n1889 0.15
R3479 GND.n2070 GND.n1851 0.15
R3480 GND.n2070 GND.n1852 0.15
R3481 GND.n1881 GND.n1849 0.15
R3482 GND.n1650 GND.n1641 0.15
R3483 GND.n1815 GND.n1639 0.15
R3484 GND.n1815 GND.n1640 0.15
R3485 GND.n1821 GND.n1602 0.15
R3486 GND.n1821 GND.n1603 0.15
R3487 GND.n1632 GND.n1600 0.15
R3488 GND.n2114 GND.n2109 0.148
R3489 GND.n2122 GND.n2115 0.148
R3490 GND.n2319 GND.n2314 0.148
R3491 GND.n2106 GND.n2100 0.148
R3492 GND.n1405 GND.n1402 0.148
R3493 GND.n1407 GND.n1398 0.148
R3494 GND.n1398 GND.n1396 0.148
R3495 GND.n1573 GND.n1360 0.148
R3496 GND.n1573 GND.n1361 0.148
R3497 GND.n1565 GND.n1358 0.148
R3498 GND.n2294 GND.n2293 0.145
R3499 GND.n2146 GND.n2145 0.145
R3500 GND.n1487 GND.n1376 0.145
R3501 GND.n156 GND.n152 0.145
R3502 GND.n158 GND.n156 0.145
R3503 GND.n2220 GND.n2216 0.145
R3504 GND.n2222 GND.n2220 0.145
R3505 GND.n535 GND.n423 0.145
R3506 GND.n549 GND.n423 0.145
R3507 GND.n2008 GND.n1923 0.145
R3508 GND.n2001 GND.n1923 0.145
R3509 GND.n880 GND.n768 0.145
R3510 GND.n894 GND.n768 0.145
R3511 GND.n1759 GND.n1674 0.145
R3512 GND.n1752 GND.n1674 0.145
R3513 GND.n1232 GND.n1229 0.145
R3514 GND.n1232 GND.n1231 0.145
R3515 GND.n1523 GND.n1522 0.145
R3516 GND.n1522 GND.n1447 0.145
R3517 GND.n277 GND.n275 0.144
R3518 GND.n297 GND.n295 0.144
R3519 GND.n317 GND.n315 0.144
R3520 GND.n339 GND.n337 0.144
R3521 GND.n359 GND.n358 0.144
R3522 GND.n641 GND.n640 0.144
R3523 GND.n661 GND.n660 0.144
R3524 GND.n683 GND.n682 0.144
R3525 GND.n704 GND.n703 0.144
R3526 GND.n986 GND.n985 0.144
R3527 GND.n1006 GND.n1005 0.144
R3528 GND.n1028 GND.n1027 0.144
R3529 GND.n1049 GND.n1048 0.144
R3530 GND.n1330 GND.n1329 0.144
R3531 GND.n1350 GND.n1349 0.144
R3532 GND.n2361 GND.n2359 0.144
R3533 GND.n1591 GND.n1590 0.144
R3534 GND.n1840 GND.n1839 0.144
R3535 GND.n2089 GND.n2088 0.144
R3536 GND.n2339 GND.n2337 0.144
R3537 GND.n1964 GND.n1873 0.144
R3538 GND.n2049 GND.n1857 0.144
R3539 GND.n1715 GND.n1624 0.144
R3540 GND.n1800 GND.n1608 0.144
R3541 GND.n1269 GND.n1083 0.144
R3542 GND.n233 GND.n232 0.142
R3543 GND.n599 GND.n395 0.142
R3544 GND.n944 GND.n740 0.142
R3545 GND.n15 GND.n13 0.132
R3546 GND.n724 GND.n723 0.132
R3547 GND.n1069 GND.n1068 0.132
R3548 GND.n379 GND.n378 0.129
R3549 GND.n62 GND.n52 0.11
R3550 GND.n76 GND.n66 0.11
R3551 GND.n90 GND.n80 0.11
R3552 GND.n104 GND.n94 0.11
R3553 GND.n118 GND.n108 0.11
R3554 GND.n132 GND.n122 0.11
R3555 GND.n148 GND.n136 0.11
R3556 GND.n174 GND.n172 0.11
R3557 GND.n188 GND.n186 0.11
R3558 GND.n200 GND.n198 0.11
R3559 GND.n212 GND.n210 0.11
R3560 GND.n225 GND.n223 0.11
R3561 GND.n237 GND.n235 0.11
R3562 GND.n250 GND.n248 0.11
R3563 GND.n2136 GND.n2127 0.11
R3564 GND.n2148 GND.n2140 0.11
R3565 GND.n2161 GND.n2152 0.11
R3566 GND.n2173 GND.n2165 0.11
R3567 GND.n2186 GND.n2177 0.11
R3568 GND.n2198 GND.n2190 0.11
R3569 GND.n2212 GND.n2202 0.11
R3570 GND.n2236 GND.n2234 0.11
R3571 GND.n2248 GND.n2246 0.11
R3572 GND.n2261 GND.n2259 0.11
R3573 GND.n2273 GND.n2271 0.11
R3574 GND.n2286 GND.n2284 0.11
R3575 GND.n2298 GND.n2296 0.11
R3576 GND.n2311 GND.n2309 0.11
R3577 GND.n486 GND.n458 0.11
R3578 GND.n488 GND.n453 0.11
R3579 GND.n500 GND.n499 0.11
R3580 GND.n512 GND.n510 0.11
R3581 GND.n521 GND.n437 0.11
R3582 GND.n523 GND.n432 0.11
R3583 GND.n537 GND.n534 0.11
R3584 GND.n551 GND.n417 0.11
R3585 GND.n563 GND.n562 0.11
R3586 GND.n615 GND.n573 0.11
R3587 GND.n613 GND.n574 0.11
R3588 GND.n604 GND.n603 0.11
R3589 GND.n597 GND.n596 0.11
R3590 GND.n590 GND.n589 0.11
R3591 GND.n2061 GND.n1900 0.11
R3592 GND.n2052 GND.n2051 0.11
R3593 GND.n2042 GND.n1910 0.11
R3594 GND.n2040 GND.n1911 0.11
R3595 GND.n2026 GND.n1916 0.11
R3596 GND.n2024 GND.n1917 0.11
R3597 GND.n2010 GND.n1922 0.11
R3598 GND.n1999 GND.n1926 0.11
R3599 GND.n1990 GND.n1989 0.11
R3600 GND.n1983 GND.n1982 0.11
R3601 GND.n1976 GND.n1975 0.11
R3602 GND.n1969 GND.n1968 0.11
R3603 GND.n1962 GND.n1961 0.11
R3604 GND.n1955 GND.n1954 0.11
R3605 GND.n831 GND.n803 0.11
R3606 GND.n833 GND.n798 0.11
R3607 GND.n845 GND.n844 0.11
R3608 GND.n857 GND.n855 0.11
R3609 GND.n866 GND.n782 0.11
R3610 GND.n868 GND.n777 0.11
R3611 GND.n882 GND.n879 0.11
R3612 GND.n896 GND.n762 0.11
R3613 GND.n908 GND.n907 0.11
R3614 GND.n960 GND.n918 0.11
R3615 GND.n958 GND.n919 0.11
R3616 GND.n949 GND.n948 0.11
R3617 GND.n942 GND.n941 0.11
R3618 GND.n935 GND.n934 0.11
R3619 GND.n1812 GND.n1651 0.11
R3620 GND.n1803 GND.n1802 0.11
R3621 GND.n1793 GND.n1661 0.11
R3622 GND.n1791 GND.n1662 0.11
R3623 GND.n1777 GND.n1667 0.11
R3624 GND.n1775 GND.n1668 0.11
R3625 GND.n1761 GND.n1673 0.11
R3626 GND.n1750 GND.n1677 0.11
R3627 GND.n1741 GND.n1740 0.11
R3628 GND.n1734 GND.n1733 0.11
R3629 GND.n1727 GND.n1726 0.11
R3630 GND.n1720 GND.n1719 0.11
R3631 GND.n1713 GND.n1712 0.11
R3632 GND.n1706 GND.n1705 0.11
R3633 GND.n1169 GND.n1168 0.11
R3634 GND.n1181 GND.n1179 0.11
R3635 GND.n1190 GND.n1134 0.11
R3636 GND.n1192 GND.n1129 0.11
R3637 GND.n1204 GND.n1203 0.11
R3638 GND.n1218 GND.n1214 0.11
R3639 GND.n1216 GND.n1114 0.11
R3640 GND.n1243 GND.n1241 0.11
R3641 GND.n1254 GND.n1100 0.11
R3642 GND.n1258 GND.n1257 0.11
R3643 GND.n1296 GND.n1267 0.11
R3644 GND.n1294 GND.n1268 0.11
R3645 GND.n1286 GND.n1285 0.11
R3646 GND.n1280 GND.n1279 0.11
R3647 GND.n1558 GND.n1417 0.11
R3648 GND.n1556 GND.n1418 0.11
R3649 GND.n1548 GND.n1547 0.11
R3650 GND.n1543 GND.n1542 0.11
R3651 GND.n1538 GND.n1537 0.11
R3652 GND.n1533 GND.n1532 0.11
R3653 GND.n1528 GND.n1527 0.11
R3654 GND.n1516 GND.n1515 0.11
R3655 GND.n1510 GND.n1509 0.11
R3656 GND.n1504 GND.n1503 0.11
R3657 GND.n1498 GND.n1497 0.11
R3658 GND.n1492 GND.n1491 0.11
R3659 GND.n1486 GND.n1485 0.11
R3660 GND.n1480 GND.n1479 0.11
R3661 GND.n1481 GND.n1378 0.088
R3662 GND.n1281 GND.n1085 0.087
R3663 GND GND.n2366 0.084
R3664 GND.n2097 GND.n344 0.061
R3665 GND.n1848 GND.n689 0.061
R3666 GND.n1599 GND.n1034 0.061
R3667 GND.n2345 GND.n261 0.051
R3668 GND.n2096 GND.n626 0.051
R3669 GND.n1847 GND.n971 0.051
R3670 GND.n1598 GND.n1315 0.051
R3671 GND.n1597 GND.n1576 0.05
R3672 GND.n1846 GND.n1825 0.05
R3673 GND.n2095 GND.n2074 0.05
R3674 GND.n2344 GND.n2323 0.05
R3675 GND.n1825 GND.n1824 0.049
R3676 GND.n2074 GND.n2073 0.049
R3677 GND.n2323 GND.n2322 0.049
R3678 GND.n2323 GND.n322 0.048
R3679 GND.n2074 GND.n667 0.048
R3680 GND.n1825 GND.n1012 0.048
R3681 GND.n1576 GND.n1356 0.048
R3682 GND GND.n1598 0.048
R3683 GND GND.n1847 0.048
R3684 GND GND.n2345 0.048
R3685 GND GND.n2096 0.047
R3686 GND.n1598 GND.n1597 0.044
R3687 GND.n1847 GND.n1846 0.044
R3688 GND.n2096 GND.n2095 0.044
R3689 GND.n2345 GND.n2344 0.044
R3690 GND.n275 GND.n268 0.04
R3691 GND.n295 GND.n288 0.04
R3692 GND.n315 GND.n308 0.04
R3693 GND.n337 GND.n330 0.04
R3694 GND.n358 GND.n349 0.04
R3695 GND.n640 GND.n631 0.04
R3696 GND.n660 GND.n651 0.04
R3697 GND.n682 GND.n673 0.04
R3698 GND.n703 GND.n694 0.04
R3699 GND.n985 GND.n976 0.04
R3700 GND.n1005 GND.n996 0.04
R3701 GND.n1027 GND.n1018 0.04
R3702 GND.n1048 GND.n1039 0.04
R3703 GND.n1329 GND.n1320 0.04
R3704 GND.n1349 GND.n1340 0.04
R3705 GND.n2359 GND.n2352 0.04
R3706 GND.n1590 GND.n1581 0.04
R3707 GND.n1839 GND.n1830 0.04
R3708 GND.n2088 GND.n2079 0.04
R3709 GND.n2337 GND.n2330 0.04
R3710 GND.n13 GND.n6 0.037
R3711 GND.n723 GND.n714 0.037
R3712 GND.n1068 GND.n1059 0.037
R3713 GND.n1824 GND.n1599 0.037
R3714 GND.n2073 GND.n1848 0.037
R3715 GND.n378 GND.n369 0.036
R3716 GND.n281 GND.n279 0.035
R3717 GND.n301 GND.n299 0.035
R3718 GND.n321 GND.n319 0.035
R3719 GND.n343 GND.n341 0.035
R3720 GND.n364 GND.n345 0.035
R3721 GND.n646 GND.n627 0.035
R3722 GND.n666 GND.n647 0.035
R3723 GND.n688 GND.n669 0.035
R3724 GND.n709 GND.n690 0.035
R3725 GND.n991 GND.n972 0.035
R3726 GND.n1011 GND.n992 0.035
R3727 GND.n1033 GND.n1014 0.035
R3728 GND.n1054 GND.n1035 0.035
R3729 GND.n1335 GND.n1316 0.035
R3730 GND.n1355 GND.n1336 0.035
R3731 GND.n2365 GND.n2363 0.035
R3732 GND.n1596 GND.n1577 0.035
R3733 GND.n1845 GND.n1826 0.035
R3734 GND.n2094 GND.n2075 0.035
R3735 GND.n2343 GND.n2341 0.035
R3736 GND.n52 GND.n50 0.033
R3737 GND.n252 GND.n250 0.033
R3738 GND.n2127 GND.n2125 0.033
R3739 GND.n2313 GND.n2311 0.033
R3740 GND.n476 GND.n458 0.033
R3741 GND.n589 GND.n386 0.033
R3742 GND.n2062 GND.n2061 0.033
R3743 GND.n1954 GND.n1850 0.033
R3744 GND.n821 GND.n803 0.033
R3745 GND.n934 GND.n731 0.033
R3746 GND.n1813 GND.n1812 0.033
R3747 GND.n1705 GND.n1601 0.033
R3748 GND.n1168 GND.n1148 0.033
R3749 GND.n1279 GND.n1076 0.033
R3750 GND.n1417 GND.n1395 0.033
R3751 GND.n1479 GND.n1359 0.033
R3752 GND.n19 GND.n17 0.032
R3753 GND.n729 GND.n710 0.032
R3754 GND.n1074 GND.n1055 0.032
R3755 GND.n2322 GND.n2097 0.032
R3756 GND.n150 GND.n148 0.031
R3757 GND.n172 GND.n160 0.031
R3758 GND.n2214 GND.n2212 0.031
R3759 GND.n2234 GND.n2224 0.031
R3760 GND.n537 GND.n536 0.031
R3761 GND.n551 GND.n550 0.031
R3762 GND.n384 GND.n365 0.031
R3763 GND.n2010 GND.n2009 0.031
R3764 GND.n2000 GND.n1999 0.031
R3765 GND.n882 GND.n881 0.031
R3766 GND.n896 GND.n895 0.031
R3767 GND.n1761 GND.n1760 0.031
R3768 GND.n1751 GND.n1750 0.031
R3769 GND.n1228 GND.n1114 0.031
R3770 GND.n1241 GND.n1107 0.031
R3771 GND.n1527 GND.n1442 0.031
R3772 GND.n1516 GND.n1452 0.031
R3773 GND.n2318 GND.n2317 0.03
R3774 GND.n1572 GND.n1571 0.03
R3775 GND.n2069 GND.n2068 0.029
R3776 GND.n1820 GND.n1819 0.029
R3777 GND.n1311 GND.n1310 0.029
R3778 GND.n257 GND.n256 0.029
R3779 GND.n622 GND.n621 0.029
R3780 GND.n967 GND.n966 0.029
R3781 GND.n66 GND.n64 0.029
R3782 GND.n239 GND.n237 0.029
R3783 GND.n2140 GND.n2138 0.029
R3784 GND.n2300 GND.n2298 0.029
R3785 GND.n488 GND.n487 0.029
R3786 GND.n596 GND.n582 0.029
R3787 GND.n2053 GND.n2052 0.029
R3788 GND.n1961 GND.n1947 0.029
R3789 GND.n833 GND.n832 0.029
R3790 GND.n941 GND.n927 0.029
R3791 GND.n1804 GND.n1803 0.029
R3792 GND.n1712 GND.n1698 0.029
R3793 GND.n1179 GND.n1142 0.029
R3794 GND.n1285 GND.n1271 0.029
R3795 GND.n1557 GND.n1556 0.029
R3796 GND.n1485 GND.n1473 0.029
R3797 GND.n134 GND.n132 0.027
R3798 GND.n186 GND.n176 0.027
R3799 GND.n2200 GND.n2198 0.027
R3800 GND.n2246 GND.n2238 0.027
R3801 GND.n432 GND.n430 0.027
R3802 GND.n562 GND.n561 0.027
R3803 GND.n1921 GND.n1917 0.027
R3804 GND.n1990 GND.n1930 0.027
R3805 GND.n777 GND.n775 0.027
R3806 GND.n907 GND.n906 0.027
R3807 GND.n1672 GND.n1668 0.027
R3808 GND.n1741 GND.n1681 0.027
R3809 GND.n1218 GND.n1217 0.027
R3810 GND.n1242 GND.n1100 0.027
R3811 GND.n1532 GND.n1437 0.027
R3812 GND.n1510 GND.n1453 0.027
R3813 GND.n80 GND.n78 0.025
R3814 GND.n227 GND.n225 0.025
R3815 GND.n2152 GND.n2150 0.025
R3816 GND.n2288 GND.n2286 0.025
R3817 GND.n499 GND.n451 0.025
R3818 GND.n603 GND.n576 0.025
R3819 GND.n1910 GND.n1902 0.025
R3820 GND.n1968 GND.n1944 0.025
R3821 GND.n844 GND.n796 0.025
R3822 GND.n948 GND.n921 0.025
R3823 GND.n1661 GND.n1653 0.025
R3824 GND.n1719 GND.n1695 0.025
R3825 GND.n1180 GND.n1134 0.025
R3826 GND.n1287 GND.n1268 0.025
R3827 GND.n1549 GND.n1548 0.025
R3828 GND.n1491 GND.n1469 0.025
R3829 GND.n1599 GND 0.023
R3830 GND.n1848 GND 0.023
R3831 GND.n2097 GND 0.023
R3832 GND.n120 GND.n118 0.022
R3833 GND.n198 GND.n190 0.022
R3834 GND.n2188 GND.n2186 0.022
R3835 GND.n2259 GND.n2250 0.022
R3836 GND.n522 GND.n521 0.022
R3837 GND.n573 GND.n411 0.022
R3838 GND.n2026 GND.n2025 0.022
R3839 GND.n1983 GND.n1931 0.022
R3840 GND.n867 GND.n866 0.022
R3841 GND.n918 GND.n756 0.022
R3842 GND.n1777 GND.n1776 0.022
R3843 GND.n1734 GND.n1682 0.022
R3844 GND.n1204 GND.n1121 0.022
R3845 GND.n1258 GND.n1255 0.022
R3846 GND.n1537 GND.n1432 0.022
R3847 GND.n1504 GND.n1457 0.022
R3848 GND.n94 GND.n92 0.02
R3849 GND.n214 GND.n212 0.02
R3850 GND.n2165 GND.n2163 0.02
R3851 GND.n2275 GND.n2273 0.02
R3852 GND.n510 GND.n445 0.02
R3853 GND.n605 GND.n574 0.02
R3854 GND.n2041 GND.n2040 0.02
R3855 GND.n1975 GND.n1939 0.02
R3856 GND.n855 GND.n790 0.02
R3857 GND.n950 GND.n919 0.02
R3858 GND.n1792 GND.n1791 0.02
R3859 GND.n1726 GND.n1690 0.02
R3860 GND.n1192 GND.n1191 0.02
R3861 GND.n1296 GND.n1295 0.02
R3862 GND.n1543 GND.n1420 0.02
R3863 GND.n1497 GND.n1465 0.02
R3864 GND.n106 GND.n104 0.018
R3865 GND.n210 GND.n202 0.018
R3866 GND.n2175 GND.n2173 0.018
R3867 GND.n2271 GND.n2263 0.018
R3868 GND.n512 GND.n511 0.018
R3869 GND.n614 GND.n613 0.018
R3870 GND.n1915 GND.n1911 0.018
R3871 GND.n1976 GND.n1936 0.018
R3872 GND.n857 GND.n856 0.018
R3873 GND.n959 GND.n958 0.018
R3874 GND.n1666 GND.n1662 0.018
R3875 GND.n1727 GND.n1687 0.018
R3876 GND.n1129 GND.n1127 0.018
R3877 GND.n1267 GND.n1092 0.018
R3878 GND.n1542 GND.n1427 0.018
R3879 GND.n1498 GND.n1461 0.018
R3880 GND.n108 GND.n106 0.016
R3881 GND.n202 GND.n200 0.016
R3882 GND.n2177 GND.n2175 0.016
R3883 GND.n2263 GND.n2261 0.016
R3884 GND.n511 GND.n437 0.016
R3885 GND.n615 GND.n614 0.016
R3886 GND.n1916 GND.n1915 0.016
R3887 GND.n1982 GND.n1936 0.016
R3888 GND.n856 GND.n782 0.016
R3889 GND.n960 GND.n959 0.016
R3890 GND.n1667 GND.n1666 0.016
R3891 GND.n1733 GND.n1687 0.016
R3892 GND.n1203 GND.n1127 0.016
R3893 GND.n1257 GND.n1092 0.016
R3894 GND.n1538 GND.n1427 0.016
R3895 GND.n1503 GND.n1461 0.016
R3896 GND.n92 GND.n90 0.014
R3897 GND.n223 GND.n214 0.014
R3898 GND.n2163 GND.n2161 0.014
R3899 GND.n2284 GND.n2275 0.014
R3900 GND.n500 GND.n445 0.014
R3901 GND.n605 GND.n604 0.014
R3902 GND.n2042 GND.n2041 0.014
R3903 GND.n1969 GND.n1939 0.014
R3904 GND.n845 GND.n790 0.014
R3905 GND.n950 GND.n949 0.014
R3906 GND.n1793 GND.n1792 0.014
R3907 GND.n1720 GND.n1690 0.014
R3908 GND.n1191 GND.n1190 0.014
R3909 GND.n1295 GND.n1294 0.014
R3910 GND.n1547 GND.n1420 0.014
R3911 GND.n1492 GND.n1465 0.014
R3912 GND.n122 GND.n120 0.012
R3913 GND.n190 GND.n188 0.012
R3914 GND.n2190 GND.n2188 0.012
R3915 GND.n2250 GND.n2248 0.012
R3916 GND.n523 GND.n522 0.012
R3917 GND.n563 GND.n411 0.012
R3918 GND.n2025 GND.n2024 0.012
R3919 GND.n1989 GND.n1931 0.012
R3920 GND.n868 GND.n867 0.012
R3921 GND.n908 GND.n756 0.012
R3922 GND.n1776 GND.n1775 0.012
R3923 GND.n1740 GND.n1682 0.012
R3924 GND.n1214 GND.n1121 0.012
R3925 GND.n1255 GND.n1254 0.012
R3926 GND.n1533 GND.n1432 0.012
R3927 GND.n1509 GND.n1457 0.012
R3928 GND.n78 GND.n76 0.01
R3929 GND.n235 GND.n227 0.01
R3930 GND.n17 GND.n15 0.01
R3931 GND.n279 GND.n277 0.01
R3932 GND.n299 GND.n297 0.01
R3933 GND.n319 GND.n317 0.01
R3934 GND.n2150 GND.n2148 0.01
R3935 GND.n2296 GND.n2288 0.01
R3936 GND.n341 GND.n339 0.01
R3937 GND.n453 GND.n451 0.01
R3938 GND.n597 GND.n576 0.01
R3939 GND.n359 GND.n345 0.01
R3940 GND.n641 GND.n627 0.01
R3941 GND.n661 GND.n647 0.01
R3942 GND.n2051 GND.n1902 0.01
R3943 GND.n1962 GND.n1944 0.01
R3944 GND.n683 GND.n669 0.01
R3945 GND.n798 GND.n796 0.01
R3946 GND.n942 GND.n921 0.01
R3947 GND.n724 GND.n710 0.01
R3948 GND.n704 GND.n690 0.01
R3949 GND.n986 GND.n972 0.01
R3950 GND.n1006 GND.n992 0.01
R3951 GND.n1802 GND.n1653 0.01
R3952 GND.n1713 GND.n1695 0.01
R3953 GND.n1028 GND.n1014 0.01
R3954 GND.n1181 GND.n1180 0.01
R3955 GND.n1287 GND.n1286 0.01
R3956 GND.n1069 GND.n1055 0.01
R3957 GND.n1049 GND.n1035 0.01
R3958 GND.n1330 GND.n1316 0.01
R3959 GND.n1350 GND.n1336 0.01
R3960 GND.n1549 GND.n1418 0.01
R3961 GND.n1486 GND.n1469 0.01
R3962 GND.n2363 GND.n2361 0.01
R3963 GND.n1591 GND.n1577 0.01
R3964 GND.n1840 GND.n1826 0.01
R3965 GND.n2089 GND.n2075 0.01
R3966 GND.n2341 GND.n2339 0.01
R3967 GND.n379 GND.n365 0.009
R3968 GND.n136 GND.n134 0.008
R3969 GND.n176 GND.n174 0.008
R3970 GND.n2202 GND.n2200 0.008
R3971 GND.n2238 GND.n2236 0.008
R3972 GND.n534 GND.n430 0.008
R3973 GND.n561 GND.n417 0.008
R3974 GND.n1922 GND.n1921 0.008
R3975 GND.n1930 GND.n1926 0.008
R3976 GND.n879 GND.n775 0.008
R3977 GND.n906 GND.n762 0.008
R3978 GND.n1673 GND.n1672 0.008
R3979 GND.n1681 GND.n1677 0.008
R3980 GND.n1217 GND.n1216 0.008
R3981 GND.n1243 GND.n1242 0.008
R3982 GND.n1528 GND.n1437 0.008
R3983 GND.n1515 GND.n1453 0.008
R3984 GND.n2323 GND.n323 0.007
R3985 GND.n2074 GND.n668 0.007
R3986 GND.n1825 GND.n1013 0.007
R3987 GND.n1576 GND.n1357 0.007
R3988 GND.n64 GND.n62 0.006
R3989 GND.n248 GND.n239 0.006
R3990 GND.n2138 GND.n2136 0.006
R3991 GND.n2309 GND.n2300 0.006
R3992 GND.n487 GND.n486 0.006
R3993 GND.n590 GND.n582 0.006
R3994 GND.n2053 GND.n1900 0.006
R3995 GND.n1955 GND.n1947 0.006
R3996 GND.n832 GND.n831 0.006
R3997 GND.n935 GND.n927 0.006
R3998 GND.n1804 GND.n1651 0.006
R3999 GND.n1706 GND.n1698 0.006
R4000 GND.n1169 GND.n1142 0.006
R4001 GND.n1280 GND.n1271 0.006
R4002 GND.n1558 GND.n1557 0.006
R4003 GND.n1480 GND.n1473 0.006
R4004 GND.n6 GND.n4 0.005
R4005 GND.n268 GND.n266 0.005
R4006 GND.n288 GND.n286 0.005
R4007 GND.n308 GND.n306 0.005
R4008 GND.n330 GND.n328 0.005
R4009 GND.n352 GND.n349 0.005
R4010 GND.n634 GND.n631 0.005
R4011 GND.n654 GND.n651 0.005
R4012 GND.n676 GND.n673 0.005
R4013 GND.n717 GND.n714 0.005
R4014 GND.n697 GND.n694 0.005
R4015 GND.n979 GND.n976 0.005
R4016 GND.n999 GND.n996 0.005
R4017 GND.n1021 GND.n1018 0.005
R4018 GND.n1062 GND.n1059 0.005
R4019 GND.n1042 GND.n1039 0.005
R4020 GND.n1323 GND.n1320 0.005
R4021 GND.n1343 GND.n1340 0.005
R4022 GND.n2352 GND.n2350 0.005
R4023 GND.n1584 GND.n1581 0.005
R4024 GND.n1833 GND.n1830 0.005
R4025 GND.n2082 GND.n2079 0.005
R4026 GND.n2330 GND.n2328 0.005
R4027 GND.n152 GND.n150 0.004
R4028 GND.n160 GND.n158 0.004
R4029 GND.n2216 GND.n2214 0.004
R4030 GND.n2224 GND.n2222 0.004
R4031 GND.n536 GND.n535 0.004
R4032 GND.n550 GND.n549 0.004
R4033 GND.n372 GND.n369 0.004
R4034 GND.n2009 GND.n2008 0.004
R4035 GND.n2001 GND.n2000 0.004
R4036 GND.n881 GND.n880 0.004
R4037 GND.n895 GND.n894 0.004
R4038 GND.n1760 GND.n1759 0.004
R4039 GND.n1752 GND.n1751 0.004
R4040 GND.n1229 GND.n1228 0.004
R4041 GND.n1231 GND.n1107 0.004
R4042 GND.n1523 GND.n1442 0.004
R4043 GND.n1452 GND.n1447 0.004
R4044 GND.n50 GND.n48 0.002
R4045 GND.n259 GND.n252 0.002
R4046 GND.n2125 GND.n2123 0.002
R4047 GND.n2320 GND.n2313 0.002
R4048 GND.n477 GND.n476 0.002
R4049 GND.n624 GND.n386 0.002
R4050 GND.n2063 GND.n2062 0.002
R4051 GND.n2071 GND.n1850 0.002
R4052 GND.n822 GND.n821 0.002
R4053 GND.n969 GND.n731 0.002
R4054 GND.n1814 GND.n1813 0.002
R4055 GND.n1822 GND.n1601 0.002
R4056 GND.n1150 GND.n1148 0.002
R4057 GND.n1313 GND.n1076 0.002
R4058 GND.n1401 GND.n1395 0.002
R4059 GND.n1574 GND.n1359 0.002
R4060 fout5.n510 fout5.t3 1038.92
R4061 fout5.n388 fout5.t13 1037.29
R4062 fout5.n389 fout5.t7 797.185
R4063 fout5.n525 fout5.t4 795.549
R4064 fout5.n367 fout5.t5 732.331
R4065 fout5.n479 fout5.t8 731.671
R4066 fout5.n417 fout5.t11 731.671
R4067 fout5.n497 fout5.t14 730.667
R4068 fout5.n496 fout5.t6 400.619
R4069 fout5.n453 fout5.t12 400.601
R4070 fout5.n11 fout5.t9 397.315
R4071 fout5.n497 fout5.t10 395.829
R4072 fout5.n244 fout5.n243 13.176
R4073 fout5.n14 fout5.t2 11.721
R4074 fout5.n14 fout5.t1 10.994
R4075 fout5.n23 fout5.n22 9.3
R4076 fout5.n322 fout5.n321 9.3
R4077 fout5.n288 fout5.n287 9.3
R4078 fout5.n285 fout5.n284 9.3
R4079 fout5.n222 fout5.n221 9.3
R4080 fout5.n336 fout5.n335 9.3
R4081 fout5.n338 fout5.n337 9.3
R4082 fout5.n220 fout5.n219 9.3
R4083 fout5.n253 fout5.n252 9.3
R4084 fout5.n266 fout5.n265 9.3
R4085 fout5.n274 fout5.n273 9.3
R4086 fout5.n277 fout5.n276 9.3
R4087 fout5.n137 fout5.n136 9.3
R4088 fout5.n134 fout5.n133 9.3
R4089 fout5.n50 fout5.n49 9.3
R4090 fout5.n48 fout5.n47 9.3
R4091 fout5.n41 fout5.n40 8.097
R4092 fout5.n276 fout5.n275 5.457
R4093 fout5.n136 fout5.n135 5.08
R4094 fout5.n39 fout5.n38 4.65
R4095 fout5.n146 fout5.n145 4.65
R4096 fout5.n55 fout5.n53 4.5
R4097 fout5.n107 fout5.n103 4.5
R4098 fout5.n111 fout5.n100 4.5
R4099 fout5.n126 fout5.n125 4.5
R4100 fout5.n81 fout5.n80 4.5
R4101 fout5.n255 fout5.n247 4.5
R4102 fout5.n262 fout5.n245 4.5
R4103 fout5.n271 fout5.n242 4.5
R4104 fout5.n294 fout5.n293 4.5
R4105 fout5.n342 fout5.n341 4.5
R4106 fout5.n330 fout5.n329 4.5
R4107 fout5.n230 fout5.n229 4.5
R4108 fout5.n237 fout5.n236 4.5
R4109 fout5.n302 fout5.n301 4.5
R4110 fout5.n282 fout5.n281 4.5
R4111 fout5.n119 fout5.n118 4.5
R4112 fout5.n213 fout5.n212 4.5
R4113 fout5.n27 fout5.n25 4.5
R4114 fout5.n229 fout5.n227 4.314
R4115 fout5.n301 fout5.n298 3.944
R4116 fout5.n103 fout5.n102 3.937
R4117 fout5.n118 fout5.n117 3.567
R4118 fout5.n147 fout5.n140 3.033
R4119 fout5.n43 fout5.n42 3.033
R4120 fout5.n40 fout5.t0 2.9
R4121 fout5.n300 fout5.n299 2.258
R4122 fout5.n116 fout5.n115 2.258
R4123 fout5.n235 fout5.n234 1.882
R4124 fout5.n236 fout5.n235 1.882
R4125 fout5.n99 fout5.n98 1.882
R4126 fout5.n350 fout5.n14 1.518
R4127 fout5.n118 fout5.n116 1.505
R4128 fout5.n100 fout5.n99 1.505
R4129 fout5.n56 fout5.n55 1.5
R4130 fout5.n343 fout5.n342 1.5
R4131 fout5.n82 fout5.n81 1.5
R4132 fout5.n148 fout5.n147 1.5
R4133 fout5.n127 fout5.n126 1.5
R4134 fout5.n214 fout5.n213 1.5
R4135 fout5.n28 fout5.n27 1.5
R4136 fout5.n465 fout5.n464 1.435
R4137 fout5.n448 fout5.n447 1.435
R4138 fout5.n402 fout5.n388 1.388
R4139 fout5.n390 fout5.n389 1.355
R4140 fout5.n527 fout5.n525 1.355
R4141 fout5.n511 fout5.n510 1.355
R4142 fout5.n369 fout5.n367 1.354
R4143 fout5.n419 fout5.n417 1.354
R4144 fout5.n12 fout5.n11 1.354
R4145 fout5.n481 fout5.n479 1.354
R4146 fout5.n13 fout5.n12 1.142
R4147 fout5.n482 fout5.n481 1.142
R4148 fout5.n528 fout5.n527 1.142
R4149 fout5.n420 fout5.n419 1.14
R4150 fout5.n362 fout5.n13 1.138
R4151 fout5.n483 fout5.n482 1.138
R4152 fout5.n529 fout5.n528 1.138
R4153 fout5.n359 fout5.n358 1.137
R4154 fout5.n375 fout5.n374 1.137
R4155 fout5.n354 fout5.n353 1.137
R4156 fout5.n3 fout5.n2 1.137
R4157 fout5.n370 fout5.n369 1.137
R4158 fout5.n512 fout5.n511 1.137
R4159 fout5.n538 fout5.n537 1.137
R4160 fout5.n503 fout5.n502 1.137
R4161 fout5.n533 fout5.n532 1.137
R4162 fout5.n518 fout5.n517 1.137
R4163 fout5.n466 fout5.n465 1.137
R4164 fout5.n492 fout5.n491 1.137
R4165 fout5.n458 fout5.n457 1.137
R4166 fout5.n488 fout5.n487 1.137
R4167 fout5.n472 fout5.n471 1.137
R4168 fout5.n449 fout5.n448 1.137
R4169 fout5.n440 fout5.n439 1.137
R4170 fout5.n425 fout5.n424 1.137
R4171 fout5.n430 fout5.n429 1.137
R4172 fout5.n434 fout5.n433 1.137
R4173 fout5.n540 fout5.n539 1.136
R4174 fout5.n494 fout5.n493 1.136
R4175 fout5.n378 fout5.n377 1.136
R4176 fout5.n361 fout5.n360 1.136
R4177 fout5.n468 fout5.n467 1.136
R4178 fout5.n514 fout5.n513 1.136
R4179 fout5.n451 fout5.n450 1.136
R4180 fout5.n341 fout5.n340 1.129
R4181 fout5.n301 fout5.n300 1.129
R4182 fout5.n293 fout5.n292 1.129
R4183 fout5.n303 fout5.n302 1.042
R4184 fout5.n58 fout5.n57 0.853
R4185 fout5.n192 fout5.n191 0.853
R4186 fout5.n150 fout5.n149 0.853
R4187 fout5.n345 fout5.n344 0.853
R4188 fout5.n410 fout5.n409 0.823
R4189 fout5.n212 fout5.n211 0.752
R4190 fout5.n80 fout5.n79 0.752
R4191 fout5.n125 fout5.n124 0.752
R4192 fout5.n103 fout5.n101 0.752
R4193 fout5.n53 fout5.n52 0.752
R4194 fout5.n25 fout5.n24 0.752
R4195 fout5.n30 fout5.n29 0.716
R4196 fout5.n350 fout5.n349 0.69
R4197 fout5.n351 fout5.n350 0.68
R4198 fout5.n252 fout5.n251 0.536
R4199 fout5.n265 fout5.n264 0.536
R4200 fout5.n145 fout5.n144 0.476
R4201 fout5.n287 fout5.n286 0.475
R4202 fout5.n410 fout5.n379 0.468
R4203 fout5.n403 fout5.n402 0.44
R4204 fout5.n42 fout5.n41 0.382
R4205 fout5.n328 fout5.n327 0.382
R4206 fout5.n329 fout5.n328 0.376
R4207 fout5.n229 fout5.n228 0.376
R4208 fout5.n281 fout5.n280 0.376
R4209 fout5.n242 fout5.n241 0.376
R4210 fout5.n245 fout5.n244 0.376
R4211 fout5.n247 fout5.n246 0.376
R4212 fout5.n52 fout5.n51 0.35
R4213 fout5.n340 fout5.n339 0.349
R4214 fout5 fout5.n410 0.234
R4215 fout5.n499 fout5.n498 0.152
R4216 fout5.n496 fout5.n495 0.123
R4217 fout5.n453 fout5.n452 0.123
R4218 fout5.n454 fout5.n453 0.091
R4219 fout5.n367 fout5.n366 0.083
R4220 fout5.n11 fout5.n10 0.083
R4221 fout5.n479 fout5.n478 0.083
R4222 fout5.n417 fout5.n416 0.083
R4223 fout5.n388 fout5.n387 0.075
R4224 fout5.n525 fout5.n524 0.075
R4225 fout5.n510 fout5.n509 0.075
R4226 fout5.n498 fout5.n496 0.07
R4227 fout5.n444 fout5.n443 0.064
R4228 fout5.n384 fout5.n383 0.058
R4229 fout5.n324 fout5.n323 0.047
R4230 fout5.n278 fout5.n277 0.047
R4231 fout5.n268 fout5.n267 0.047
R4232 fout5.n259 fout5.n258 0.047
R4233 fout5.n249 fout5.n248 0.047
R4234 fout5.n138 fout5.n137 0.047
R4235 fout5.n21 fout5.n20 0.047
R4236 fout5 fout5.n541 0.045
R4237 fout5.n106 fout5.n105 0.043
R4238 fout5.n88 fout5.n87 0.043
R4239 fout5.n226 fout5.n225 0.041
R4240 fout5.n311 fout5.n310 0.041
R4241 fout5.n45 fout5.n44 0.035
R4242 fout5.n181 fout5.n180 0.035
R4243 fout5.n176 fout5.n175 0.035
R4244 fout5.n35 fout5.n34 0.035
R4245 fout5.n333 fout5.n332 0.034
R4246 fout5.n261 fout5.n260 0.034
R4247 fout5.n257 fout5.n256 0.034
R4248 fout5.n48 fout5.n46 0.034
R4249 fout5.n320 fout5.n319 0.034
R4250 fout5.n318 fout5.n317 0.034
R4251 fout5.n170 fout5.n169 0.034
R4252 fout5.n189 fout5.n188 0.034
R4253 fout5.n82 fout5.n75 0.034
R4254 fout5.n84 fout5.n83 0.034
R4255 fout5.n132 fout5.n131 0.034
R4256 fout5.n37 fout5.n36 0.034
R4257 fout5.n336 fout5.n334 0.032
R4258 fout5.n147 fout5.n146 0.032
R4259 fout5.n43 fout5.n39 0.032
R4260 fout5.n187 fout5.n186 0.032
R4261 fout5.n56 fout5.n37 0.032
R4262 fout5.n358 fout5.n356 0.032
R4263 fout5.n397 fout5.n396 0.032
R4264 fout5.n398 fout5.n397 0.032
R4265 fout5.n537 fout5.n535 0.032
R4266 fout5.n487 fout5.n486 0.032
R4267 fout5.n433 fout5.n432 0.032
R4268 fout5.n402 fout5.n401 0.032
R4269 fout5.n71 fout5.n70 0.031
R4270 fout5.n60 fout5.n59 0.031
R4271 fout5.n347 fout5.n346 0.031
R4272 fout5.n205 fout5.n204 0.031
R4273 fout5.n285 fout5.n283 0.03
R4274 fout5.n270 fout5.n269 0.03
R4275 fout5.n77 fout5.n76 0.03
R4276 fout5.n20 fout5.n19 0.03
R4277 fout5.n343 fout5.n320 0.03
R4278 fout5.n315 fout5.n314 0.03
R4279 fout5.n185 fout5.n184 0.03
R4280 fout5.n73 fout5.n72 0.03
R4281 fout5.n85 fout5.n84 0.03
R4282 fout5.n32 fout5.n31 0.03
R4283 fout5.n194 fout5.n193 0.03
R4284 fout5.n163 fout5.n162 0.03
R4285 fout5.n152 fout5.n151 0.03
R4286 fout5.n392 fout5.n391 0.03
R4287 fout5.n325 fout5.n324 0.028
R4288 fout5.n224 fout5.n223 0.028
R4289 fout5.n239 fout5.n238 0.028
R4290 fout5.n302 fout5.n240 0.028
R4291 fout5.n291 fout5.n290 0.028
R4292 fout5.n147 fout5.n139 0.028
R4293 fout5.n113 fout5.n112 0.028
R4294 fout5.n105 fout5.n104 0.028
R4295 fout5.n55 fout5.n50 0.028
R4296 fout5.n27 fout5.n23 0.028
R4297 fout5.n215 fout5.n214 0.028
R4298 fout5.n344 fout5.n218 0.028
R4299 fout5.n313 fout5.n312 0.028
R4300 fout5.n306 fout5.n305 0.028
R4301 fout5.n304 fout5.n303 0.028
R4302 fout5.n168 fout5.n167 0.028
R4303 fout5.n190 fout5.n189 0.028
R4304 fout5.n183 fout5.n182 0.028
R4305 fout5.n174 fout5.n173 0.028
R4306 fout5.n149 fout5.n148 0.028
R4307 fout5.n93 fout5.n92 0.028
R4308 fout5.n87 fout5.n86 0.028
R4309 fout5.n28 fout5.n18 0.028
R4310 fout5.n366 fout5.n365 0.028
R4311 fout5.n364 fout5.n363 0.028
R4312 fout5.n8 fout5.n7 0.028
R4313 fout5.n10 fout5.n9 0.028
R4314 fout5.n374 fout5.n373 0.028
R4315 fout5.n353 fout5.n352 0.028
R4316 fout5.n358 fout5.n357 0.028
R4317 fout5.n2 fout5.n0 0.028
R4318 fout5.n394 fout5.n393 0.028
R4319 fout5.n396 fout5.n395 0.028
R4320 fout5.n399 fout5.n398 0.028
R4321 fout5.n401 fout5.n400 0.028
R4322 fout5.n517 fout5.n516 0.028
R4323 fout5.n532 fout5.n531 0.028
R4324 fout5.n537 fout5.n536 0.028
R4325 fout5.n502 fout5.n500 0.028
R4326 fout5.n478 fout5.n477 0.028
R4327 fout5.n476 fout5.n475 0.028
R4328 fout5.n462 fout5.n461 0.028
R4329 fout5.n464 fout5.n463 0.028
R4330 fout5.n471 fout5.n470 0.028
R4331 fout5.n487 fout5.n485 0.028
R4332 fout5.n491 fout5.n490 0.028
R4333 fout5.n457 fout5.n455 0.028
R4334 fout5.n416 fout5.n415 0.028
R4335 fout5.n445 fout5.n444 0.028
R4336 fout5.n447 fout5.n446 0.028
R4337 fout5.n429 fout5.n428 0.028
R4338 fout5.n439 fout5.n437 0.028
R4339 fout5.n67 fout5.n66 0.027
R4340 fout5.n64 fout5.n63 0.027
R4341 fout5.n342 fout5.n338 0.026
R4342 fout5.n282 fout5.n279 0.026
R4343 fout5.n142 fout5.n141 0.026
R4344 fout5.n119 fout5.n114 0.026
R4345 fout5.n165 fout5.n164 0.026
R4346 fout5.n191 fout5.n171 0.026
R4347 fout5.n130 fout5.n129 0.026
R4348 fout5.n95 fout5.n94 0.026
R4349 fout5.n90 fout5.n89 0.026
R4350 fout5.n17 fout5.n16 0.026
R4351 fout5.n201 fout5.n200 0.026
R4352 fout5.n198 fout5.n197 0.026
R4353 fout5.n159 fout5.n158 0.026
R4354 fout5.n156 fout5.n155 0.026
R4355 fout5.n381 fout5.n380 0.025
R4356 fout5.n383 fout5.n382 0.025
R4357 fout5.n385 fout5.n384 0.025
R4358 fout5.n387 fout5.n386 0.025
R4359 fout5.n524 fout5.n523 0.025
R4360 fout5.n522 fout5.n521 0.025
R4361 fout5.n507 fout5.n506 0.025
R4362 fout5.n509 fout5.n508 0.025
R4363 fout5.n29 fout5.n28 0.024
R4364 fout5.n289 fout5.n288 0.024
R4365 fout5.n146 fout5.n143 0.024
R4366 fout5.n217 fout5.n216 0.024
R4367 fout5.n309 fout5.n308 0.024
R4368 fout5.n171 fout5.n170 0.024
R4369 fout5.n178 fout5.n177 0.024
R4370 fout5.n127 fout5.n97 0.024
R4371 fout5.n406 fout5.n405 0.023
R4372 fout5.n232 fout5.n231 0.022
R4373 fout5.n279 fout5.n278 0.022
R4374 fout5.n266 fout5.n263 0.022
R4375 fout5.n254 fout5.n253 0.022
R4376 fout5.n143 fout5.n142 0.022
R4377 fout5.n109 fout5.n108 0.022
R4378 fout5.n218 fout5.n217 0.022
R4379 fout5.n191 fout5.n190 0.022
R4380 fout5.n179 fout5.n178 0.022
R4381 fout5.n148 fout5.n132 0.022
R4382 fout5.n131 fout5.n130 0.022
R4383 fout5.n296 fout5.n295 0.02
R4384 fout5.n294 fout5.n291 0.02
R4385 fout5.n290 fout5.n289 0.02
R4386 fout5.n139 fout5.n138 0.02
R4387 fout5.n123 fout5.n122 0.02
R4388 fout5.n214 fout5.n208 0.02
R4389 fout5.n344 fout5.n343 0.02
R4390 fout5.n169 fout5.n168 0.02
R4391 fout5.n149 fout5.n85 0.02
R4392 fout5.n16 fout5.n15 0.02
R4393 fout5.n59 fout5.n58 0.019
R4394 fout5.n58 fout5.n30 0.019
R4395 fout5.n346 fout5.n345 0.019
R4396 fout5.n345 fout5.n205 0.019
R4397 fout5.n308 fout5.n307 0.018
R4398 fout5.n57 fout5.n56 0.018
R4399 fout5.n150 fout5.n71 0.018
R4400 fout5.n193 fout5.n192 0.018
R4401 fout5.n192 fout5.n163 0.018
R4402 fout5.n151 fout5.n150 0.018
R4403 fout5.n210 fout5.n209 0.017
R4404 fout5.n223 fout5.n222 0.017
R4405 fout5.n272 fout5.n271 0.017
R4406 fout5.n269 fout5.n268 0.017
R4407 fout5.n208 fout5.n207 0.017
R4408 fout5.n314 fout5.n313 0.017
R4409 fout5.n167 fout5.n166 0.017
R4410 fout5.n188 fout5.n187 0.017
R4411 fout5.n186 fout5.n185 0.017
R4412 fout5.n184 fout5.n183 0.017
R4413 fout5.n129 fout5.n128 0.017
R4414 fout5.n97 fout5.n96 0.017
R4415 fout5.n91 fout5.n90 0.017
R4416 fout5.n369 fout5.n368 0.017
R4417 fout5.n374 fout5.n372 0.017
R4418 fout5.n2 fout5.n1 0.017
R4419 fout5.n12 fout5.n6 0.017
R4420 fout5.n391 fout5.n390 0.017
R4421 fout5.n393 fout5.n392 0.017
R4422 fout5.n527 fout5.n526 0.017
R4423 fout5.n517 fout5.n515 0.017
R4424 fout5.n502 fout5.n501 0.017
R4425 fout5.n511 fout5.n505 0.017
R4426 fout5.n481 fout5.n480 0.017
R4427 fout5.n471 fout5.n469 0.017
R4428 fout5.n457 fout5.n456 0.017
R4429 fout5.n465 fout5.n460 0.017
R4430 fout5.n419 fout5.n418 0.017
R4431 fout5.n424 fout5.n423 0.017
R4432 fout5.n439 fout5.n438 0.017
R4433 fout5.n448 fout5.n442 0.017
R4434 fout5.n359 fout5.n355 0.016
R4435 fout5.n533 fout5.n530 0.016
R4436 fout5.n538 fout5.n534 0.016
R4437 fout5.n488 fout5.n484 0.016
R4438 fout5.n492 fout5.n489 0.016
R4439 fout5.n430 fout5.n426 0.016
R4440 fout5.n435 fout5.n434 0.016
R4441 fout5.n326 fout5.n325 0.015
R4442 fout5.n334 fout5.n333 0.015
R4443 fout5.n240 fout5.n239 0.015
R4444 fout5.n81 fout5.n78 0.015
R4445 fout5.n114 fout5.n113 0.015
R4446 fout5.n112 fout5.n111 0.015
R4447 fout5.n319 fout5.n318 0.015
R4448 fout5.n317 fout5.n316 0.015
R4449 fout5.n305 fout5.n304 0.015
R4450 fout5.n75 fout5.n74 0.015
R4451 fout5.n83 fout5.n82 0.015
R4452 fout5.n94 fout5.n93 0.015
R4453 fout5.n92 fout5.n91 0.015
R4454 fout5.n365 fout5.n364 0.015
R4455 fout5.n9 fout5.n8 0.015
R4456 fout5.n395 fout5.n394 0.015
R4457 fout5.n400 fout5.n399 0.015
R4458 fout5.n477 fout5.n476 0.015
R4459 fout5.n463 fout5.n462 0.015
R4460 fout5.n415 fout5.n414 0.015
R4461 fout5.n446 fout5.n445 0.015
R4462 fout5.n428 fout5.n427 0.015
R4463 fout5.n437 fout5.n436 0.015
R4464 fout5.n332 fout5.n331 0.013
R4465 fout5.n238 fout5.n237 0.013
R4466 fout5.n274 fout5.n272 0.013
R4467 fout5.n44 fout5.n43 0.013
R4468 fout5.n46 fout5.n45 0.013
R4469 fout5.n307 fout5.n306 0.013
R4470 fout5.n34 fout5.n33 0.013
R4471 fout5.n36 fout5.n35 0.013
R4472 fout5.n349 fout5.n348 0.013
R4473 fout5.n382 fout5.n381 0.013
R4474 fout5.n386 fout5.n385 0.013
R4475 fout5.n523 fout5.n522 0.013
R4476 fout5.n508 fout5.n507 0.013
R4477 fout5.n66 fout5.n65 0.012
R4478 fout5.n65 fout5.n64 0.012
R4479 fout5.n360 fout5.n354 0.012
R4480 fout5.n360 fout5.n359 0.012
R4481 fout5.n539 fout5.n533 0.012
R4482 fout5.n539 fout5.n538 0.012
R4483 fout5.n493 fout5.n488 0.012
R4484 fout5.n493 fout5.n492 0.012
R4485 fout5.n431 fout5.n430 0.012
R4486 fout5.n434 fout5.n431 0.012
R4487 fout5.n297 fout5.n296 0.011
R4488 fout5.n122 fout5.n121 0.011
R4489 fout5.n69 fout5.n68 0.011
R4490 fout5.n62 fout5.n61 0.011
R4491 fout5.n200 fout5.n199 0.011
R4492 fout5.n199 fout5.n198 0.011
R4493 fout5.n196 fout5.n195 0.011
R4494 fout5.n161 fout5.n160 0.011
R4495 fout5.n158 fout5.n157 0.011
R4496 fout5.n157 fout5.n156 0.011
R4497 fout5.n154 fout5.n153 0.011
R4498 fout5.n203 fout5.n202 0.011
R4499 fout5.n377 fout5.n376 0.011
R4500 fout5.n5 fout5.n4 0.011
R4501 fout5.n520 fout5.n519 0.011
R4502 fout5.n513 fout5.n504 0.011
R4503 fout5.n474 fout5.n473 0.011
R4504 fout5.n467 fout5.n459 0.011
R4505 fout5.n422 fout5.n421 0.011
R4506 fout5.n450 fout5.n441 0.011
R4507 fout5.n375 fout5.n371 0.01
R4508 fout5.n426 fout5.n425 0.01
R4509 fout5.n440 fout5.n435 0.01
R4510 fout5.n405 fout5.n404 0.01
R4511 fout5.n404 fout5.n403 0.01
R4512 fout5.n323 fout5.n322 0.009
R4513 fout5.n233 fout5.n232 0.009
R4514 fout5.n237 fout5.n233 0.009
R4515 fout5.n260 fout5.n259 0.009
R4516 fout5.n110 fout5.n109 0.009
R4517 fout5.n216 fout5.n215 0.009
R4518 fout5.n180 fout5.n179 0.009
R4519 fout5.n408 fout5.n407 0.009
R4520 fout5.n230 fout5.n226 0.007
R4521 fout5.n263 fout5.n262 0.007
R4522 fout5.n258 fout5.n257 0.007
R4523 fout5.n255 fout5.n254 0.007
R4524 fout5.n111 fout5.n110 0.007
R4525 fout5.n23 fout5.n21 0.007
R4526 fout5.n310 fout5.n309 0.007
R4527 fout5.n182 fout5.n181 0.007
R4528 fout5.n177 fout5.n176 0.007
R4529 fout5.n175 fout5.n174 0.007
R4530 fout5.n18 fout5.n17 0.007
R4531 fout5.n70 fout5.n69 0.006
R4532 fout5.n68 fout5.n67 0.006
R4533 fout5.n63 fout5.n62 0.006
R4534 fout5.n61 fout5.n60 0.006
R4535 fout5.n197 fout5.n196 0.006
R4536 fout5.n195 fout5.n194 0.006
R4537 fout5.n162 fout5.n161 0.006
R4538 fout5.n160 fout5.n159 0.006
R4539 fout5.n155 fout5.n154 0.006
R4540 fout5.n153 fout5.n152 0.006
R4541 fout5.n348 fout5.n347 0.006
R4542 fout5.n204 fout5.n203 0.006
R4543 fout5.n202 fout5.n201 0.006
R4544 fout5.n377 fout5.n370 0.006
R4545 fout5.n376 fout5.n375 0.006
R4546 fout5.n4 fout5.n3 0.006
R4547 fout5.n519 fout5.n518 0.006
R4548 fout5.n504 fout5.n503 0.006
R4549 fout5.n513 fout5.n512 0.006
R4550 fout5.n473 fout5.n472 0.006
R4551 fout5.n459 fout5.n458 0.006
R4552 fout5.n467 fout5.n466 0.006
R4553 fout5.n425 fout5.n422 0.006
R4554 fout5.n441 fout5.n440 0.006
R4555 fout5.n450 fout5.n449 0.006
R4556 fout5.n342 fout5.n326 0.005
R4557 fout5.n338 fout5.n336 0.005
R4558 fout5.n302 fout5.n297 0.005
R4559 fout5.n295 fout5.n294 0.005
R4560 fout5.n267 fout5.n266 0.005
R4561 fout5.n253 fout5.n250 0.005
R4562 fout5.n121 fout5.n120 0.005
R4563 fout5.n107 fout5.n106 0.005
R4564 fout5.n207 fout5.n206 0.005
R4565 fout5.n128 fout5.n127 0.005
R4566 fout5.n89 fout5.n88 0.005
R4567 fout5.n409 fout5.n408 0.005
R4568 fout5.n407 fout5.n406 0.005
R4569 fout5.n541 fout5.n540 0.004
R4570 fout5.n495 fout5.n494 0.004
R4571 fout5.n421 fout5.n420 0.003
R4572 fout5.n361 fout5.n351 0.003
R4573 fout5.n379 fout5.n378 0.003
R4574 fout5.n514 fout5.n499 0.003
R4575 fout5.n468 fout5.n454 0.003
R4576 fout5.n452 fout5.n451 0.003
R4577 fout5.n213 fout5.n210 0.003
R4578 fout5.n81 fout5.n77 0.003
R4579 fout5.n137 fout5.n134 0.003
R4580 fout5.n126 fout5.n123 0.003
R4581 fout5.n108 fout5.n107 0.003
R4582 fout5.n50 fout5.n48 0.003
R4583 fout5.n55 fout5.n54 0.003
R4584 fout5.n27 fout5.n26 0.003
R4585 fout5.n166 fout5.n165 0.003
R4586 fout5.n33 fout5.n32 0.003
R4587 fout5.n13 fout5.n5 0.003
R4588 fout5.n528 fout5.n520 0.003
R4589 fout5.n482 fout5.n474 0.003
R4590 fout5.n412 fout5.n411 0.003
R4591 fout5.n413 fout5.n412 0.002
R4592 fout5.n494 fout5.n483 0.002
R4593 fout5.n540 fout5.n529 0.002
R4594 fout5.n378 fout5.n362 0.002
R4595 fout5.n362 fout5.n361 0.002
R4596 fout5.n451 fout5.n413 0.002
R4597 fout5.n483 fout5.n468 0.002
R4598 fout5.n529 fout5.n514 0.002
R4599 fout5.n331 fout5.n330 0.001
R4600 fout5.n222 fout5.n220 0.001
R4601 fout5.n225 fout5.n224 0.001
R4602 fout5.n231 fout5.n230 0.001
R4603 fout5.n288 fout5.n285 0.001
R4604 fout5.n283 fout5.n282 0.001
R4605 fout5.n277 fout5.n274 0.001
R4606 fout5.n271 fout5.n270 0.001
R4607 fout5.n262 fout5.n261 0.001
R4608 fout5.n256 fout5.n255 0.001
R4609 fout5.n250 fout5.n249 0.001
R4610 fout5.n120 fout5.n119 0.001
R4611 fout5.n316 fout5.n315 0.001
R4612 fout5.n312 fout5.n311 0.001
R4613 fout5.n173 fout5.n172 0.001
R4614 fout5.n74 fout5.n73 0.001
R4615 fout5.n96 fout5.n95 0.001
R4616 fout5.n498 fout5.n497 0.001
R4617 a_n14423_5865.n97 a_n14423_5865.t4 1040.28
R4618 a_n14423_5865.n97 a_n14423_5865.t5 796.134
R4619 a_n14423_5865.n41 a_n14423_5865.n40 13.176
R4620 a_n14423_5865.n95 a_n14423_5865.t0 11.611
R4621 a_n14423_5865.n95 a_n14423_5865.t2 11.295
R4622 a_n14423_5865.n96 a_n14423_5865.t1 10.06
R4623 a_n14423_5865.n151 a_n14423_5865.n34 9.3
R4624 a_n14423_5865.n151 a_n14423_5865.n142 9.3
R4625 a_n14423_5865.n151 a_n14423_5865.n136 9.3
R4626 a_n14423_5865.n151 a_n14423_5865.n49 9.3
R4627 a_n14423_5865.n151 a_n14423_5865.n54 9.3
R4628 a_n14423_5865.n151 a_n14423_5865.n124 9.3
R4629 a_n14423_5865.n151 a_n14423_5865.n150 8.469
R4630 a_n14423_5865.n151 a_n14423_5865.n114 8.469
R4631 a_n14423_5865.n151 a_n14423_5865.n119 8.125
R4632 a_n14423_5865.n151 a_n14423_5865.n29 8.124
R4633 a_n14423_5865.n151 a_n14423_5865.n111 8.097
R4634 a_n14423_5865.n151 a_n14423_5865.n147 8.096
R4635 a_n14423_5865.n151 a_n14423_5865.n127 8.016
R4636 a_n14423_5865.n151 a_n14423_5865.n39 8.016
R4637 a_n14423_5865.n151 a_n14423_5865.n131 7.964
R4638 a_n14423_5865.n151 a_n14423_5865.n44 7.964
R4639 a_n14423_5865.n126 a_n14423_5865.n125 6.4
R4640 a_n14423_5865.n110 a_n14423_5865.n55 6.4
R4641 a_n14423_5865.n145 a_n14423_5865.n144 6.023
R4642 a_n14423_5865.n37 a_n14423_5865.n36 6.023
R4643 a_n14423_5865.n136 a_n14423_5865.n135 6.023
R4644 a_n14423_5865.n43 a_n14423_5865.n42 6.023
R4645 a_n14423_5865.n130 a_n14423_5865.n129 6.023
R4646 a_n14423_5865.n149 a_n14423_5865.n148 5.647
R4647 a_n14423_5865.n49 a_n14423_5865.n46 5.647
R4648 a_n14423_5865.n117 a_n14423_5865.n116 5.647
R4649 a_n14423_5865.n113 a_n14423_5865.n112 5.647
R4650 a_n14423_5865.n133 a_n14423_5865.n132 5.457
R4651 a_n14423_5865.n27 a_n14423_5865.n26 5.27
R4652 a_n14423_5865.n48 a_n14423_5865.n47 5.08
R4653 a_n14423_5865.n34 a_n14423_5865.n33 4.517
R4654 a_n14423_5865.n124 a_n14423_5865.n121 4.517
R4655 a_n14423_5865.n63 a_n14423_5865.n62 4.5
R4656 a_n14423_5865.n2 a_n14423_5865.n1 4.5
R4657 a_n14423_5865.n31 a_n14423_5865.n30 4.314
R4658 a_n14423_5865.n141 a_n14423_5865.n140 4.141
R4659 a_n14423_5865.n51 a_n14423_5865.n50 4.141
R4660 a_n14423_5865.n138 a_n14423_5865.n137 3.944
R4661 a_n14423_5865.n123 a_n14423_5865.n122 3.937
R4662 a_n14423_5865.n53 a_n14423_5865.n52 3.567
R4663 a_n14423_5865.n98 a_n14423_5865.n97 3.395
R4664 a_n14423_5865.n110 a_n14423_5865.n109 3.033
R4665 a_n14423_5865.t3 a_n14423_5865.n151 2.9
R4666 a_n14423_5865.n142 a_n14423_5865.n141 2.258
R4667 a_n14423_5865.n54 a_n14423_5865.n51 2.258
R4668 a_n14423_5865.n99 a_n14423_5865.n98 2.146
R4669 a_n14423_5865.n33 a_n14423_5865.n32 1.882
R4670 a_n14423_5865.n121 a_n14423_5865.n120 1.882
R4671 a_n14423_5865.n54 a_n14423_5865.n53 1.505
R4672 a_n14423_5865.n82 a_n14423_5865.n103 1.5
R4673 a_n14423_5865.n64 a_n14423_5865.n66 1.5
R4674 a_n14423_5865.n63 a_n14423_5865.n61 1.5
R4675 a_n14423_5865.n21 a_n14423_5865.n24 1.5
R4676 a_n14423_5865.n12 a_n14423_5865.n11 1.5
R4677 a_n14423_5865.n109 a_n14423_5865.n80 1.5
R4678 a_n14423_5865.n28 a_n14423_5865.n27 1.129
R4679 a_n14423_5865.n26 a_n14423_5865.n25 1.129
R4680 a_n14423_5865.n142 a_n14423_5865.n138 1.129
R4681 a_n14423_5865.n140 a_n14423_5865.n139 1.129
R4682 a_n14423_5865.n98 a_n14423_5865.n96 1.029
R4683 a_n14423_5865.n102 a_n14423_5865.n101 0.853
R4684 a_n14423_5865.n150 a_n14423_5865.n149 0.752
R4685 a_n14423_5865.n46 a_n14423_5865.n45 0.752
R4686 a_n14423_5865.n49 a_n14423_5865.n48 0.752
R4687 a_n14423_5865.n124 a_n14423_5865.n123 0.752
R4688 a_n14423_5865.n116 a_n14423_5865.n115 0.752
R4689 a_n14423_5865.n118 a_n14423_5865.n117 0.752
R4690 a_n14423_5865.n114 a_n14423_5865.n113 0.752
R4691 a_n14423_5865.n89 a_n14423_5865.n88 0.716
R4692 a_n14423_5865.n131 a_n14423_5865.n130 0.536
R4693 a_n14423_5865.n44 a_n14423_5865.n43 0.536
R4694 a_n14423_5865.n127 a_n14423_5865.n126 0.476
R4695 a_n14423_5865.n39 a_n14423_5865.n38 0.475
R4696 a_n14423_5865.n111 a_n14423_5865.n110 0.382
R4697 a_n14423_5865.n147 a_n14423_5865.n146 0.382
R4698 a_n14423_5865.n146 a_n14423_5865.n145 0.376
R4699 a_n14423_5865.n144 a_n14423_5865.n143 0.376
R4700 a_n14423_5865.n34 a_n14423_5865.n31 0.376
R4701 a_n14423_5865.n38 a_n14423_5865.n37 0.376
R4702 a_n14423_5865.n36 a_n14423_5865.n35 0.376
R4703 a_n14423_5865.n136 a_n14423_5865.n133 0.376
R4704 a_n14423_5865.n135 a_n14423_5865.n134 0.376
R4705 a_n14423_5865.n42 a_n14423_5865.n41 0.376
R4706 a_n14423_5865.n129 a_n14423_5865.n128 0.376
R4707 a_n14423_5865.n119 a_n14423_5865.n118 0.35
R4708 a_n14423_5865.n29 a_n14423_5865.n28 0.349
R4709 a_n14423_5865.n96 a_n14423_5865.n95 0.308
R4710 a_n14423_5865.n2 a_n14423_5865.n0 0.066
R4711 a_n14423_5865.n87 a_n14423_5865.n86 0.047
R4712 a_n14423_5865.n72 a_n14423_5865.n71 0.043
R4713 a_n14423_5865.n68 a_n14423_5865.n67 0.043
R4714 a_n14423_5865.n64 a_n14423_5865.n63 0.041
R4715 a_n14423_5865.n79 a_n14423_5865.n78 0.035
R4716 a_n14423_5865.n108 a_n14423_5865.n107 0.035
R4717 a_n14423_5865.n19 a_n14423_5865.n18 0.034
R4718 a_n14423_5865.n23 a_n14423_5865.n22 0.034
R4719 a_n14423_5865.n8 a_n14423_5865.n7 0.034
R4720 a_n14423_5865.n77 a_n14423_5865.n76 0.034
R4721 a_n14423_5865.n106 a_n14423_5865.n105 0.034
R4722 a_n14423_5865.n12 a_n14423_5865.n6 0.032
R4723 a_n14423_5865.n109 a_n14423_5865.n70 0.032
R4724 a_n14423_5865.n100 a_n14423_5865.n99 0.031
R4725 a_n14423_5865.n9 a_n14423_5865.n8 0.03
R4726 a_n14423_5865.n75 a_n14423_5865.n74 0.03
R4727 a_n14423_5865.n102 a_n14423_5865.n94 0.03
R4728 a_n14423_5865.n81 a_n14423_5865.n87 0.03
R4729 a_n14423_5865.n11 a_n14423_5865.n10 0.028
R4730 a_n14423_5865.n60 a_n14423_5865.n58 0.028
R4731 a_n14423_5865.n73 a_n14423_5865.n72 0.028
R4732 a_n14423_5865.n91 a_n14423_5865.n90 0.028
R4733 a_n14423_5865.n13 a_n14423_5865.n12 0.028
R4734 a_n14423_5865.n57 a_n14423_5865.n56 0.028
R4735 a_n14423_5865.n69 a_n14423_5865.n68 0.028
R4736 a_n14423_5865.n104 a_n14423_5865.n82 0.028
R4737 a_n14423_5865.n85 a_n14423_5865.n83 0.028
R4738 a_n14423_5865.n17 a_n14423_5865.n15 0.026
R4739 a_n14423_5865.n66 a_n14423_5865.n65 0.026
R4740 a_n14423_5865.n93 a_n14423_5865.n92 0.026
R4741 a_n14423_5865.n4 a_n14423_5865.n3 0.026
R4742 a_n14423_5865.n90 a_n14423_5865.n89 0.024
R4743 a_n14423_5865.n18 a_n14423_5865.n17 0.024
R4744 a_n14423_5865.n6 a_n14423_5865.n5 0.024
R4745 a_n14423_5865.n15 a_n14423_5865.n16 0.022
R4746 a_n14423_5865.n5 a_n14423_5865.n4 0.022
R4747 a_n14423_5865.n3 a_n14423_5865.n2 0.022
R4748 a_n14423_5865.n20 a_n14423_5865.n19 0.02
R4749 a_n14423_5865.n10 a_n14423_5865.n9 0.02
R4750 a_n14423_5865.n94 a_n14423_5865.n93 0.02
R4751 a_n14423_5865.n14 a_n14423_5865.n13 0.02
R4752 a_n14423_5865.n101 a_n14423_5865.n100 0.019
R4753 a_n14423_5865.n82 a_n14423_5865.n81 0.018
R4754 a_n14423_5865.n103 a_n14423_5865.n102 0.018
R4755 a_n14423_5865.n70 a_n14423_5865.n69 0.018
R4756 a_n14423_5865.n24 a_n14423_5865.n23 0.017
R4757 a_n14423_5865.n74 a_n14423_5865.n73 0.017
R4758 a_n14423_5865.n58 a_n14423_5865.n59 0.015
R4759 a_n14423_5865.n61 a_n14423_5865.n60 0.015
R4760 a_n14423_5865.n56 a_n14423_5865.n0 0.015
R4761 a_n14423_5865.n63 a_n14423_5865.n57 0.015
R4762 a_n14423_5865.n80 a_n14423_5865.n79 0.013
R4763 a_n14423_5865.n78 a_n14423_5865.n77 0.013
R4764 a_n14423_5865.n109 a_n14423_5865.n108 0.013
R4765 a_n14423_5865.n107 a_n14423_5865.n106 0.013
R4766 a_n14423_5865.n92 a_n14423_5865.n91 0.007
R4767 a_n14423_5865.n86 a_n14423_5865.n85 0.007
R4768 a_n14423_5865.n21 a_n14423_5865.n20 1.424
R4769 a_n14423_5865.n67 a_n14423_5865.n64 0.005
R4770 a_n14423_5865.n80 a_n14423_5865.n75 0.003
R4771 a_n14423_5865.n105 a_n14423_5865.n104 0.003
R4772 a_n14423_5865.n83 a_n14423_5865.n84 0.003
R4773 a_n14423_5865.n14 a_n14423_5865.n21 0.47
R4774 fout6.n510 fout6.t5 1038.95
R4775 fout6.n388 fout6.t11 1037.29
R4776 fout6.n389 fout6.t10 798.832
R4777 fout6.n525 fout6.t14 795.565
R4778 fout6.n367 fout6.t4 732.329
R4779 fout6.n472 fout6.t9 731.671
R4780 fout6.n457 fout6.t13 731.671
R4781 fout6.n497 fout6.t8 730.672
R4782 fout6.n496 fout6.t7 400.616
R4783 fout6.n466 fout6.t12 400.613
R4784 fout6.n11 fout6.t3 397.313
R4785 fout6.n497 fout6.t6 395.84
R4786 fout6.n244 fout6.n243 13.176
R4787 fout6.n14 fout6.t0 11.731
R4788 fout6.n14 fout6.t1 10.988
R4789 fout6.n23 fout6.n22 9.3
R4790 fout6.n322 fout6.n321 9.3
R4791 fout6.n288 fout6.n287 9.3
R4792 fout6.n285 fout6.n284 9.3
R4793 fout6.n222 fout6.n221 9.3
R4794 fout6.n336 fout6.n335 9.3
R4795 fout6.n338 fout6.n337 9.3
R4796 fout6.n220 fout6.n219 9.3
R4797 fout6.n253 fout6.n252 9.3
R4798 fout6.n266 fout6.n265 9.3
R4799 fout6.n274 fout6.n273 9.3
R4800 fout6.n277 fout6.n276 9.3
R4801 fout6.n137 fout6.n136 9.3
R4802 fout6.n134 fout6.n133 9.3
R4803 fout6.n50 fout6.n49 9.3
R4804 fout6.n48 fout6.n47 9.3
R4805 fout6.n41 fout6.n40 8.097
R4806 fout6.n276 fout6.n275 5.457
R4807 fout6.n136 fout6.n135 5.08
R4808 fout6.n39 fout6.n38 4.65
R4809 fout6.n146 fout6.n145 4.65
R4810 fout6.n55 fout6.n53 4.5
R4811 fout6.n107 fout6.n103 4.5
R4812 fout6.n111 fout6.n100 4.5
R4813 fout6.n126 fout6.n125 4.5
R4814 fout6.n81 fout6.n80 4.5
R4815 fout6.n255 fout6.n247 4.5
R4816 fout6.n262 fout6.n245 4.5
R4817 fout6.n271 fout6.n242 4.5
R4818 fout6.n294 fout6.n293 4.5
R4819 fout6.n342 fout6.n341 4.5
R4820 fout6.n330 fout6.n329 4.5
R4821 fout6.n230 fout6.n229 4.5
R4822 fout6.n237 fout6.n236 4.5
R4823 fout6.n302 fout6.n301 4.5
R4824 fout6.n282 fout6.n281 4.5
R4825 fout6.n119 fout6.n118 4.5
R4826 fout6.n213 fout6.n212 4.5
R4827 fout6.n27 fout6.n25 4.5
R4828 fout6.n229 fout6.n227 4.314
R4829 fout6.n301 fout6.n298 3.944
R4830 fout6.n103 fout6.n102 3.937
R4831 fout6.n118 fout6.n117 3.567
R4832 fout6.n147 fout6.n140 3.033
R4833 fout6.n43 fout6.n42 3.033
R4834 fout6.n40 fout6.t2 2.9
R4835 fout6.n300 fout6.n299 2.258
R4836 fout6.n116 fout6.n115 2.258
R4837 fout6.n235 fout6.n234 1.882
R4838 fout6.n236 fout6.n235 1.882
R4839 fout6.n99 fout6.n98 1.882
R4840 fout6.n350 fout6.n14 1.64
R4841 fout6.n118 fout6.n116 1.505
R4842 fout6.n100 fout6.n99 1.505
R4843 fout6.n56 fout6.n55 1.5
R4844 fout6.n343 fout6.n342 1.5
R4845 fout6.n82 fout6.n81 1.5
R4846 fout6.n148 fout6.n147 1.5
R4847 fout6.n127 fout6.n126 1.5
R4848 fout6.n214 fout6.n213 1.5
R4849 fout6.n28 fout6.n27 1.5
R4850 fout6.n422 fout6.n421 1.435
R4851 fout6.n440 fout6.n439 1.435
R4852 fout6.n402 fout6.n388 1.388
R4853 fout6.n527 fout6.n525 1.354
R4854 fout6.n511 fout6.n510 1.354
R4855 fout6.n390 fout6.n389 1.354
R4856 fout6.n474 fout6.n472 1.354
R4857 fout6.n369 fout6.n367 1.354
R4858 fout6.n459 fout6.n457 1.354
R4859 fout6.n12 fout6.n11 1.354
R4860 fout6.n460 fout6.n459 1.142
R4861 fout6.n528 fout6.n527 1.142
R4862 fout6.n423 fout6.n422 1.142
R4863 fout6.n441 fout6.n440 1.142
R4864 fout6.n13 fout6.n12 1.142
R4865 fout6.n483 fout6.n423 1.138
R4866 fout6.n463 fout6.n441 1.138
R4867 fout6.n463 fout6.n460 1.138
R4868 fout6.n529 fout6.n528 1.138
R4869 fout6.n362 fout6.n13 1.138
R4870 fout6.n512 fout6.n511 1.137
R4871 fout6.n538 fout6.n537 1.137
R4872 fout6.n503 fout6.n502 1.137
R4873 fout6.n533 fout6.n532 1.137
R4874 fout6.n518 fout6.n517 1.137
R4875 fout6.n492 fout6.n491 1.137
R4876 fout6.n479 fout6.n478 1.137
R4877 fout6.n487 fout6.n486 1.137
R4878 fout6.n414 fout6.n413 1.137
R4879 fout6.n475 fout6.n474 1.137
R4880 fout6.n426 fout6.n425 1.137
R4881 fout6.n444 fout6.n443 1.137
R4882 fout6.n432 fout6.n431 1.137
R4883 fout6.n450 fout6.n449 1.137
R4884 fout6.n359 fout6.n358 1.137
R4885 fout6.n375 fout6.n374 1.137
R4886 fout6.n355 fout6.n354 1.137
R4887 fout6.n3 fout6.n2 1.137
R4888 fout6.n370 fout6.n369 1.137
R4889 fout6.n540 fout6.n539 1.136
R4890 fout6.n482 fout6.n481 1.136
R4891 fout6.n494 fout6.n493 1.136
R4892 fout6.n514 fout6.n513 1.136
R4893 fout6.n378 fout6.n377 1.136
R4894 fout6.n361 fout6.n360 1.136
R4895 fout6.n341 fout6.n340 1.129
R4896 fout6.n301 fout6.n300 1.129
R4897 fout6.n293 fout6.n292 1.129
R4898 fout6.n303 fout6.n302 1.042
R4899 fout6.n58 fout6.n57 0.853
R4900 fout6.n192 fout6.n191 0.853
R4901 fout6.n150 fout6.n149 0.853
R4902 fout6.n345 fout6.n344 0.853
R4903 fout6.n410 fout6.n409 0.826
R4904 fout6.n212 fout6.n211 0.752
R4905 fout6.n80 fout6.n79 0.752
R4906 fout6.n125 fout6.n124 0.752
R4907 fout6.n103 fout6.n101 0.752
R4908 fout6.n53 fout6.n52 0.752
R4909 fout6.n25 fout6.n24 0.752
R4910 fout6.n30 fout6.n29 0.716
R4911 fout6.n350 fout6.n349 0.69
R4912 fout6.n351 fout6.n350 0.68
R4913 fout6.n252 fout6.n251 0.536
R4914 fout6.n265 fout6.n264 0.536
R4915 fout6.n145 fout6.n144 0.476
R4916 fout6.n287 fout6.n286 0.475
R4917 fout6.n410 fout6.n379 0.471
R4918 fout6.n403 fout6.n402 0.44
R4919 fout6.n42 fout6.n41 0.382
R4920 fout6.n328 fout6.n327 0.382
R4921 fout6.n329 fout6.n328 0.376
R4922 fout6.n229 fout6.n228 0.376
R4923 fout6.n281 fout6.n280 0.376
R4924 fout6.n242 fout6.n241 0.376
R4925 fout6.n245 fout6.n244 0.376
R4926 fout6.n247 fout6.n246 0.376
R4927 fout6.n52 fout6.n51 0.35
R4928 fout6.n340 fout6.n339 0.349
R4929 fout6 fout6.n541 0.176
R4930 fout6.n499 fout6.n498 0.152
R4931 fout6.n496 fout6.n495 0.123
R4932 fout6.n466 fout6.n465 0.123
R4933 fout6 fout6.n410 0.094
R4934 fout6.n467 fout6.n466 0.091
R4935 fout6.n472 fout6.n471 0.083
R4936 fout6.n457 fout6.n456 0.083
R4937 fout6.n367 fout6.n366 0.083
R4938 fout6.n11 fout6.n10 0.083
R4939 fout6.n525 fout6.n524 0.076
R4940 fout6.n510 fout6.n509 0.076
R4941 fout6.n388 fout6.n387 0.076
R4942 fout6.n498 fout6.n496 0.07
R4943 fout6.n384 fout6.n383 0.059
R4944 fout6.n324 fout6.n323 0.047
R4945 fout6.n278 fout6.n277 0.047
R4946 fout6.n268 fout6.n267 0.047
R4947 fout6.n259 fout6.n258 0.047
R4948 fout6.n249 fout6.n248 0.047
R4949 fout6.n138 fout6.n137 0.047
R4950 fout6.n21 fout6.n20 0.047
R4951 fout6.n106 fout6.n105 0.043
R4952 fout6.n88 fout6.n87 0.043
R4953 fout6.n226 fout6.n225 0.041
R4954 fout6.n311 fout6.n310 0.041
R4955 fout6.n45 fout6.n44 0.035
R4956 fout6.n181 fout6.n180 0.035
R4957 fout6.n176 fout6.n175 0.035
R4958 fout6.n35 fout6.n34 0.035
R4959 fout6.n333 fout6.n332 0.034
R4960 fout6.n261 fout6.n260 0.034
R4961 fout6.n257 fout6.n256 0.034
R4962 fout6.n48 fout6.n46 0.034
R4963 fout6.n320 fout6.n319 0.034
R4964 fout6.n318 fout6.n317 0.034
R4965 fout6.n170 fout6.n169 0.034
R4966 fout6.n189 fout6.n188 0.034
R4967 fout6.n82 fout6.n75 0.034
R4968 fout6.n84 fout6.n83 0.034
R4969 fout6.n132 fout6.n131 0.034
R4970 fout6.n37 fout6.n36 0.034
R4971 fout6.n537 fout6.n535 0.032
R4972 fout6.n491 fout6.n489 0.032
R4973 fout6.n443 fout6.n442 0.032
R4974 fout6.n336 fout6.n334 0.032
R4975 fout6.n147 fout6.n146 0.032
R4976 fout6.n43 fout6.n39 0.032
R4977 fout6.n187 fout6.n186 0.032
R4978 fout6.n56 fout6.n37 0.032
R4979 fout6.n354 fout6.n353 0.032
R4980 fout6.n397 fout6.n396 0.032
R4981 fout6.n398 fout6.n397 0.032
R4982 fout6.n402 fout6.n401 0.032
R4983 fout6.n71 fout6.n70 0.031
R4984 fout6.n60 fout6.n59 0.031
R4985 fout6.n347 fout6.n346 0.031
R4986 fout6.n205 fout6.n204 0.031
R4987 fout6.n285 fout6.n283 0.03
R4988 fout6.n270 fout6.n269 0.03
R4989 fout6.n77 fout6.n76 0.03
R4990 fout6.n20 fout6.n19 0.03
R4991 fout6.n343 fout6.n320 0.03
R4992 fout6.n315 fout6.n314 0.03
R4993 fout6.n185 fout6.n184 0.03
R4994 fout6.n73 fout6.n72 0.03
R4995 fout6.n85 fout6.n84 0.03
R4996 fout6.n32 fout6.n31 0.03
R4997 fout6.n194 fout6.n193 0.03
R4998 fout6.n163 fout6.n162 0.03
R4999 fout6.n152 fout6.n151 0.03
R5000 fout6.n392 fout6.n391 0.03
R5001 fout6.n517 fout6.n516 0.028
R5002 fout6.n532 fout6.n531 0.028
R5003 fout6.n537 fout6.n536 0.028
R5004 fout6.n502 fout6.n500 0.028
R5005 fout6.n471 fout6.n470 0.028
R5006 fout6.n469 fout6.n468 0.028
R5007 fout6.n419 fout6.n418 0.028
R5008 fout6.n421 fout6.n420 0.028
R5009 fout6.n478 fout6.n477 0.028
R5010 fout6.n486 fout6.n485 0.028
R5011 fout6.n491 fout6.n490 0.028
R5012 fout6.n413 fout6.n411 0.028
R5013 fout6.n456 fout6.n455 0.028
R5014 fout6.n454 fout6.n453 0.028
R5015 fout6.n437 fout6.n436 0.028
R5016 fout6.n439 fout6.n438 0.028
R5017 fout6.n449 fout6.n448 0.028
R5018 fout6.n431 fout6.n429 0.028
R5019 fout6.n325 fout6.n324 0.028
R5020 fout6.n224 fout6.n223 0.028
R5021 fout6.n239 fout6.n238 0.028
R5022 fout6.n302 fout6.n240 0.028
R5023 fout6.n291 fout6.n290 0.028
R5024 fout6.n147 fout6.n139 0.028
R5025 fout6.n113 fout6.n112 0.028
R5026 fout6.n105 fout6.n104 0.028
R5027 fout6.n55 fout6.n50 0.028
R5028 fout6.n27 fout6.n23 0.028
R5029 fout6.n215 fout6.n214 0.028
R5030 fout6.n344 fout6.n218 0.028
R5031 fout6.n313 fout6.n312 0.028
R5032 fout6.n306 fout6.n305 0.028
R5033 fout6.n304 fout6.n303 0.028
R5034 fout6.n168 fout6.n167 0.028
R5035 fout6.n190 fout6.n189 0.028
R5036 fout6.n183 fout6.n182 0.028
R5037 fout6.n174 fout6.n173 0.028
R5038 fout6.n149 fout6.n148 0.028
R5039 fout6.n93 fout6.n92 0.028
R5040 fout6.n87 fout6.n86 0.028
R5041 fout6.n28 fout6.n18 0.028
R5042 fout6.n366 fout6.n365 0.028
R5043 fout6.n364 fout6.n363 0.028
R5044 fout6.n8 fout6.n7 0.028
R5045 fout6.n10 fout6.n9 0.028
R5046 fout6.n374 fout6.n373 0.028
R5047 fout6.n354 fout6.n352 0.028
R5048 fout6.n358 fout6.n357 0.028
R5049 fout6.n2 fout6.n0 0.028
R5050 fout6.n394 fout6.n393 0.028
R5051 fout6.n396 fout6.n395 0.028
R5052 fout6.n399 fout6.n398 0.028
R5053 fout6.n401 fout6.n400 0.028
R5054 fout6.n67 fout6.n66 0.027
R5055 fout6.n64 fout6.n63 0.027
R5056 fout6.n524 fout6.n523 0.026
R5057 fout6.n522 fout6.n521 0.026
R5058 fout6.n507 fout6.n506 0.026
R5059 fout6.n509 fout6.n508 0.026
R5060 fout6.n342 fout6.n338 0.026
R5061 fout6.n282 fout6.n279 0.026
R5062 fout6.n142 fout6.n141 0.026
R5063 fout6.n119 fout6.n114 0.026
R5064 fout6.n165 fout6.n164 0.026
R5065 fout6.n191 fout6.n171 0.026
R5066 fout6.n130 fout6.n129 0.026
R5067 fout6.n95 fout6.n94 0.026
R5068 fout6.n90 fout6.n89 0.026
R5069 fout6.n17 fout6.n16 0.026
R5070 fout6.n201 fout6.n200 0.026
R5071 fout6.n198 fout6.n197 0.026
R5072 fout6.n159 fout6.n158 0.026
R5073 fout6.n156 fout6.n155 0.026
R5074 fout6.n381 fout6.n380 0.026
R5075 fout6.n383 fout6.n382 0.026
R5076 fout6.n385 fout6.n384 0.026
R5077 fout6.n387 fout6.n386 0.026
R5078 fout6.n29 fout6.n28 0.024
R5079 fout6.n289 fout6.n288 0.024
R5080 fout6.n146 fout6.n143 0.024
R5081 fout6.n217 fout6.n216 0.024
R5082 fout6.n309 fout6.n308 0.024
R5083 fout6.n171 fout6.n170 0.024
R5084 fout6.n178 fout6.n177 0.024
R5085 fout6.n127 fout6.n97 0.024
R5086 fout6.n406 fout6.n405 0.023
R5087 fout6.n232 fout6.n231 0.022
R5088 fout6.n279 fout6.n278 0.022
R5089 fout6.n266 fout6.n263 0.022
R5090 fout6.n254 fout6.n253 0.022
R5091 fout6.n143 fout6.n142 0.022
R5092 fout6.n109 fout6.n108 0.022
R5093 fout6.n218 fout6.n217 0.022
R5094 fout6.n191 fout6.n190 0.022
R5095 fout6.n179 fout6.n178 0.022
R5096 fout6.n148 fout6.n132 0.022
R5097 fout6.n131 fout6.n130 0.022
R5098 fout6.n296 fout6.n295 0.02
R5099 fout6.n294 fout6.n291 0.02
R5100 fout6.n290 fout6.n289 0.02
R5101 fout6.n139 fout6.n138 0.02
R5102 fout6.n123 fout6.n122 0.02
R5103 fout6.n214 fout6.n208 0.02
R5104 fout6.n344 fout6.n343 0.02
R5105 fout6.n169 fout6.n168 0.02
R5106 fout6.n149 fout6.n85 0.02
R5107 fout6.n16 fout6.n15 0.02
R5108 fout6.n59 fout6.n58 0.019
R5109 fout6.n58 fout6.n30 0.019
R5110 fout6.n346 fout6.n345 0.019
R5111 fout6.n345 fout6.n205 0.019
R5112 fout6.n308 fout6.n307 0.018
R5113 fout6.n57 fout6.n56 0.018
R5114 fout6.n150 fout6.n71 0.018
R5115 fout6.n193 fout6.n192 0.018
R5116 fout6.n192 fout6.n163 0.018
R5117 fout6.n151 fout6.n150 0.018
R5118 fout6.n527 fout6.n526 0.017
R5119 fout6.n517 fout6.n515 0.017
R5120 fout6.n502 fout6.n501 0.017
R5121 fout6.n511 fout6.n505 0.017
R5122 fout6.n474 fout6.n473 0.017
R5123 fout6.n478 fout6.n476 0.017
R5124 fout6.n413 fout6.n412 0.017
R5125 fout6.n422 fout6.n417 0.017
R5126 fout6.n459 fout6.n458 0.017
R5127 fout6.n449 fout6.n446 0.017
R5128 fout6.n431 fout6.n430 0.017
R5129 fout6.n440 fout6.n435 0.017
R5130 fout6.n210 fout6.n209 0.017
R5131 fout6.n223 fout6.n222 0.017
R5132 fout6.n272 fout6.n271 0.017
R5133 fout6.n269 fout6.n268 0.017
R5134 fout6.n208 fout6.n207 0.017
R5135 fout6.n314 fout6.n313 0.017
R5136 fout6.n167 fout6.n166 0.017
R5137 fout6.n188 fout6.n187 0.017
R5138 fout6.n186 fout6.n185 0.017
R5139 fout6.n184 fout6.n183 0.017
R5140 fout6.n129 fout6.n128 0.017
R5141 fout6.n97 fout6.n96 0.017
R5142 fout6.n91 fout6.n90 0.017
R5143 fout6.n369 fout6.n368 0.017
R5144 fout6.n374 fout6.n372 0.017
R5145 fout6.n2 fout6.n1 0.017
R5146 fout6.n12 fout6.n6 0.017
R5147 fout6.n391 fout6.n390 0.017
R5148 fout6.n393 fout6.n392 0.017
R5149 fout6.n533 fout6.n530 0.016
R5150 fout6.n538 fout6.n534 0.016
R5151 fout6.n487 fout6.n484 0.016
R5152 fout6.n492 fout6.n488 0.016
R5153 fout6.n445 fout6.n444 0.016
R5154 fout6.n427 fout6.n426 0.016
R5155 fout6.n359 fout6.n356 0.016
R5156 fout6.n470 fout6.n469 0.015
R5157 fout6.n420 fout6.n419 0.015
R5158 fout6.n455 fout6.n454 0.015
R5159 fout6.n438 fout6.n437 0.015
R5160 fout6.n448 fout6.n447 0.015
R5161 fout6.n429 fout6.n428 0.015
R5162 fout6.n326 fout6.n325 0.015
R5163 fout6.n334 fout6.n333 0.015
R5164 fout6.n240 fout6.n239 0.015
R5165 fout6.n81 fout6.n78 0.015
R5166 fout6.n114 fout6.n113 0.015
R5167 fout6.n112 fout6.n111 0.015
R5168 fout6.n319 fout6.n318 0.015
R5169 fout6.n317 fout6.n316 0.015
R5170 fout6.n305 fout6.n304 0.015
R5171 fout6.n75 fout6.n74 0.015
R5172 fout6.n83 fout6.n82 0.015
R5173 fout6.n94 fout6.n93 0.015
R5174 fout6.n92 fout6.n91 0.015
R5175 fout6.n365 fout6.n364 0.015
R5176 fout6.n9 fout6.n8 0.015
R5177 fout6.n395 fout6.n394 0.015
R5178 fout6.n400 fout6.n399 0.015
R5179 fout6.n523 fout6.n522 0.013
R5180 fout6.n508 fout6.n507 0.013
R5181 fout6.n332 fout6.n331 0.013
R5182 fout6.n238 fout6.n237 0.013
R5183 fout6.n274 fout6.n272 0.013
R5184 fout6.n44 fout6.n43 0.013
R5185 fout6.n46 fout6.n45 0.013
R5186 fout6.n307 fout6.n306 0.013
R5187 fout6.n34 fout6.n33 0.013
R5188 fout6.n36 fout6.n35 0.013
R5189 fout6.n349 fout6.n348 0.013
R5190 fout6.n382 fout6.n381 0.013
R5191 fout6.n386 fout6.n385 0.013
R5192 fout6.n539 fout6.n533 0.012
R5193 fout6.n539 fout6.n538 0.012
R5194 fout6.n493 fout6.n487 0.012
R5195 fout6.n493 fout6.n492 0.012
R5196 fout6.n426 fout6.n424 0.012
R5197 fout6.n66 fout6.n65 0.012
R5198 fout6.n65 fout6.n64 0.012
R5199 fout6.n360 fout6.n355 0.012
R5200 fout6.n360 fout6.n359 0.012
R5201 fout6.n520 fout6.n519 0.011
R5202 fout6.n513 fout6.n504 0.011
R5203 fout6.n481 fout6.n480 0.011
R5204 fout6.n416 fout6.n415 0.011
R5205 fout6.n452 fout6.n451 0.011
R5206 fout6.n434 fout6.n433 0.011
R5207 fout6.n297 fout6.n296 0.011
R5208 fout6.n122 fout6.n121 0.011
R5209 fout6.n69 fout6.n68 0.011
R5210 fout6.n62 fout6.n61 0.011
R5211 fout6.n200 fout6.n199 0.011
R5212 fout6.n199 fout6.n198 0.011
R5213 fout6.n196 fout6.n195 0.011
R5214 fout6.n161 fout6.n160 0.011
R5215 fout6.n158 fout6.n157 0.011
R5216 fout6.n157 fout6.n156 0.011
R5217 fout6.n154 fout6.n153 0.011
R5218 fout6.n203 fout6.n202 0.011
R5219 fout6.n377 fout6.n376 0.011
R5220 fout6.n5 fout6.n4 0.011
R5221 fout6.n450 fout6.n445 0.01
R5222 fout6.n432 fout6.n427 0.01
R5223 fout6.n375 fout6.n371 0.01
R5224 fout6.n405 fout6.n404 0.01
R5225 fout6.n404 fout6.n403 0.01
R5226 fout6.n323 fout6.n322 0.009
R5227 fout6.n233 fout6.n232 0.009
R5228 fout6.n237 fout6.n233 0.009
R5229 fout6.n260 fout6.n259 0.009
R5230 fout6.n110 fout6.n109 0.009
R5231 fout6.n216 fout6.n215 0.009
R5232 fout6.n180 fout6.n179 0.009
R5233 fout6.n408 fout6.n407 0.009
R5234 fout6.n230 fout6.n226 0.007
R5235 fout6.n263 fout6.n262 0.007
R5236 fout6.n258 fout6.n257 0.007
R5237 fout6.n255 fout6.n254 0.007
R5238 fout6.n111 fout6.n110 0.007
R5239 fout6.n23 fout6.n21 0.007
R5240 fout6.n310 fout6.n309 0.007
R5241 fout6.n182 fout6.n181 0.007
R5242 fout6.n177 fout6.n176 0.007
R5243 fout6.n175 fout6.n174 0.007
R5244 fout6.n18 fout6.n17 0.007
R5245 fout6.n519 fout6.n518 0.006
R5246 fout6.n504 fout6.n503 0.006
R5247 fout6.n513 fout6.n512 0.006
R5248 fout6.n481 fout6.n475 0.006
R5249 fout6.n480 fout6.n479 0.006
R5250 fout6.n415 fout6.n414 0.006
R5251 fout6.n451 fout6.n450 0.006
R5252 fout6.n433 fout6.n432 0.006
R5253 fout6.n70 fout6.n69 0.006
R5254 fout6.n68 fout6.n67 0.006
R5255 fout6.n63 fout6.n62 0.006
R5256 fout6.n61 fout6.n60 0.006
R5257 fout6.n197 fout6.n196 0.006
R5258 fout6.n195 fout6.n194 0.006
R5259 fout6.n162 fout6.n161 0.006
R5260 fout6.n160 fout6.n159 0.006
R5261 fout6.n155 fout6.n154 0.006
R5262 fout6.n153 fout6.n152 0.006
R5263 fout6.n348 fout6.n347 0.006
R5264 fout6.n204 fout6.n203 0.006
R5265 fout6.n202 fout6.n201 0.006
R5266 fout6.n377 fout6.n370 0.006
R5267 fout6.n376 fout6.n375 0.006
R5268 fout6.n4 fout6.n3 0.006
R5269 fout6.n342 fout6.n326 0.005
R5270 fout6.n338 fout6.n336 0.005
R5271 fout6.n302 fout6.n297 0.005
R5272 fout6.n295 fout6.n294 0.005
R5273 fout6.n267 fout6.n266 0.005
R5274 fout6.n253 fout6.n250 0.005
R5275 fout6.n121 fout6.n120 0.005
R5276 fout6.n107 fout6.n106 0.005
R5277 fout6.n207 fout6.n206 0.005
R5278 fout6.n128 fout6.n127 0.005
R5279 fout6.n89 fout6.n88 0.005
R5280 fout6.n409 fout6.n408 0.005
R5281 fout6.n407 fout6.n406 0.005
R5282 fout6.n541 fout6.n540 0.004
R5283 fout6.n514 fout6.n499 0.003
R5284 fout6.n495 fout6.n494 0.003
R5285 fout6.n482 fout6.n467 0.003
R5286 fout6.n361 fout6.n351 0.003
R5287 fout6.n379 fout6.n378 0.003
R5288 fout6.n213 fout6.n210 0.003
R5289 fout6.n81 fout6.n77 0.003
R5290 fout6.n137 fout6.n134 0.003
R5291 fout6.n126 fout6.n123 0.003
R5292 fout6.n108 fout6.n107 0.003
R5293 fout6.n50 fout6.n48 0.003
R5294 fout6.n55 fout6.n54 0.003
R5295 fout6.n27 fout6.n26 0.003
R5296 fout6.n166 fout6.n165 0.003
R5297 fout6.n33 fout6.n32 0.003
R5298 fout6.n528 fout6.n520 0.003
R5299 fout6.n460 fout6.n452 0.003
R5300 fout6.n423 fout6.n416 0.003
R5301 fout6.n441 fout6.n434 0.003
R5302 fout6.n13 fout6.n5 0.003
R5303 fout6.n464 fout6.n463 0.002
R5304 fout6.n462 fout6.n461 0.002
R5305 fout6.n465 fout6.n464 0.002
R5306 fout6.n463 fout6.n462 0.002
R5307 fout6.n540 fout6.n529 0.002
R5308 fout6.n483 fout6.n482 0.002
R5309 fout6.n494 fout6.n483 0.002
R5310 fout6.n529 fout6.n514 0.002
R5311 fout6.n378 fout6.n362 0.002
R5312 fout6.n362 fout6.n361 0.002
R5313 fout6.n331 fout6.n330 0.001
R5314 fout6.n222 fout6.n220 0.001
R5315 fout6.n225 fout6.n224 0.001
R5316 fout6.n231 fout6.n230 0.001
R5317 fout6.n288 fout6.n285 0.001
R5318 fout6.n283 fout6.n282 0.001
R5319 fout6.n277 fout6.n274 0.001
R5320 fout6.n271 fout6.n270 0.001
R5321 fout6.n262 fout6.n261 0.001
R5322 fout6.n256 fout6.n255 0.001
R5323 fout6.n250 fout6.n249 0.001
R5324 fout6.n120 fout6.n119 0.001
R5325 fout6.n316 fout6.n315 0.001
R5326 fout6.n312 fout6.n311 0.001
R5327 fout6.n173 fout6.n172 0.001
R5328 fout6.n74 fout6.n73 0.001
R5329 fout6.n96 fout6.n95 0.001
R5330 fout6.n498 fout6.n497 0.001
R5331 fin fin.t4 1038.73
R5332 fin.n121 fin.t0 795.567
R5333 fin.n80 fin.t5 731.671
R5334 fin.n51 fin.t3 731.671
R5335 fin.n14 fin.t2 730.672
R5336 fin.n100 fin.t1 400.619
R5337 fin.n57 fin.t6 400.618
R5338 fin.n14 fin.t7 395.84
R5339 fin.n89 fin.n87 1.435
R5340 fin.n22 fin.n21 1.435
R5341 fin.n130 fin.n120 1.354
R5342 fin.n81 fin.n80 1.354
R5343 fin.n52 fin.n51 1.354
R5344 fin.n82 fin.n81 1.142
R5345 fin.n23 fin.n22 1.14
R5346 fin.n83 fin.n82 1.138
R5347 fin.n90 fin.n89 1.137
R5348 fin.n66 fin.n65 1.137
R5349 fin.n72 fin.n71 1.137
R5350 fin.n61 fin.n60 1.137
R5351 fin.n95 fin.n94 1.137
R5352 fin.n28 fin.n27 1.137
R5353 fin.n33 fin.n32 1.137
R5354 fin.n53 fin.n52 1.137
R5355 fin.n43 fin.n42 1.137
R5356 fin.n37 fin.n36 1.137
R5357 fin.n120 fin.n119 1.137
R5358 fin.n68 fin.n67 1.136
R5359 fin.n55 fin.n54 1.136
R5360 fin.n118 fin.n106 1.136
R5361 fin.n98 fin.n97 1.136
R5362 fin fin.n130 0.225
R5363 fin.n102 fin.n101 0.154
R5364 fin.n57 fin.n56 0.123
R5365 fin.n100 fin.n99 0.123
R5366 fin.n58 fin.n57 0.091
R5367 fin.n80 fin.n79 0.083
R5368 fin.n51 fin.n50 0.083
R5369 fin.n130 fin.n129 0.076
R5370 fin.n122 fin.n121 0.076
R5371 fin.n101 fin.n100 0.072
R5372 fin.n47 fin.n46 0.064
R5373 fin.n126 fin.n125 0.059
R5374 fin.n65 fin.n63 0.032
R5375 fin.n36 fin.n35 0.032
R5376 fin.n8 fin.n7 0.032
R5377 fin.n7 fin.n6 0.032
R5378 fin.n13 fin.n12 0.03
R5379 fin.n2 fin.n1 0.03
R5380 fin.n87 fin.n86 0.028
R5381 fin.n85 fin.n84 0.028
R5382 fin.n77 fin.n76 0.028
R5383 fin.n79 fin.n78 0.028
R5384 fin.n94 fin.n93 0.028
R5385 fin.n60 fin.n59 0.028
R5386 fin.n65 fin.n64 0.028
R5387 fin.n71 fin.n69 0.028
R5388 fin.n21 fin.n20 0.028
R5389 fin.n48 fin.n47 0.028
R5390 fin.n50 fin.n49 0.028
R5391 fin.n32 fin.n31 0.028
R5392 fin.n42 fin.n40 0.028
R5393 fin.n11 fin.n10 0.028
R5394 fin.n9 fin.n8 0.028
R5395 fin.n6 fin.n5 0.028
R5396 fin.n4 fin.n3 0.028
R5397 fin.n129 fin.n128 0.026
R5398 fin.n127 fin.n126 0.026
R5399 fin.n125 fin.n124 0.026
R5400 fin.n123 fin.n122 0.026
R5401 fin.n89 fin.n88 0.017
R5402 fin.n94 fin.n92 0.017
R5403 fin.n71 fin.n70 0.017
R5404 fin.n81 fin.n75 0.017
R5405 fin.n22 fin.n18 0.017
R5406 fin.n27 fin.n26 0.017
R5407 fin.n42 fin.n41 0.017
R5408 fin.n52 fin.n45 0.017
R5409 fin.n120 fin.n13 0.017
R5410 fin.n12 fin.n11 0.017
R5411 fin.n3 fin.n2 0.017
R5412 fin.n1 fin.n0 0.017
R5413 fin.n115 fin.n114 0.016
R5414 fin.n112 fin.n111 0.016
R5415 fin.n66 fin.n62 0.016
R5416 fin.n33 fin.n29 0.016
R5417 fin.n38 fin.n37 0.016
R5418 fin.n86 fin.n85 0.015
R5419 fin.n78 fin.n77 0.015
R5420 fin.n20 fin.n19 0.015
R5421 fin.n49 fin.n48 0.015
R5422 fin.n31 fin.n30 0.015
R5423 fin.n40 fin.n39 0.015
R5424 fin.n10 fin.n9 0.015
R5425 fin.n5 fin.n4 0.015
R5426 fin.n128 fin.n127 0.013
R5427 fin.n124 fin.n123 0.013
R5428 fin.n114 fin.n113 0.012
R5429 fin.n113 fin.n112 0.012
R5430 fin.n67 fin.n61 0.012
R5431 fin.n67 fin.n66 0.012
R5432 fin.n34 fin.n33 0.012
R5433 fin.n37 fin.n34 0.012
R5434 fin.n118 fin.n117 0.011
R5435 fin.n109 fin.n108 0.011
R5436 fin.n97 fin.n96 0.011
R5437 fin.n74 fin.n73 0.011
R5438 fin.n25 fin.n24 0.011
R5439 fin.n54 fin.n44 0.011
R5440 fin.n116 fin.n115 0.01
R5441 fin.n111 fin.n110 0.01
R5442 fin.n95 fin.n91 0.01
R5443 fin.n29 fin.n28 0.01
R5444 fin.n43 fin.n38 0.01
R5445 fin.n119 fin.n118 0.006
R5446 fin.n117 fin.n116 0.006
R5447 fin.n110 fin.n109 0.006
R5448 fin.n97 fin.n90 0.006
R5449 fin.n96 fin.n95 0.006
R5450 fin.n73 fin.n72 0.006
R5451 fin.n28 fin.n25 0.006
R5452 fin.n44 fin.n43 0.006
R5453 fin.n54 fin.n53 0.006
R5454 fin.n103 fin.n102 0.004
R5455 fin.n68 fin.n58 0.004
R5456 fin.n24 fin.n23 0.003
R5457 fin.n56 fin.n55 0.003
R5458 fin.n99 fin.n98 0.003
R5459 fin.n106 fin.n105 0.003
R5460 fin.n82 fin.n74 0.003
R5461 fin.n16 fin.n15 0.003
R5462 fin.n108 fin.n107 0.002
R5463 fin.n17 fin.n16 0.002
R5464 fin.n104 fin.n103 0.002
R5465 fin.n83 fin.n68 0.002
R5466 fin.n106 fin.n104 0.002
R5467 fin.n98 fin.n83 0.002
R5468 fin.n55 fin.n17 0.002
R5469 fin.n101 fin.n14 0.002
R5470 a_n24539_11543.n97 a_n24539_11543.t5 1040.28
R5471 a_n24539_11543.n97 a_n24539_11543.t4 796.134
R5472 a_n24539_11543.n50 a_n24539_11543.n49 13.176
R5473 a_n24539_11543.n98 a_n24539_11543.t1 11.611
R5474 a_n24539_11543.n98 a_n24539_11543.t0 11.295
R5475 a_n24539_11543.n99 a_n24539_11543.t3 10.373
R5476 a_n24539_11543.n138 a_n24539_11543.n39 9.3
R5477 a_n24539_11543.n138 a_n24539_11543.n134 9.3
R5478 a_n24539_11543.n138 a_n24539_11543.n128 9.3
R5479 a_n24539_11543.n138 a_n24539_11543.n58 9.3
R5480 a_n24539_11543.n138 a_n24539_11543.n66 9.3
R5481 a_n24539_11543.n138 a_n24539_11543.n123 9.3
R5482 a_n24539_11543.n138 a_n24539_11543.n118 8.47
R5483 a_n24539_11543.n138 a_n24539_11543.n137 8.469
R5484 a_n24539_11543.n138 a_n24539_11543.n115 8.124
R5485 a_n24539_11543.n138 a_n24539_11543.n29 8.124
R5486 a_n24539_11543.n138 a_n24539_11543.n34 8.097
R5487 a_n24539_11543.n138 a_n24539_11543.n110 8.097
R5488 a_n24539_11543.n138 a_n24539_11543.n61 8.016
R5489 a_n24539_11543.n138 a_n24539_11543.n44 8.016
R5490 a_n24539_11543.n138 a_n24539_11543.n53 7.964
R5491 a_n24539_11543.n138 a_n24539_11543.n48 7.964
R5492 a_n24539_11543.n60 a_n24539_11543.n59 6.4
R5493 a_n24539_11543.n109 a_n24539_11543.n67 6.4
R5494 a_n24539_11543.n32 a_n24539_11543.n31 6.023
R5495 a_n24539_11543.n42 a_n24539_11543.n41 6.023
R5496 a_n24539_11543.n128 a_n24539_11543.n127 6.023
R5497 a_n24539_11543.n47 a_n24539_11543.n46 6.023
R5498 a_n24539_11543.n52 a_n24539_11543.n51 6.023
R5499 a_n24539_11543.n136 a_n24539_11543.n135 5.647
R5500 a_n24539_11543.n58 a_n24539_11543.n55 5.647
R5501 a_n24539_11543.n113 a_n24539_11543.n112 5.647
R5502 a_n24539_11543.n117 a_n24539_11543.n116 5.647
R5503 a_n24539_11543.n125 a_n24539_11543.n124 5.457
R5504 a_n24539_11543.n27 a_n24539_11543.n26 5.27
R5505 a_n24539_11543.n57 a_n24539_11543.n56 5.08
R5506 a_n24539_11543.n39 a_n24539_11543.n38 4.517
R5507 a_n24539_11543.n123 a_n24539_11543.n120 4.517
R5508 a_n24539_11543.n75 a_n24539_11543.n74 4.5
R5509 a_n24539_11543.n2 a_n24539_11543.n1 4.5
R5510 a_n24539_11543.n36 a_n24539_11543.n35 4.314
R5511 a_n24539_11543.n133 a_n24539_11543.n132 4.141
R5512 a_n24539_11543.n63 a_n24539_11543.n62 4.141
R5513 a_n24539_11543.n130 a_n24539_11543.n129 3.944
R5514 a_n24539_11543.n122 a_n24539_11543.n121 3.937
R5515 a_n24539_11543.n65 a_n24539_11543.n64 3.567
R5516 a_n24539_11543.n100 a_n24539_11543.n97 3.395
R5517 a_n24539_11543.n109 a_n24539_11543.n108 3.033
R5518 a_n24539_11543.t2 a_n24539_11543.n138 2.9
R5519 a_n24539_11543.n101 a_n24539_11543.n100 2.4
R5520 a_n24539_11543.n134 a_n24539_11543.n133 2.258
R5521 a_n24539_11543.n66 a_n24539_11543.n63 2.258
R5522 a_n24539_11543.n38 a_n24539_11543.n37 1.882
R5523 a_n24539_11543.n120 a_n24539_11543.n119 1.882
R5524 a_n24539_11543.n66 a_n24539_11543.n65 1.505
R5525 a_n24539_11543.n94 a_n24539_11543.n102 1.5
R5526 a_n24539_11543.n76 a_n24539_11543.n78 1.5
R5527 a_n24539_11543.n75 a_n24539_11543.n73 1.5
R5528 a_n24539_11543.n21 a_n24539_11543.n24 1.5
R5529 a_n24539_11543.n12 a_n24539_11543.n11 1.5
R5530 a_n24539_11543.n108 a_n24539_11543.n92 1.5
R5531 a_n24539_11543.n28 a_n24539_11543.n27 1.129
R5532 a_n24539_11543.n26 a_n24539_11543.n25 1.129
R5533 a_n24539_11543.n134 a_n24539_11543.n130 1.129
R5534 a_n24539_11543.n132 a_n24539_11543.n131 1.129
R5535 a_n24539_11543.n100 a_n24539_11543.n99 1.022
R5536 a_n24539_11543.n137 a_n24539_11543.n136 0.752
R5537 a_n24539_11543.n55 a_n24539_11543.n54 0.752
R5538 a_n24539_11543.n58 a_n24539_11543.n57 0.752
R5539 a_n24539_11543.n123 a_n24539_11543.n122 0.752
R5540 a_n24539_11543.n112 a_n24539_11543.n111 0.752
R5541 a_n24539_11543.n114 a_n24539_11543.n113 0.752
R5542 a_n24539_11543.n118 a_n24539_11543.n117 0.752
R5543 a_n24539_11543.n53 a_n24539_11543.n52 0.536
R5544 a_n24539_11543.n48 a_n24539_11543.n47 0.536
R5545 a_n24539_11543.n61 a_n24539_11543.n60 0.475
R5546 a_n24539_11543.n44 a_n24539_11543.n43 0.475
R5547 a_n24539_11543.n34 a_n24539_11543.n33 0.382
R5548 a_n24539_11543.n110 a_n24539_11543.n109 0.382
R5549 a_n24539_11543.n33 a_n24539_11543.n32 0.376
R5550 a_n24539_11543.n31 a_n24539_11543.n30 0.376
R5551 a_n24539_11543.n39 a_n24539_11543.n36 0.376
R5552 a_n24539_11543.n43 a_n24539_11543.n42 0.376
R5553 a_n24539_11543.n41 a_n24539_11543.n40 0.376
R5554 a_n24539_11543.n128 a_n24539_11543.n125 0.376
R5555 a_n24539_11543.n127 a_n24539_11543.n126 0.376
R5556 a_n24539_11543.n46 a_n24539_11543.n45 0.376
R5557 a_n24539_11543.n51 a_n24539_11543.n50 0.376
R5558 a_n24539_11543.n29 a_n24539_11543.n28 0.349
R5559 a_n24539_11543.n115 a_n24539_11543.n114 0.349
R5560 a_n24539_11543.n99 a_n24539_11543.n98 0.316
R5561 a_n24539_11543.n94 a_n24539_11543.n93 0.15
R5562 a_n24539_11543.n101 a_n24539_11543.n95 0.148
R5563 a_n24539_11543.n2 a_n24539_11543.n0 0.066
R5564 a_n24539_11543.n84 a_n24539_11543.n83 0.043
R5565 a_n24539_11543.n80 a_n24539_11543.n79 0.043
R5566 a_n24539_11543.n76 a_n24539_11543.n75 0.041
R5567 a_n24539_11543.n91 a_n24539_11543.n90 0.035
R5568 a_n24539_11543.n107 a_n24539_11543.n106 0.035
R5569 a_n24539_11543.n19 a_n24539_11543.n18 0.034
R5570 a_n24539_11543.n23 a_n24539_11543.n22 0.034
R5571 a_n24539_11543.n8 a_n24539_11543.n7 0.034
R5572 a_n24539_11543.n89 a_n24539_11543.n88 0.034
R5573 a_n24539_11543.n105 a_n24539_11543.n104 0.034
R5574 a_n24539_11543.n12 a_n24539_11543.n6 0.032
R5575 a_n24539_11543.n108 a_n24539_11543.n82 0.032
R5576 a_n24539_11543.n9 a_n24539_11543.n8 0.03
R5577 a_n24539_11543.n87 a_n24539_11543.n86 0.03
R5578 a_n24539_11543.n11 a_n24539_11543.n10 0.028
R5579 a_n24539_11543.n72 a_n24539_11543.n70 0.028
R5580 a_n24539_11543.n85 a_n24539_11543.n84 0.028
R5581 a_n24539_11543.n13 a_n24539_11543.n12 0.028
R5582 a_n24539_11543.n69 a_n24539_11543.n68 0.028
R5583 a_n24539_11543.n81 a_n24539_11543.n80 0.028
R5584 a_n24539_11543.n103 a_n24539_11543.n94 0.028
R5585 a_n24539_11543.n17 a_n24539_11543.n15 0.026
R5586 a_n24539_11543.n78 a_n24539_11543.n77 0.026
R5587 a_n24539_11543.n4 a_n24539_11543.n3 0.026
R5588 a_n24539_11543.n18 a_n24539_11543.n17 0.024
R5589 a_n24539_11543.n6 a_n24539_11543.n5 0.024
R5590 a_n24539_11543.n15 a_n24539_11543.n16 0.022
R5591 a_n24539_11543.n5 a_n24539_11543.n4 0.022
R5592 a_n24539_11543.n3 a_n24539_11543.n2 0.022
R5593 a_n24539_11543.n20 a_n24539_11543.n19 0.02
R5594 a_n24539_11543.n10 a_n24539_11543.n9 0.02
R5595 a_n24539_11543.n14 a_n24539_11543.n13 0.02
R5596 a_n24539_11543.n102 a_n24539_11543.n101 0.018
R5597 a_n24539_11543.n82 a_n24539_11543.n81 0.018
R5598 a_n24539_11543.n24 a_n24539_11543.n23 0.017
R5599 a_n24539_11543.n86 a_n24539_11543.n85 0.017
R5600 a_n24539_11543.n70 a_n24539_11543.n71 0.015
R5601 a_n24539_11543.n73 a_n24539_11543.n72 0.015
R5602 a_n24539_11543.n68 a_n24539_11543.n0 0.015
R5603 a_n24539_11543.n75 a_n24539_11543.n69 0.015
R5604 a_n24539_11543.n92 a_n24539_11543.n91 0.013
R5605 a_n24539_11543.n90 a_n24539_11543.n89 0.013
R5606 a_n24539_11543.n108 a_n24539_11543.n107 0.013
R5607 a_n24539_11543.n106 a_n24539_11543.n105 0.013
R5608 a_n24539_11543.n95 a_n24539_11543.n96 0.007
R5609 a_n24539_11543.n21 a_n24539_11543.n20 1.424
R5610 a_n24539_11543.n79 a_n24539_11543.n76 0.005
R5611 a_n24539_11543.n92 a_n24539_11543.n87 0.003
R5612 a_n24539_11543.n104 a_n24539_11543.n103 0.003
R5613 a_n24539_11543.n14 a_n24539_11543.n21 0.47
R5614 VDD.n536 VDD.t90 423.114
R5615 VDD.n2125 VDD.t186 422.222
R5616 VDD.n1736 VDD.t61 417.901
R5617 VDD.n1017 VDD.t232 386.053
R5618 VDD.n177 VDD.t23 374.317
R5619 VDD.n2939 VDD.t192 353.086
R5620 VDD.t125 VDD.t73 282.098
R5621 VDD.t11 VDD.t228 281.664
R5622 VDD.t173 VDD.t41 244.603
R5623 VDD.t39 VDD.t202 244.603
R5624 VDD.t217 VDD.t111 244.444
R5625 VDD.t144 VDD.t63 244.444
R5626 VDD.t216 VDD.t49 244.444
R5627 VDD.t55 VDD.t1 243.985
R5628 VDD.t143 VDD.t194 243.985
R5629 VDD.t145 VDD.t59 243.985
R5630 VDD.t0 VDD.t148 243.985
R5631 VDD.t213 VDD.t108 243.985
R5632 VDD.t201 VDD.t81 243.985
R5633 VDD.t7 VDD.t183 243.827
R5634 VDD.t162 VDD.t69 243.827
R5635 VDD.t167 VDD.t222 243.827
R5636 VDD.t223 VDD.t236 243.827
R5637 VDD.t215 VDD.t35 243.827
R5638 VDD.t113 VDD.t15 192.1
R5639 VDD.t234 VDD.t208 192.1
R5640 VDD.t25 VDD.t53 192.1
R5641 VDD.t119 VDD.t230 192.1
R5642 VDD.t224 VDD.t190 191.975
R5643 VDD.t133 VDD.t37 191.975
R5644 VDD.t115 VDD.t129 191.975
R5645 VDD.t67 VDD.t178 191.358
R5646 VDD.t208 VDD.t19 189.629
R5647 VDD.t27 VDD.t119 189.629
R5648 VDD.t178 VDD.t226 189.506
R5649 VDD.t15 VDD.t181 189.011
R5650 VDD.t184 VDD.t25 189.011
R5651 VDD.t139 VDD.t224 188.888
R5652 VDD.t131 VDD.t133 188.888
R5653 VDD.t129 VDD.t51 188.888
R5654 VDD.t1 VDD.t11 176.657
R5655 VDD.t169 VDD.t55 176.657
R5656 VDD.t194 VDD.t12 176.657
R5657 VDD.t181 VDD.t143 176.657
R5658 VDD.t59 VDD.t212 176.657
R5659 VDD.t47 VDD.t145 176.657
R5660 VDD.t148 VDD.t85 176.657
R5661 VDD.t29 VDD.t0 176.657
R5662 VDD.t198 VDD.t213 176.657
R5663 VDD.t108 VDD.t184 176.657
R5664 VDD.t81 VDD.t118 176.657
R5665 VDD.t83 VDD.t201 176.657
R5666 VDD.t183 VDD.t139 176.543
R5667 VDD.t98 VDD.t7 176.543
R5668 VDD.t79 VDD.t162 176.543
R5669 VDD.t69 VDD.t99 176.543
R5670 VDD.t222 VDD.t131 176.543
R5671 VDD.t136 VDD.t167 176.543
R5672 VDD.t160 VDD.t223 176.543
R5673 VDD.t236 VDD.t135 176.543
R5674 VDD.t51 VDD.t215 176.543
R5675 VDD.t35 VDD.t128 176.543
R5676 VDD.t41 VDD.t207 176.04
R5677 VDD.t19 VDD.t173 176.04
R5678 VDD.t117 VDD.t39 176.04
R5679 VDD.t202 VDD.t27 176.04
R5680 VDD.t226 VDD.t217 175.925
R5681 VDD.t111 VDD.t180 175.925
R5682 VDD.t152 VDD.t144 175.925
R5683 VDD.t63 VDD.t58 175.925
R5684 VDD.t65 VDD.t216 175.925
R5685 VDD.t49 VDD.t125 175.925
R5686 VDD.t56 VDD.t188 174.187
R5687 VDD.t232 VDD.t17 174.187
R5688 VDD.t207 VDD.n535 174.187
R5689 VDD.t90 VDD.t210 174.187
R5690 VDD.t23 VDD.t196 174.187
R5691 VDD.n2692 VDD.t117 174.187
R5692 VDD.t180 VDD.n1469 174.074
R5693 VDD.t61 VDD.t31 174.074
R5694 VDD.t186 VDD.t137 174.074
R5695 VDD.t192 VDD.t126 174.074
R5696 VDD.t9 VDD.t171 174.074
R5697 VDD.t12 VDD.n1016 173.569
R5698 VDD.n178 VDD.t198 173.569
R5699 VDD.n1737 VDD.t98 173.456
R5700 VDD.n2259 VDD.t136 173.456
R5701 VDD.t128 VDD.n2938 173.456
R5702 VDD.t228 VDD.t56 161.215
R5703 VDD.t210 VDD.t21 161.215
R5704 VDD.t53 VDD.t154 161.215
R5705 VDD.t203 VDD.t67 161.111
R5706 VDD.t190 VDD.t163 161.111
R5707 VDD.t137 VDD.t45 161.111
R5708 VDD.t126 VDD.t88 161.111
R5709 VDD.t109 VDD.t115 161.111
R5710 VDD.t73 VDD.t9 161.111
R5711 VDD.t156 VDD.t113 160.598
R5712 VDD.t17 VDD.t158 160.598
R5713 VDD.t165 VDD.t234 160.598
R5714 VDD.t196 VDD.t100 160.598
R5715 VDD.t230 VDD.t71 160.598
R5716 VDD.t31 VDD.t5 160.493
R5717 VDD.t37 VDD.t92 160.493
R5718 VDD.n1017 VDD.t75 158.127
R5719 VDD.n536 VDD.t96 158.127
R5720 VDD.t43 VDD.n177 158.127
R5721 VDD.t238 VDD.n2691 158.127
R5722 VDD.n1528 VDD.t146 158.024
R5723 VDD.t220 VDD.n1736 158.024
R5724 VDD.t77 VDD.n2125 158.024
R5725 VDD.n2939 VDD.t104 158.024
R5726 VDD.t94 VDD.t156 150.097
R5727 VDD.t199 VDD.t165 150.097
R5728 VDD.t71 VDD.t150 150.097
R5729 VDD.t218 VDD.t203 150
R5730 VDD.t92 VDD.t3 150
R5731 VDD.t174 VDD.t109 150
R5732 VDD.t154 VDD.t102 149.479
R5733 VDD.t163 VDD.t106 149.382
R5734 VDD.t13 VDD.t94 123.537
R5735 VDD.t75 VDD.t13 123.537
R5736 VDD.t205 VDD.t199 123.537
R5737 VDD.t96 VDD.t205 123.537
R5738 VDD.t102 VDD.t86 123.537
R5739 VDD.t86 VDD.t43 123.537
R5740 VDD.t150 VDD.t121 123.537
R5741 VDD.t121 VDD.t238 123.537
R5742 VDD.t146 VDD.t176 123.456
R5743 VDD.t176 VDD.t218 123.456
R5744 VDD.t33 VDD.t220 123.456
R5745 VDD.t106 VDD.t33 123.456
R5746 VDD.t141 VDD.t77 123.456
R5747 VDD.t3 VDD.t141 123.456
R5748 VDD.t104 VDD.t123 123.456
R5749 VDD.t123 VDD.t174 123.456
R5750 VDD.n1016 VDD.t169 117.36
R5751 VDD.n178 VDD.t29 117.36
R5752 VDD.n1469 VDD.t152 117.283
R5753 VDD.n1737 VDD.t79 117.283
R5754 VDD.n2259 VDD.t160 117.283
R5755 VDD.n2938 VDD.t65 117.283
R5756 VDD.n535 VDD.t47 116.742
R5757 VDD.n2692 VDD.t83 116.742
R5758 VDD.n111 VDD.n110 34.302
R5759 VDD.n617 VDD.n616 34.302
R5760 VDD.n1098 VDD.n1097 34.302
R5761 VDD.n2576 VDD.n2575 34.302
R5762 VDD.n765 VDD.n764 34.302
R5763 VDD.n2030 VDD.n2029 34.302
R5764 VDD.n3037 VDD.n3036 34.096
R5765 VDD.n1252 VDD.n1251 34.096
R5766 VDD.n2421 VDD.n2410 34.096
R5767 VDD.n944 VDD.n943 33.892
R5768 VDD.n476 VDD.n475 33.892
R5769 VDD.n259 VDD.n258 33.892
R5770 VDD.n2775 VDD.n2774 33.892
R5771 VDD.n2164 VDD.n2163 33.892
R5772 VDD.n1374 VDD.n1373 33.892
R5773 VDD.n1835 VDD.n1834 33.892
R5774 VDD.n109 VDD.n102 18.461
R5775 VDD.n618 VDD.n615 18.461
R5776 VDD.n1099 VDD.n1096 18.461
R5777 VDD.n2574 VDD.n2567 18.461
R5778 VDD.n2646 VDD.n2640 18.461
R5779 VDD.n2031 VDD.n2028 18.461
R5780 VDD.n763 VDD.n756 18.461
R5781 VDD.n1250 VDD.n1243 18.285
R5782 VDD.n3038 VDD.n3035 18.285
R5783 VDD.n2420 VDD.n2413 18.285
R5784 VDD.n942 VDD.n935 18.113
R5785 VDD.n474 VDD.n467 18.113
R5786 VDD.n260 VDD.n257 18.113
R5787 VDD.n2776 VDD.n2773 18.113
R5788 VDD.n2793 VDD.n2792 18.113
R5789 VDD.n1836 VDD.n1833 18.113
R5790 VDD.n1375 VDD.n1372 18.113
R5791 VDD.n2162 VDD.n2155 18.113
R5792 VDD.n120 VDD.n114 16.153
R5793 VDD.n604 VDD.n603 16.153
R5794 VDD.n1085 VDD.n1084 16.153
R5795 VDD.n2017 VDD.n2016 16.153
R5796 VDD.n1713 VDD.n1707 16.153
R5797 VDD.n41 VDD.n40 16.053
R5798 VDD.n634 VDD.n633 16.053
R5799 VDD.n1115 VDD.n1114 16.053
R5800 VDD.n2047 VDD.n2046 16.053
R5801 VDD.n774 VDD.n773 16.053
R5802 VDD.n1505 VDD.n1499 16
R5803 VDD.n3050 VDD.n3049 16
R5804 VDD.n2399 VDD.n2393 16
R5805 VDD.n1261 VDD.n1260 15.913
R5806 VDD.n3018 VDD.n3017 15.913
R5807 VDD.n2409 VDD.n2402 15.913
R5808 VDD.n953 VDD.n947 15.849
R5809 VDD.n485 VDD.n479 15.849
R5810 VDD.n246 VDD.n245 15.849
R5811 VDD.n1848 VDD.n1847 15.849
R5812 VDD.n1361 VDD.n1360 15.849
R5813 VDD.n2236 VDD.n2230 15.849
R5814 VDD.n874 VDD.n873 15.776
R5815 VDD.n406 VDD.n405 15.776
R5816 VDD.n276 VDD.n275 15.776
R5817 VDD.n1816 VDD.n1815 15.776
R5818 VDD.n1391 VDD.n1390 15.776
R5819 VDD.n2173 VDD.n2172 15.776
R5820 VDD.n67 VDD.n66 15
R5821 VDD.n705 VDD.n704 15
R5822 VDD.n1186 VDD.n1185 15
R5823 VDD.n2117 VDD.n2116 15
R5824 VDD.n800 VDD.n799 15
R5825 VDD.n1287 VDD.n1286 14.857
R5826 VDD.n2945 VDD.n2944 14.857
R5827 VDD.n2345 VDD.n2344 14.857
R5828 VDD.n900 VDD.n899 14.716
R5829 VDD.n432 VDD.n431 14.716
R5830 VDD.n347 VDD.n346 14.716
R5831 VDD.n2698 VDD.n2697 14.716
R5832 VDD.n1743 VDD.n1742 14.716
R5833 VDD.n1461 VDD.n1460 14.716
R5834 VDD.n2199 VDD.n2198 14.716
R5835 VDD.n99 VDD.n98 14.2
R5836 VDD.n646 VDD.n645 14.2
R5837 VDD.n1127 VDD.n1126 14.2
R5838 VDD.n2564 VDD.n2557 14.2
R5839 VDD.n2585 VDD.n2584 14.2
R5840 VDD.n2059 VDD.n2058 14.2
R5841 VDD.n1704 VDD.n1703 14.2
R5842 VDD.n1496 VDD.n1495 14.076
R5843 VDD.n3006 VDD.n3005 14.076
R5844 VDD.n2430 VDD.n2429 14.076
R5845 VDD.n932 VDD.n931 13.953
R5846 VDD.n464 VDD.n463 13.953
R5847 VDD.n288 VDD.n287 13.953
R5848 VDD.n2761 VDD.n2760 13.953
R5849 VDD.n2804 VDD.n2803 13.953
R5850 VDD.n1804 VDD.n1803 13.953
R5851 VDD.n1403 VDD.n1402 13.953
R5852 VDD.n2227 VDD.n2226 13.953
R5853 VDD.n32 VDD.n26 13.846
R5854 VDD.n592 VDD.n591 13.846
R5855 VDD.n1073 VDD.n1072 13.846
R5856 VDD.n2554 VDD.n2548 13.846
R5857 VDD.n2594 VDD.n2588 13.846
R5858 VDD.n2005 VDD.n2004 13.846
R5859 VDD.n753 VDD.n747 13.846
R5860 VDD.n1240 VDD.n1234 13.714
R5861 VDD.n3062 VDD.n3061 13.714
R5862 VDD.n2439 VDD.n2433 13.714
R5863 VDD.n865 VDD.n859 13.584
R5864 VDD.n397 VDD.n391 13.584
R5865 VDD.n234 VDD.n233 13.584
R5866 VDD.n2750 VDD.n2748 13.584
R5867 VDD.n2818 VDD.n2816 13.584
R5868 VDD.n1860 VDD.n1859 13.584
R5869 VDD.n1349 VDD.n1348 13.584
R5870 VDD.n2152 VDD.n2146 13.584
R5871 VDD.n80 VDD.n79 12.692
R5872 VDD.n693 VDD.n692 12.692
R5873 VDD.n1174 VDD.n1173 12.692
R5874 VDD.n2519 VDD.n2518 12.692
R5875 VDD.n2622 VDD.n2621 12.692
R5876 VDD.n2106 VDD.n2105 12.692
R5877 VDD.n1685 VDD.n1684 12.692
R5878 VDD.n1477 VDD.n1476 12.571
R5879 VDD.n2957 VDD.n2956 12.571
R5880 VDD.n2467 VDD.n2466 12.571
R5881 VDD.n913 VDD.n912 12.452
R5882 VDD.n445 VDD.n444 12.452
R5883 VDD.n335 VDD.n334 12.452
R5884 VDD.n2710 VDD.n2709 12.452
R5885 VDD.n2853 VDD.n2852 12.452
R5886 VDD.n1755 VDD.n1754 12.452
R5887 VDD.n1450 VDD.n1449 12.452
R5888 VDD.n2208 VDD.n2207 12.452
R5889 VDD.n50 VDD.n49 12.307
R5890 VDD.n658 VDD.n657 12.307
R5891 VDD.n1139 VDD.n1138 12.307
R5892 VDD.n2071 VDD.n2070 12.307
R5893 VDD.n783 VDD.n782 12.307
R5894 VDD.n1270 VDD.n1269 12.197
R5895 VDD.n2994 VDD.n2993 12.197
R5896 VDD.n2390 VDD.n2383 12.197
R5897 VDD.n883 VDD.n882 12.089
R5898 VDD.n415 VDD.n414 12.089
R5899 VDD.n300 VDD.n299 12.089
R5900 VDD.n1792 VDD.n1791 12.089
R5901 VDD.n1415 VDD.n1414 12.089
R5902 VDD.n2182 VDD.n2181 12.089
R5903 VDD.n129 VDD.n123 11.538
R5904 VDD.n580 VDD.n579 11.538
R5905 VDD.n1061 VDD.n1060 11.538
R5906 VDD.n1993 VDD.n1992 11.538
R5907 VDD.n1722 VDD.n1716 11.538
R5908 VDD.n1514 VDD.n1508 11.428
R5909 VDD.n3074 VDD.n3073 11.428
R5910 VDD.n2380 VDD.n2374 11.428
R5911 VDD.n2124 VDD.n2123 11.327
R5912 VDD.n1677 VDD.n1676 11.327
R5913 VDD.n2942 VDD.n2940 11.321
R5914 VDD.n962 VDD.n956 11.32
R5915 VDD.n494 VDD.n488 11.32
R5916 VDD.n222 VDD.n221 11.32
R5917 VDD.n1872 VDD.n1871 11.32
R5918 VDD.n1337 VDD.n1336 11.32
R5919 VDD.n2245 VDD.n2239 11.32
R5920 VDD.n1740 VDD.n1738 11.316
R5921 VDD.n1530 VDD.n1529 11.312
R5922 VDD.n1468 VDD.n1467 11.307
R5923 VDD.n2261 VDD.n2260 11.307
R5924 VDD.n2695 VDD.n2693 11.307
R5925 VDD.n72 VDD.n71 10.49
R5926 VDD.n715 VDD.n714 10.49
R5927 VDD.n1196 VDD.n1195 10.49
R5928 VDD.n2343 VDD.n2342 10.475
R5929 VDD.n357 VDD.n356 10.461
R5930 VDD.n905 VDD.n904 10.461
R5931 VDD.n437 VDD.n436 10.461
R5932 VDD.n58 VDD.n57 10.384
R5933 VDD.n681 VDD.n680 10.384
R5934 VDD.n1162 VDD.n1161 10.384
R5935 VDD.n2094 VDD.n2093 10.384
R5936 VDD.n791 VDD.n790 10.384
R5937 VDD.n90 VDD.n89 10.371
R5938 VDD.n670 VDD.n669 10.371
R5939 VDD.n1151 VDD.n1150 10.371
R5940 VDD.n2545 VDD.n2538 10.371
R5941 VDD.n2604 VDD.n2603 10.371
R5942 VDD.n2083 VDD.n2082 10.371
R5943 VDD.n1695 VDD.n1694 10.371
R5944 VDD.n1278 VDD.n1277 10.285
R5945 VDD.n2969 VDD.n2968 10.285
R5946 VDD.n2364 VDD.n2363 10.285
R5947 VDD.n1487 VDD.n1486 10.277
R5948 VDD.n2982 VDD.n2981 10.277
R5949 VDD.n2449 VDD.n2448 10.277
R5950 VDD.n891 VDD.n890 10.188
R5951 VDD.n423 VDD.n422 10.188
R5952 VDD.n323 VDD.n322 10.188
R5953 VDD.n1767 VDD.n1766 10.188
R5954 VDD.n1438 VDD.n1437 10.188
R5955 VDD.n2190 VDD.n2189 10.188
R5956 VDD.n923 VDD.n922 10.185
R5957 VDD.n455 VDD.n454 10.185
R5958 VDD.n312 VDD.n311 10.185
R5959 VDD.n2736 VDD.n2735 10.185
R5960 VDD.n2829 VDD.n2828 10.185
R5961 VDD.n1780 VDD.n1779 10.185
R5962 VDD.n1427 VDD.n1426 10.185
R5963 VDD.n2218 VDD.n2217 10.185
R5964 VDD.n1598 VDD.t112 9.544
R5965 VDD.n2883 VDD.t36 9.541
R5966 VDD.n821 VDD.t8 9.537
R5967 VDD.n0 VDD.t168 9.536
R5968 VDD.n825 VDD.t42 9.536
R5969 VDD.n2887 VDD.t40 9.536
R5970 VDD.n1602 VDD.t195 9.533
R5971 VDD.n3137 VDD.t214 9.533
R5972 VDD.n2310 VDD.t237 9.532
R5973 VDD.n1924 VDD.t70 9.532
R5974 VDD.n1608 VDD.t64 9.532
R5975 VDD.n2498 VDD.t50 9.532
R5976 VDD.n2503 VDD.t82 9.53
R5977 VDD.n833 VDD.t60 9.53
R5978 VDD.n1209 VDD.t2 9.53
R5979 VDD.n365 VDD.t149 9.53
R5980 VDD.n2491 VDD.t74 9.51
R5981 VDD.n725 VDD.t46 9.51
R5982 VDD.n1613 VDD.t6 9.51
R5983 VDD.n1584 VDD.t229 9.51
R5984 VDD.n1939 VDD.t22 9.51
R5985 VDD.n2329 VDD.t89 9.507
R5986 VDD.n1625 VDD.t159 9.507
R5987 VDD.n2333 VDD.t101 9.507
R5988 VDD.n818 VDD.t48 9.407
R5989 VDD.n2878 VDD.t84 9.407
R5990 VDD.n1918 VDD.t80 9.407
R5991 VDD.n1207 VDD.t153 9.407
R5992 VDD.n2307 VDD.t161 9.407
R5993 VDD.n1595 VDD.t170 9.404
R5994 VDD.n359 VDD.t30 9.404
R5995 VDD.n2890 VDD.t66 9.404
R5996 VDD.n2326 VDD.t26 9.396
R5997 VDD.n1203 VDD.t16 9.396
R5998 VDD.n2337 VDD.t130 9.396
R5999 VDD.n722 VDD.t209 9.393
R6000 VDD.n2488 VDD.t120 9.393
R6001 VDD.n1936 VDD.t134 9.393
R6002 VDD.n1622 VDD.t225 9.393
R6003 VDD.n1581 VDD.t179 9.393
R6004 VDD.n2325 VDD.t185 9.38
R6005 VDD.n721 VDD.t20 9.38
R6006 VDD.n1202 VDD.t182 9.38
R6007 VDD.n2487 VDD.t28 9.38
R6008 VDD.n1935 VDD.t132 9.38
R6009 VDD.n1621 VDD.t140 9.38
R6010 VDD.n1580 VDD.t227 9.38
R6011 VDD.n2336 VDD.t52 9.38
R6012 VDD.n2332 VDD.t24 9.363
R6013 VDD.n370 VDD.t187 9.363
R6014 VDD.n838 VDD.t62 9.363
R6015 VDD.n2331 VDD.t193 9.363
R6016 VDD.n1211 VDD.t189 9.361
R6017 VDD.n837 VDD.t233 9.361
R6018 VDD.n369 VDD.t91 9.361
R6019 VDD.n2324 VDD.t103 9.361
R6020 VDD.n2323 VDD.t87 9.361
R6021 VDD.n2322 VDD.t44 9.361
R6022 VDD.n1201 VDD.t95 9.361
R6023 VDD.n1200 VDD.t14 9.361
R6024 VDD.n1199 VDD.t76 9.361
R6025 VDD.n2493 VDD.t172 9.361
R6026 VDD.n3121 VDD.t105 9.361
R6027 VDD.n3123 VDD.t175 9.361
R6028 VDD.n3122 VDD.t124 9.361
R6029 VDD.n2327 VDD.t54 9.358
R6030 VDD.n2328 VDD.t155 9.358
R6031 VDD.n720 VDD.t200 9.358
R6032 VDD.n719 VDD.t206 9.358
R6033 VDD.n718 VDD.t97 9.358
R6034 VDD.n1204 VDD.t114 9.358
R6035 VDD.n1205 VDD.t157 9.358
R6036 VDD.n2486 VDD.t151 9.358
R6037 VDD.n2485 VDD.t122 9.358
R6038 VDD.n2484 VDD.t239 9.358
R6039 VDD.n370 VDD.t138 9.358
R6040 VDD.n838 VDD.t32 9.358
R6041 VDD.n1943 VDD.t78 9.358
R6042 VDD.n1941 VDD.t4 9.358
R6043 VDD.n1942 VDD.t142 9.358
R6044 VDD.n1629 VDD.t221 9.358
R6045 VDD.n1623 VDD.t191 9.358
R6046 VDD.n1624 VDD.t164 9.358
R6047 VDD.n1627 VDD.t107 9.358
R6048 VDD.n1628 VDD.t34 9.358
R6049 VDD.n1577 VDD.t147 9.358
R6050 VDD.n1582 VDD.t68 9.358
R6051 VDD.n1583 VDD.t204 9.358
R6052 VDD.n1579 VDD.t219 9.358
R6053 VDD.n1578 VDD.t177 9.358
R6054 VDD.n2338 VDD.t116 9.358
R6055 VDD.n2339 VDD.t110 9.358
R6056 VDD.n2332 VDD.t197 9.355
R6057 VDD.n1211 VDD.t57 9.355
R6058 VDD.n837 VDD.t18 9.355
R6059 VDD.n369 VDD.t211 9.355
R6060 VDD.n723 VDD.t235 9.355
R6061 VDD.n724 VDD.t166 9.355
R6062 VDD.n2489 VDD.t231 9.355
R6063 VDD.n2490 VDD.t72 9.355
R6064 VDD.n2493 VDD.t10 9.355
R6065 VDD.n2331 VDD.t127 9.355
R6066 VDD.n1937 VDD.t38 9.355
R6067 VDD.n1938 VDD.t93 9.355
R6068 VDD.n181 VDD.n179 9.312
R6069 VDD.n2937 VDD.n2936 9.312
R6070 VDD.n1015 VDD.n1014 9.303
R6071 VDD.n534 VDD.n533 9.303
R6072 VDD.n713 VDD.n712 9.3
R6073 VDD.n701 VDD.n700 9.3
R6074 VDD.n689 VDD.n688 9.3
R6075 VDD.n677 VDD.n676 9.3
R6076 VDD.n665 VDD.n664 9.3
R6077 VDD.n653 VDD.n652 9.3
R6078 VDD.n641 VDD.n640 9.3
R6079 VDD.n629 VDD.n628 9.3
R6080 VDD.n622 VDD.n621 9.3
R6081 VDD.n608 VDD.n607 9.3
R6082 VDD.n596 VDD.n595 9.3
R6083 VDD.n584 VDD.n583 9.3
R6084 VDD.n572 VDD.n571 9.3
R6085 VDD.n560 VDD.n559 9.3
R6086 VDD.n548 VDD.n547 9.3
R6087 VDD.n624 VDD.n623 9.3
R6088 VDD.n610 VDD.n609 9.3
R6089 VDD.n598 VDD.n597 9.3
R6090 VDD.n586 VDD.n585 9.3
R6091 VDD.n574 VDD.n573 9.3
R6092 VDD.n562 VDD.n561 9.3
R6093 VDD.n550 VDD.n549 9.3
R6094 VDD.n627 VDD.n626 9.3
R6095 VDD.n639 VDD.n638 9.3
R6096 VDD.n651 VDD.n650 9.3
R6097 VDD.n663 VDD.n662 9.3
R6098 VDD.n675 VDD.n674 9.3
R6099 VDD.n687 VDD.n686 9.3
R6100 VDD.n699 VDD.n698 9.3
R6101 VDD.n711 VDD.n710 9.3
R6102 VDD.n1194 VDD.n1193 9.3
R6103 VDD.n1182 VDD.n1181 9.3
R6104 VDD.n1170 VDD.n1169 9.3
R6105 VDD.n1158 VDD.n1157 9.3
R6106 VDD.n1146 VDD.n1145 9.3
R6107 VDD.n1134 VDD.n1133 9.3
R6108 VDD.n1122 VDD.n1121 9.3
R6109 VDD.n1110 VDD.n1109 9.3
R6110 VDD.n1103 VDD.n1102 9.3
R6111 VDD.n1089 VDD.n1088 9.3
R6112 VDD.n1077 VDD.n1076 9.3
R6113 VDD.n1065 VDD.n1064 9.3
R6114 VDD.n1053 VDD.n1052 9.3
R6115 VDD.n1041 VDD.n1040 9.3
R6116 VDD.n1029 VDD.n1028 9.3
R6117 VDD.n1105 VDD.n1104 9.3
R6118 VDD.n1091 VDD.n1090 9.3
R6119 VDD.n1079 VDD.n1078 9.3
R6120 VDD.n1067 VDD.n1066 9.3
R6121 VDD.n1055 VDD.n1054 9.3
R6122 VDD.n1043 VDD.n1042 9.3
R6123 VDD.n1031 VDD.n1030 9.3
R6124 VDD.n1108 VDD.n1107 9.3
R6125 VDD.n1120 VDD.n1119 9.3
R6126 VDD.n1132 VDD.n1131 9.3
R6127 VDD.n1144 VDD.n1143 9.3
R6128 VDD.n1156 VDD.n1155 9.3
R6129 VDD.n1168 VDD.n1167 9.3
R6130 VDD.n1180 VDD.n1179 9.3
R6131 VDD.n1192 VDD.n1191 9.3
R6132 VDD.n355 VDD.n354 9.3
R6133 VDD.n343 VDD.n342 9.3
R6134 VDD.n331 VDD.n330 9.3
R6135 VDD.n319 VDD.n318 9.3
R6136 VDD.n307 VDD.n306 9.3
R6137 VDD.n295 VDD.n294 9.3
R6138 VDD.n283 VDD.n282 9.3
R6139 VDD.n271 VDD.n270 9.3
R6140 VDD.n264 VDD.n263 9.3
R6141 VDD.n250 VDD.n249 9.3
R6142 VDD.n238 VDD.n237 9.3
R6143 VDD.n226 VDD.n225 9.3
R6144 VDD.n214 VDD.n213 9.3
R6145 VDD.n202 VDD.n201 9.3
R6146 VDD.n190 VDD.n189 9.3
R6147 VDD.n266 VDD.n265 9.3
R6148 VDD.n252 VDD.n251 9.3
R6149 VDD.n240 VDD.n239 9.3
R6150 VDD.n228 VDD.n227 9.3
R6151 VDD.n216 VDD.n215 9.3
R6152 VDD.n204 VDD.n203 9.3
R6153 VDD.n192 VDD.n191 9.3
R6154 VDD.n269 VDD.n268 9.3
R6155 VDD.n281 VDD.n280 9.3
R6156 VDD.n293 VDD.n292 9.3
R6157 VDD.n305 VDD.n304 9.3
R6158 VDD.n317 VDD.n316 9.3
R6159 VDD.n329 VDD.n328 9.3
R6160 VDD.n341 VDD.n340 9.3
R6161 VDD.n353 VDD.n352 9.3
R6162 VDD.n2525 VDD.n2524 9.3
R6163 VDD.n2535 VDD.n2534 9.3
R6164 VDD.n2544 VDD.n2543 9.3
R6165 VDD.n2554 VDD.n2553 9.3
R6166 VDD.n2563 VDD.n2562 9.3
R6167 VDD.n2574 VDD.n2573 9.3
R6168 VDD.n2646 VDD.n2645 9.3
R6169 VDD.n2691 VDD.n2646 9.3
R6170 VDD.n2582 VDD.n2581 9.3
R6171 VDD.n2594 VDD.n2593 9.3
R6172 VDD.n2601 VDD.n2600 9.3
R6173 VDD.n2613 VDD.n2612 9.3
R6174 VDD.n2620 VDD.n2619 9.3
R6175 VDD.n2632 VDD.n2631 9.3
R6176 VDD.n2516 VDD.n2515 9.3
R6177 VDD.n358 VDD.n357 9.3
R6178 VDD.n188 VDD.n187 9.3
R6179 VDD.n187 VDD.n186 9.3
R6180 VDD.n200 VDD.n199 9.3
R6181 VDD.n199 VDD.n198 9.3
R6182 VDD.n212 VDD.n211 9.3
R6183 VDD.n211 VDD.n210 9.3
R6184 VDD.n224 VDD.n223 9.3
R6185 VDD.n223 VDD.n222 9.3
R6186 VDD.n236 VDD.n235 9.3
R6187 VDD.n235 VDD.n234 9.3
R6188 VDD.n248 VDD.n247 9.3
R6189 VDD.n247 VDD.n246 9.3
R6190 VDD.n262 VDD.n261 9.3
R6191 VDD.n261 VDD.n260 9.3
R6192 VDD.n279 VDD.n278 9.3
R6193 VDD.n278 VDD.n277 9.3
R6194 VDD.n291 VDD.n290 9.3
R6195 VDD.n290 VDD.n289 9.3
R6196 VDD.n303 VDD.n302 9.3
R6197 VDD.n302 VDD.n301 9.3
R6198 VDD.n315 VDD.n314 9.3
R6199 VDD.n314 VDD.n313 9.3
R6200 VDD.n327 VDD.n326 9.3
R6201 VDD.n326 VDD.n325 9.3
R6202 VDD.n339 VDD.n338 9.3
R6203 VDD.n338 VDD.n337 9.3
R6204 VDD.n351 VDD.n350 9.3
R6205 VDD.n350 VDD.n349 9.3
R6206 VDD.n379 VDD.n378 9.3
R6207 VDD.n535 VDD.n379 9.3
R6208 VDD.n503 VDD.n502 9.3
R6209 VDD.n535 VDD.n503 9.3
R6210 VDD.n388 VDD.n387 9.3
R6211 VDD.n535 VDD.n388 9.3
R6212 VDD.n494 VDD.n493 9.3
R6213 VDD.n535 VDD.n494 9.3
R6214 VDD.n397 VDD.n396 9.3
R6215 VDD.n535 VDD.n397 9.3
R6216 VDD.n485 VDD.n484 9.3
R6217 VDD.n535 VDD.n485 9.3
R6218 VDD.n474 VDD.n473 9.3
R6219 VDD.n403 VDD.n402 9.3
R6220 VDD.n461 VDD.n460 9.3
R6221 VDD.n412 VDD.n411 9.3
R6222 VDD.n452 VDD.n451 9.3
R6223 VDD.n421 VDD.n420 9.3
R6224 VDD.n443 VDD.n442 9.3
R6225 VDD.n430 VDD.n429 9.3
R6226 VDD.n847 VDD.n846 9.3
R6227 VDD.n1016 VDD.n847 9.3
R6228 VDD.n971 VDD.n970 9.3
R6229 VDD.n1016 VDD.n971 9.3
R6230 VDD.n856 VDD.n855 9.3
R6231 VDD.n1016 VDD.n856 9.3
R6232 VDD.n962 VDD.n961 9.3
R6233 VDD.n1016 VDD.n962 9.3
R6234 VDD.n865 VDD.n864 9.3
R6235 VDD.n1016 VDD.n865 9.3
R6236 VDD.n953 VDD.n952 9.3
R6237 VDD.n1016 VDD.n953 9.3
R6238 VDD.n942 VDD.n941 9.3
R6239 VDD.n871 VDD.n870 9.3
R6240 VDD.n929 VDD.n928 9.3
R6241 VDD.n880 VDD.n879 9.3
R6242 VDD.n920 VDD.n919 9.3
R6243 VDD.n889 VDD.n888 9.3
R6244 VDD.n911 VDD.n910 9.3
R6245 VDD.n898 VDD.n897 9.3
R6246 VDD.n1197 VDD.n1196 9.3
R6247 VDD.n1027 VDD.n1026 9.3
R6248 VDD.n1026 VDD.n1025 9.3
R6249 VDD.n1039 VDD.n1038 9.3
R6250 VDD.n1038 VDD.n1037 9.3
R6251 VDD.n1051 VDD.n1050 9.3
R6252 VDD.n1050 VDD.n1049 9.3
R6253 VDD.n1063 VDD.n1062 9.3
R6254 VDD.n1062 VDD.n1061 9.3
R6255 VDD.n1075 VDD.n1074 9.3
R6256 VDD.n1074 VDD.n1073 9.3
R6257 VDD.n1087 VDD.n1086 9.3
R6258 VDD.n1086 VDD.n1085 9.3
R6259 VDD.n1101 VDD.n1100 9.3
R6260 VDD.n1100 VDD.n1099 9.3
R6261 VDD.n1118 VDD.n1117 9.3
R6262 VDD.n1117 VDD.n1116 9.3
R6263 VDD.n1130 VDD.n1129 9.3
R6264 VDD.n1129 VDD.n1128 9.3
R6265 VDD.n1142 VDD.n1141 9.3
R6266 VDD.n1141 VDD.n1140 9.3
R6267 VDD.n1154 VDD.n1153 9.3
R6268 VDD.n1153 VDD.n1152 9.3
R6269 VDD.n1166 VDD.n1165 9.3
R6270 VDD.n1165 VDD.n1164 9.3
R6271 VDD.n1178 VDD.n1177 9.3
R6272 VDD.n1177 VDD.n1176 9.3
R6273 VDD.n1190 VDD.n1189 9.3
R6274 VDD.n1189 VDD.n1188 9.3
R6275 VDD.n716 VDD.n715 9.3
R6276 VDD.n546 VDD.n545 9.3
R6277 VDD.n545 VDD.n544 9.3
R6278 VDD.n558 VDD.n557 9.3
R6279 VDD.n557 VDD.n556 9.3
R6280 VDD.n570 VDD.n569 9.3
R6281 VDD.n569 VDD.n568 9.3
R6282 VDD.n582 VDD.n581 9.3
R6283 VDD.n581 VDD.n580 9.3
R6284 VDD.n594 VDD.n593 9.3
R6285 VDD.n593 VDD.n592 9.3
R6286 VDD.n606 VDD.n605 9.3
R6287 VDD.n605 VDD.n604 9.3
R6288 VDD.n620 VDD.n619 9.3
R6289 VDD.n619 VDD.n618 9.3
R6290 VDD.n637 VDD.n636 9.3
R6291 VDD.n636 VDD.n635 9.3
R6292 VDD.n649 VDD.n648 9.3
R6293 VDD.n648 VDD.n647 9.3
R6294 VDD.n661 VDD.n660 9.3
R6295 VDD.n660 VDD.n659 9.3
R6296 VDD.n673 VDD.n672 9.3
R6297 VDD.n672 VDD.n671 9.3
R6298 VDD.n685 VDD.n684 9.3
R6299 VDD.n684 VDD.n683 9.3
R6300 VDD.n697 VDD.n696 9.3
R6301 VDD.n696 VDD.n695 9.3
R6302 VDD.n709 VDD.n708 9.3
R6303 VDD.n708 VDD.n707 9.3
R6304 VDD.n14 VDD.n13 9.3
R6305 VDD.n177 VDD.n14 9.3
R6306 VDD.n138 VDD.n137 9.3
R6307 VDD.n177 VDD.n138 9.3
R6308 VDD.n23 VDD.n22 9.3
R6309 VDD.n177 VDD.n23 9.3
R6310 VDD.n129 VDD.n128 9.3
R6311 VDD.n177 VDD.n129 9.3
R6312 VDD.n32 VDD.n31 9.3
R6313 VDD.n177 VDD.n32 9.3
R6314 VDD.n120 VDD.n119 9.3
R6315 VDD.n177 VDD.n120 9.3
R6316 VDD.n109 VDD.n108 9.3
R6317 VDD.n38 VDD.n37 9.3
R6318 VDD.n96 VDD.n95 9.3
R6319 VDD.n47 VDD.n46 9.3
R6320 VDD.n87 VDD.n86 9.3
R6321 VDD.n56 VDD.n55 9.3
R6322 VDD.n78 VDD.n77 9.3
R6323 VDD.n65 VDD.n64 9.3
R6324 VDD.n2874 VDD.n2873 9.3
R6325 VDD.n2861 VDD.n2860 9.3
R6326 VDD.n2849 VDD.n2848 9.3
R6327 VDD.n2836 VDD.n2835 9.3
R6328 VDD.n2824 VDD.n2823 9.3
R6329 VDD.n2811 VDD.n2810 9.3
R6330 VDD.n2799 VDD.n2798 9.3
R6331 VDD.n2787 VDD.n2786 9.3
R6332 VDD.n2780 VDD.n2779 9.3
R6333 VDD.n2766 VDD.n2765 9.3
R6334 VDD.n2754 VDD.n2753 9.3
R6335 VDD.n2741 VDD.n2740 9.3
R6336 VDD.n2729 VDD.n2728 9.3
R6337 VDD.n2716 VDD.n2715 9.3
R6338 VDD.n2704 VDD.n2703 9.3
R6339 VDD.n2877 VDD.n2876 9.3
R6340 VDD.n2782 VDD.n2781 9.3
R6341 VDD.n2768 VDD.n2767 9.3
R6342 VDD.n2756 VDD.n2755 9.3
R6343 VDD.n2743 VDD.n2742 9.3
R6344 VDD.n2731 VDD.n2730 9.3
R6345 VDD.n2718 VDD.n2717 9.3
R6346 VDD.n2706 VDD.n2705 9.3
R6347 VDD.n2702 VDD.n2701 9.3
R6348 VDD.n2701 VDD.n2700 9.3
R6349 VDD.n2714 VDD.n2713 9.3
R6350 VDD.n2713 VDD.n2712 9.3
R6351 VDD.n2727 VDD.n2726 9.3
R6352 VDD.n2726 VDD.n2725 9.3
R6353 VDD.n2739 VDD.n2738 9.3
R6354 VDD.n2738 VDD.n2737 9.3
R6355 VDD.n2752 VDD.n2751 9.3
R6356 VDD.n2751 VDD.n2750 9.3
R6357 VDD.n2764 VDD.n2763 9.3
R6358 VDD.n2763 VDD.n2762 9.3
R6359 VDD.n2778 VDD.n2777 9.3
R6360 VDD.n2777 VDD.n2776 9.3
R6361 VDD.n2785 VDD.n2784 9.3
R6362 VDD.n2795 VDD.n2794 9.3
R6363 VDD.n2794 VDD.n2793 9.3
R6364 VDD.n2797 VDD.n2796 9.3
R6365 VDD.n2807 VDD.n2806 9.3
R6366 VDD.n2806 VDD.n2805 9.3
R6367 VDD.n2809 VDD.n2808 9.3
R6368 VDD.n2820 VDD.n2819 9.3
R6369 VDD.n2819 VDD.n2818 9.3
R6370 VDD.n2822 VDD.n2821 9.3
R6371 VDD.n2832 VDD.n2831 9.3
R6372 VDD.n2831 VDD.n2830 9.3
R6373 VDD.n2834 VDD.n2833 9.3
R6374 VDD.n2845 VDD.n2844 9.3
R6375 VDD.n2844 VDD.n2843 9.3
R6376 VDD.n2847 VDD.n2846 9.3
R6377 VDD.n2857 VDD.n2856 9.3
R6378 VDD.n2856 VDD.n2855 9.3
R6379 VDD.n2859 VDD.n2858 9.3
R6380 VDD.n2870 VDD.n2869 9.3
R6381 VDD.n2869 VDD.n2868 9.3
R6382 VDD.n2872 VDD.n2871 9.3
R6383 VDD.n1914 VDD.n1913 9.3
R6384 VDD.n1902 VDD.n1901 9.3
R6385 VDD.n1890 VDD.n1889 9.3
R6386 VDD.n1878 VDD.n1877 9.3
R6387 VDD.n1866 VDD.n1865 9.3
R6388 VDD.n1854 VDD.n1853 9.3
R6389 VDD.n1842 VDD.n1841 9.3
R6390 VDD.n1828 VDD.n1827 9.3
R6391 VDD.n1821 VDD.n1820 9.3
R6392 VDD.n1809 VDD.n1808 9.3
R6393 VDD.n1797 VDD.n1796 9.3
R6394 VDD.n1785 VDD.n1784 9.3
R6395 VDD.n1773 VDD.n1772 9.3
R6396 VDD.n1761 VDD.n1760 9.3
R6397 VDD.n1749 VDD.n1748 9.3
R6398 VDD.n1912 VDD.n1911 9.3
R6399 VDD.n1900 VDD.n1899 9.3
R6400 VDD.n1888 VDD.n1887 9.3
R6401 VDD.n1876 VDD.n1875 9.3
R6402 VDD.n1864 VDD.n1863 9.3
R6403 VDD.n1852 VDD.n1851 9.3
R6404 VDD.n1840 VDD.n1839 9.3
R6405 VDD.n1826 VDD.n1825 9.3
R6406 VDD.n1823 VDD.n1822 9.3
R6407 VDD.n1811 VDD.n1810 9.3
R6408 VDD.n1799 VDD.n1798 9.3
R6409 VDD.n1787 VDD.n1786 9.3
R6410 VDD.n1775 VDD.n1774 9.3
R6411 VDD.n1763 VDD.n1762 9.3
R6412 VDD.n1751 VDD.n1750 9.3
R6413 VDD.n1293 VDD.n1292 9.3
R6414 VDD.n1305 VDD.n1304 9.3
R6415 VDD.n1317 VDD.n1316 9.3
R6416 VDD.n1329 VDD.n1328 9.3
R6417 VDD.n1341 VDD.n1340 9.3
R6418 VDD.n1353 VDD.n1352 9.3
R6419 VDD.n1365 VDD.n1364 9.3
R6420 VDD.n1379 VDD.n1378 9.3
R6421 VDD.n1386 VDD.n1385 9.3
R6422 VDD.n1398 VDD.n1397 9.3
R6423 VDD.n1410 VDD.n1409 9.3
R6424 VDD.n1422 VDD.n1421 9.3
R6425 VDD.n1434 VDD.n1433 9.3
R6426 VDD.n1446 VDD.n1445 9.3
R6427 VDD.n1458 VDD.n1457 9.3
R6428 VDD.n1295 VDD.n1294 9.3
R6429 VDD.n1307 VDD.n1306 9.3
R6430 VDD.n1319 VDD.n1318 9.3
R6431 VDD.n1331 VDD.n1330 9.3
R6432 VDD.n1343 VDD.n1342 9.3
R6433 VDD.n1355 VDD.n1354 9.3
R6434 VDD.n1367 VDD.n1366 9.3
R6435 VDD.n1382 VDD.n1381 9.3
R6436 VDD.n1384 VDD.n1383 9.3
R6437 VDD.n1396 VDD.n1395 9.3
R6438 VDD.n1408 VDD.n1407 9.3
R6439 VDD.n1420 VDD.n1419 9.3
R6440 VDD.n1432 VDD.n1431 9.3
R6441 VDD.n1444 VDD.n1443 9.3
R6442 VDD.n1456 VDD.n1455 9.3
R6443 VDD.n1949 VDD.n1948 9.3
R6444 VDD.n1961 VDD.n1960 9.3
R6445 VDD.n1973 VDD.n1972 9.3
R6446 VDD.n1985 VDD.n1984 9.3
R6447 VDD.n1997 VDD.n1996 9.3
R6448 VDD.n2009 VDD.n2008 9.3
R6449 VDD.n2021 VDD.n2020 9.3
R6450 VDD.n2035 VDD.n2034 9.3
R6451 VDD.n2042 VDD.n2041 9.3
R6452 VDD.n2054 VDD.n2053 9.3
R6453 VDD.n2066 VDD.n2065 9.3
R6454 VDD.n2078 VDD.n2077 9.3
R6455 VDD.n2090 VDD.n2089 9.3
R6456 VDD.n2102 VDD.n2101 9.3
R6457 VDD.n2114 VDD.n2113 9.3
R6458 VDD.n1951 VDD.n1950 9.3
R6459 VDD.n1963 VDD.n1962 9.3
R6460 VDD.n1975 VDD.n1974 9.3
R6461 VDD.n1987 VDD.n1986 9.3
R6462 VDD.n1999 VDD.n1998 9.3
R6463 VDD.n2011 VDD.n2010 9.3
R6464 VDD.n2023 VDD.n2022 9.3
R6465 VDD.n2038 VDD.n2037 9.3
R6466 VDD.n2040 VDD.n2039 9.3
R6467 VDD.n2052 VDD.n2051 9.3
R6468 VDD.n2064 VDD.n2063 9.3
R6469 VDD.n2076 VDD.n2075 9.3
R6470 VDD.n2088 VDD.n2087 9.3
R6471 VDD.n2100 VDD.n2099 9.3
R6472 VDD.n2112 VDD.n2111 9.3
R6473 VDD.n3116 VDD.n3115 9.3
R6474 VDD.n3104 VDD.n3103 9.3
R6475 VDD.n3092 VDD.n3091 9.3
R6476 VDD.n3080 VDD.n3079 9.3
R6477 VDD.n3068 VDD.n3067 9.3
R6478 VDD.n3056 VDD.n3055 9.3
R6479 VDD.n3044 VDD.n3043 9.3
R6480 VDD.n3030 VDD.n3029 9.3
R6481 VDD.n3023 VDD.n3022 9.3
R6482 VDD.n3011 VDD.n3010 9.3
R6483 VDD.n2999 VDD.n2998 9.3
R6484 VDD.n2987 VDD.n2986 9.3
R6485 VDD.n2975 VDD.n2974 9.3
R6486 VDD.n2963 VDD.n2962 9.3
R6487 VDD.n2951 VDD.n2950 9.3
R6488 VDD.n3114 VDD.n3113 9.3
R6489 VDD.n3102 VDD.n3101 9.3
R6490 VDD.n3090 VDD.n3089 9.3
R6491 VDD.n3078 VDD.n3077 9.3
R6492 VDD.n3066 VDD.n3065 9.3
R6493 VDD.n3054 VDD.n3053 9.3
R6494 VDD.n3042 VDD.n3041 9.3
R6495 VDD.n3028 VDD.n3027 9.3
R6496 VDD.n3025 VDD.n3024 9.3
R6497 VDD.n3013 VDD.n3012 9.3
R6498 VDD.n3001 VDD.n3000 9.3
R6499 VDD.n2989 VDD.n2988 9.3
R6500 VDD.n2977 VDD.n2976 9.3
R6501 VDD.n2965 VDD.n2964 9.3
R6502 VDD.n2953 VDD.n2952 9.3
R6503 VDD.n3112 VDD.n3111 9.3
R6504 VDD.n3111 VDD.n3110 9.3
R6505 VDD.n3100 VDD.n3099 9.3
R6506 VDD.n3099 VDD.n3098 9.3
R6507 VDD.n3088 VDD.n3087 9.3
R6508 VDD.n3087 VDD.n3086 9.3
R6509 VDD.n3076 VDD.n3075 9.3
R6510 VDD.n3075 VDD.n3074 9.3
R6511 VDD.n3064 VDD.n3063 9.3
R6512 VDD.n3063 VDD.n3062 9.3
R6513 VDD.n3052 VDD.n3051 9.3
R6514 VDD.n3051 VDD.n3050 9.3
R6515 VDD.n3040 VDD.n3039 9.3
R6516 VDD.n3039 VDD.n3038 9.3
R6517 VDD.n3021 VDD.n3020 9.3
R6518 VDD.n3020 VDD.n3019 9.3
R6519 VDD.n3009 VDD.n3008 9.3
R6520 VDD.n3008 VDD.n3007 9.3
R6521 VDD.n2997 VDD.n2996 9.3
R6522 VDD.n2996 VDD.n2995 9.3
R6523 VDD.n2985 VDD.n2984 9.3
R6524 VDD.n2984 VDD.n2983 9.3
R6525 VDD.n2973 VDD.n2972 9.3
R6526 VDD.n2972 VDD.n2971 9.3
R6527 VDD.n2961 VDD.n2960 9.3
R6528 VDD.n2960 VDD.n2959 9.3
R6529 VDD.n2949 VDD.n2948 9.3
R6530 VDD.n2948 VDD.n2947 9.3
R6531 VDD.n3119 VDD.n3118 9.3
R6532 VDD.n1222 VDD.n1221 9.3
R6533 VDD.n1528 VDD.n1222 9.3
R6534 VDD.n1523 VDD.n1522 9.3
R6535 VDD.n1528 VDD.n1523 9.3
R6536 VDD.n1231 VDD.n1230 9.3
R6537 VDD.n1528 VDD.n1231 9.3
R6538 VDD.n1514 VDD.n1513 9.3
R6539 VDD.n1528 VDD.n1514 9.3
R6540 VDD.n1240 VDD.n1239 9.3
R6541 VDD.n1528 VDD.n1240 9.3
R6542 VDD.n1505 VDD.n1504 9.3
R6543 VDD.n1528 VDD.n1505 9.3
R6544 VDD.n1250 VDD.n1249 9.3
R6545 VDD.n1258 VDD.n1257 9.3
R6546 VDD.n1493 VDD.n1492 9.3
R6547 VDD.n1267 VDD.n1266 9.3
R6548 VDD.n1484 VDD.n1483 9.3
R6549 VDD.n1276 VDD.n1275 9.3
R6550 VDD.n1475 VDD.n1474 9.3
R6551 VDD.n1285 VDD.n1284 9.3
R6552 VDD.n735 VDD.n734 9.3
R6553 VDD.n1736 VDD.n735 9.3
R6554 VDD.n1731 VDD.n1730 9.3
R6555 VDD.n1736 VDD.n1731 9.3
R6556 VDD.n744 VDD.n743 9.3
R6557 VDD.n1736 VDD.n744 9.3
R6558 VDD.n1722 VDD.n1721 9.3
R6559 VDD.n1736 VDD.n1722 9.3
R6560 VDD.n753 VDD.n752 9.3
R6561 VDD.n1736 VDD.n753 9.3
R6562 VDD.n1713 VDD.n1712 9.3
R6563 VDD.n1736 VDD.n1713 9.3
R6564 VDD.n763 VDD.n762 9.3
R6565 VDD.n771 VDD.n770 9.3
R6566 VDD.n1701 VDD.n1700 9.3
R6567 VDD.n780 VDD.n779 9.3
R6568 VDD.n1692 VDD.n1691 9.3
R6569 VDD.n789 VDD.n788 9.3
R6570 VDD.n1683 VDD.n1682 9.3
R6571 VDD.n798 VDD.n797 9.3
R6572 VDD.n1959 VDD.n1958 9.3
R6573 VDD.n1958 VDD.n1957 9.3
R6574 VDD.n1971 VDD.n1970 9.3
R6575 VDD.n1970 VDD.n1969 9.3
R6576 VDD.n1983 VDD.n1982 9.3
R6577 VDD.n1982 VDD.n1981 9.3
R6578 VDD.n1995 VDD.n1994 9.3
R6579 VDD.n1994 VDD.n1993 9.3
R6580 VDD.n2007 VDD.n2006 9.3
R6581 VDD.n2006 VDD.n2005 9.3
R6582 VDD.n2019 VDD.n2018 9.3
R6583 VDD.n2018 VDD.n2017 9.3
R6584 VDD.n2033 VDD.n2032 9.3
R6585 VDD.n2032 VDD.n2031 9.3
R6586 VDD.n2050 VDD.n2049 9.3
R6587 VDD.n2049 VDD.n2048 9.3
R6588 VDD.n2062 VDD.n2061 9.3
R6589 VDD.n2061 VDD.n2060 9.3
R6590 VDD.n2074 VDD.n2073 9.3
R6591 VDD.n2073 VDD.n2072 9.3
R6592 VDD.n2086 VDD.n2085 9.3
R6593 VDD.n2085 VDD.n2084 9.3
R6594 VDD.n2098 VDD.n2097 9.3
R6595 VDD.n2097 VDD.n2096 9.3
R6596 VDD.n2110 VDD.n2109 9.3
R6597 VDD.n2109 VDD.n2108 9.3
R6598 VDD.n2121 VDD.n2120 9.3
R6599 VDD.n2120 VDD.n2119 9.3
R6600 VDD.n1947 VDD.n1946 9.3
R6601 VDD.n2134 VDD.n2133 9.3
R6602 VDD.n2259 VDD.n2134 9.3
R6603 VDD.n2254 VDD.n2253 9.3
R6604 VDD.n2259 VDD.n2254 9.3
R6605 VDD.n2143 VDD.n2142 9.3
R6606 VDD.n2259 VDD.n2143 9.3
R6607 VDD.n2245 VDD.n2244 9.3
R6608 VDD.n2259 VDD.n2245 9.3
R6609 VDD.n2152 VDD.n2151 9.3
R6610 VDD.n2259 VDD.n2152 9.3
R6611 VDD.n2236 VDD.n2235 9.3
R6612 VDD.n2259 VDD.n2236 9.3
R6613 VDD.n2162 VDD.n2161 9.3
R6614 VDD.n2170 VDD.n2169 9.3
R6615 VDD.n2224 VDD.n2223 9.3
R6616 VDD.n2179 VDD.n2178 9.3
R6617 VDD.n2215 VDD.n2214 9.3
R6618 VDD.n2188 VDD.n2187 9.3
R6619 VDD.n2206 VDD.n2205 9.3
R6620 VDD.n2197 VDD.n2196 9.3
R6621 VDD.n1303 VDD.n1302 9.3
R6622 VDD.n1302 VDD.n1301 9.3
R6623 VDD.n1315 VDD.n1314 9.3
R6624 VDD.n1314 VDD.n1313 9.3
R6625 VDD.n1327 VDD.n1326 9.3
R6626 VDD.n1326 VDD.n1325 9.3
R6627 VDD.n1339 VDD.n1338 9.3
R6628 VDD.n1338 VDD.n1337 9.3
R6629 VDD.n1351 VDD.n1350 9.3
R6630 VDD.n1350 VDD.n1349 9.3
R6631 VDD.n1363 VDD.n1362 9.3
R6632 VDD.n1362 VDD.n1361 9.3
R6633 VDD.n1377 VDD.n1376 9.3
R6634 VDD.n1376 VDD.n1375 9.3
R6635 VDD.n1394 VDD.n1393 9.3
R6636 VDD.n1393 VDD.n1392 9.3
R6637 VDD.n1406 VDD.n1405 9.3
R6638 VDD.n1405 VDD.n1404 9.3
R6639 VDD.n1418 VDD.n1417 9.3
R6640 VDD.n1417 VDD.n1416 9.3
R6641 VDD.n1430 VDD.n1429 9.3
R6642 VDD.n1429 VDD.n1428 9.3
R6643 VDD.n1442 VDD.n1441 9.3
R6644 VDD.n1441 VDD.n1440 9.3
R6645 VDD.n1454 VDD.n1453 9.3
R6646 VDD.n1453 VDD.n1452 9.3
R6647 VDD.n1465 VDD.n1464 9.3
R6648 VDD.n1464 VDD.n1463 9.3
R6649 VDD.n1291 VDD.n1290 9.3
R6650 VDD.n1910 VDD.n1909 9.3
R6651 VDD.n1909 VDD.n1908 9.3
R6652 VDD.n1898 VDD.n1897 9.3
R6653 VDD.n1897 VDD.n1896 9.3
R6654 VDD.n1886 VDD.n1885 9.3
R6655 VDD.n1885 VDD.n1884 9.3
R6656 VDD.n1874 VDD.n1873 9.3
R6657 VDD.n1873 VDD.n1872 9.3
R6658 VDD.n1862 VDD.n1861 9.3
R6659 VDD.n1861 VDD.n1860 9.3
R6660 VDD.n1850 VDD.n1849 9.3
R6661 VDD.n1849 VDD.n1848 9.3
R6662 VDD.n1838 VDD.n1837 9.3
R6663 VDD.n1837 VDD.n1836 9.3
R6664 VDD.n1819 VDD.n1818 9.3
R6665 VDD.n1818 VDD.n1817 9.3
R6666 VDD.n1807 VDD.n1806 9.3
R6667 VDD.n1806 VDD.n1805 9.3
R6668 VDD.n1795 VDD.n1794 9.3
R6669 VDD.n1794 VDD.n1793 9.3
R6670 VDD.n1783 VDD.n1782 9.3
R6671 VDD.n1782 VDD.n1781 9.3
R6672 VDD.n1771 VDD.n1770 9.3
R6673 VDD.n1770 VDD.n1769 9.3
R6674 VDD.n1759 VDD.n1758 9.3
R6675 VDD.n1758 VDD.n1757 9.3
R6676 VDD.n1747 VDD.n1746 9.3
R6677 VDD.n1746 VDD.n1745 9.3
R6678 VDD.n1917 VDD.n1916 9.3
R6679 VDD.n2351 VDD.n2350 9.3
R6680 VDD.n2361 VDD.n2360 9.3
R6681 VDD.n2370 VDD.n2369 9.3
R6682 VDD.n2380 VDD.n2379 9.3
R6683 VDD.n2389 VDD.n2388 9.3
R6684 VDD.n2399 VDD.n2398 9.3
R6685 VDD.n2408 VDD.n2407 9.3
R6686 VDD.n2420 VDD.n2419 9.3
R6687 VDD.n2427 VDD.n2426 9.3
R6688 VDD.n2439 VDD.n2438 9.3
R6689 VDD.n2446 VDD.n2445 9.3
R6690 VDD.n2458 VDD.n2457 9.3
R6691 VDD.n2465 VDD.n2464 9.3
R6692 VDD.n2477 VDD.n2476 9.3
R6693 VDD.n2690 VDD.n2689 9.295
R6694 VDD.n176 VDD.n175 9.294
R6695 VDD.n539 VDD.n537 9.294
R6696 VDD.n1020 VDD.n1018 9.294
R6697 VDD.n23 VDD.n17 9.23
R6698 VDD.n568 VDD.n567 9.23
R6699 VDD.n1049 VDD.n1048 9.23
R6700 VDD.n2535 VDD.n2529 9.23
R6701 VDD.n2613 VDD.n2607 9.23
R6702 VDD.n1981 VDD.n1980 9.23
R6703 VDD.n744 VDD.n738 9.23
R6704 VDD.n1231 VDD.n1225 9.142
R6705 VDD.n3086 VDD.n3085 9.142
R6706 VDD.n2458 VDD.n2452 9.142
R6707 VDD.n856 VDD.n850 9.056
R6708 VDD.n388 VDD.n382 9.056
R6709 VDD.n210 VDD.n209 9.056
R6710 VDD.n2725 VDD.n2723 9.056
R6711 VDD.n2843 VDD.n2841 9.056
R6712 VDD.n1884 VDD.n1883 9.056
R6713 VDD.n1325 VDD.n1324 9.056
R6714 VDD.n2143 VDD.n2137 9.056
R6715 VDD.n535 VDD.n433 8.654
R6716 VDD.n1016 VDD.n901 8.654
R6717 VDD.n2259 VDD.n2200 8.654
R6718 VDD.n1528 VDD.n1288 8.652
R6719 VDD.n2938 VDD.n2352 8.652
R6720 VDD.n177 VDD.n68 8.65
R6721 VDD.n1736 VDD.n801 8.65
R6722 VDD.n535 VDD.n446 8.556
R6723 VDD.n1016 VDD.n914 8.556
R6724 VDD.n2259 VDD.n2209 8.556
R6725 VDD.n1528 VDD.n1478 8.554
R6726 VDD.n2938 VDD.n2468 8.554
R6727 VDD.n2691 VDD.n2526 8.551
R6728 VDD.n2691 VDD.n2623 8.551
R6729 VDD.n177 VDD.n81 8.551
R6730 VDD.n1736 VDD.n1686 8.551
R6731 VDD.n535 VDD.n424 8.461
R6732 VDD.n1016 VDD.n892 8.461
R6733 VDD.n2259 VDD.n2191 8.461
R6734 VDD.n1916 VDD.n1915 8.459
R6735 VDD.n1290 VDD.n1289 8.459
R6736 VDD.n2258 VDD.n2257 8.459
R6737 VDD.n3118 VDD.n3117 8.459
R6738 VDD.n1527 VDD.n1526 8.459
R6739 VDD.n1946 VDD.n1945 8.459
R6740 VDD.n1735 VDD.n1734 8.459
R6741 VDD.n2876 VDD.n2875 8.458
R6742 VDD.n2637 VDD.n2636 8.457
R6743 VDD.n1528 VDD.n1279 8.457
R6744 VDD.n2938 VDD.n2371 8.457
R6745 VDD.n177 VDD.n59 8.454
R6746 VDD.n1736 VDD.n792 8.454
R6747 VDD.n2938 VDD.n2937 8.453
R6748 VDD.n179 VDD.n178 8.453
R6749 VDD.n2691 VDD.n2637 8.453
R6750 VDD.n1018 VDD.n1017 8.453
R6751 VDD.n537 VDD.n536 8.453
R6752 VDD.n177 VDD.n176 8.453
R6753 VDD.n535 VDD.n534 8.453
R6754 VDD.n1016 VDD.n1015 8.453
R6755 VDD.n2691 VDD.n2690 8.451
R6756 VDD.n1736 VDD.n1735 8.451
R6757 VDD.n2259 VDD.n2258 8.451
R6758 VDD.n1528 VDD.n1527 8.451
R6759 VDD.n59 VDD.n58 8.39
R6760 VDD.n682 VDD.n681 8.39
R6761 VDD.n1163 VDD.n1162 8.39
R6762 VDD.n2095 VDD.n2094 8.39
R6763 VDD.n792 VDD.n791 8.39
R6764 VDD.n535 VDD.n455 8.368
R6765 VDD.n1016 VDD.n923 8.368
R6766 VDD.n2259 VDD.n2218 8.368
R6767 VDD.n1528 VDD.n1487 8.363
R6768 VDD.n2938 VDD.n2449 8.363
R6769 VDD.n2691 VDD.n2545 8.359
R6770 VDD.n2691 VDD.n2604 8.359
R6771 VDD.n177 VDD.n90 8.359
R6772 VDD.n1736 VDD.n1695 8.359
R6773 VDD.n1279 VDD.n1278 8.314
R6774 VDD.n2970 VDD.n2969 8.314
R6775 VDD.n2371 VDD.n2364 8.314
R6776 VDD.n535 VDD.n415 8.277
R6777 VDD.n1016 VDD.n883 8.277
R6778 VDD.n2259 VDD.n2182 8.277
R6779 VDD.n1528 VDD.n1270 8.272
R6780 VDD.n2938 VDD.n2390 8.272
R6781 VDD.n177 VDD.n50 8.266
R6782 VDD.n1736 VDD.n783 8.266
R6783 VDD.n892 VDD.n891 8.239
R6784 VDD.n424 VDD.n423 8.239
R6785 VDD.n324 VDD.n323 8.239
R6786 VDD.n1768 VDD.n1767 8.239
R6787 VDD.n1439 VDD.n1438 8.239
R6788 VDD.n2191 VDD.n2190 8.239
R6789 VDD.n535 VDD.n464 8.188
R6790 VDD.n1016 VDD.n932 8.188
R6791 VDD.n2259 VDD.n2227 8.188
R6792 VDD.n1528 VDD.n1496 8.182
R6793 VDD.n2938 VDD.n2430 8.182
R6794 VDD.n2691 VDD.n2564 8.176
R6795 VDD.n2691 VDD.n2585 8.176
R6796 VDD.n177 VDD.n99 8.176
R6797 VDD.n1736 VDD.n1704 8.176
R6798 VDD.n535 VDD.n406 8.1
R6799 VDD.n1016 VDD.n874 8.1
R6800 VDD.n2259 VDD.n2173 8.1
R6801 VDD.n1528 VDD.n1261 8.094
R6802 VDD.n2938 VDD.n2409 8.094
R6803 VDD.n177 VDD.n41 8.087
R6804 VDD.n1736 VDD.n774 8.087
R6805 VDD.n89 VDD.n88 8.076
R6806 VDD.n669 VDD.n668 8.076
R6807 VDD.n1150 VDD.n1149 8.076
R6808 VDD.n2538 VDD.n2537 8.076
R6809 VDD.n2603 VDD.n2602 8.076
R6810 VDD.n2082 VDD.n2081 8.076
R6811 VDD.n1694 VDD.n1693 8.076
R6812 VDD.n1486 VDD.n1485 8
R6813 VDD.n2981 VDD.n2980 8
R6814 VDD.n2448 VDD.n2447 8
R6815 VDD.n922 VDD.n921 7.924
R6816 VDD.n454 VDD.n453 7.924
R6817 VDD.n311 VDD.n310 7.924
R6818 VDD.n2735 VDD.n2734 7.924
R6819 VDD.n2828 VDD.n2827 7.924
R6820 VDD.n1779 VDD.n1778 7.924
R6821 VDD.n1426 VDD.n1425 7.924
R6822 VDD.n2217 VDD.n2216 7.924
R6823 VDD.n8 VDD.n7 7.208
R6824 VDD.n543 VDD.n542 7.208
R6825 VDD.n1024 VDD.n1023 7.208
R6826 VDD.n2509 VDD.n2508 7.208
R6827 VDD.n2626 VDD.n2625 7.208
R6828 VDD.n2625 VDD.n2624 7.208
R6829 VDD.n2510 VDD.n2509 7.208
R6830 VDD.n1023 VDD.n1022 7.208
R6831 VDD.n542 VDD.n541 7.208
R6832 VDD.n7 VDD.n6 7.208
R6833 VDD.n1956 VDD.n1955 7.208
R6834 VDD.n729 VDD.n728 7.208
R6835 VDD.n728 VDD.n727 7.208
R6836 VDD.n1955 VDD.n1954 7.208
R6837 VDD.n1216 VDD.n1215 7.142
R6838 VDD.n3109 VDD.n3108 7.142
R6839 VDD.n3108 VDD.n3107 7.142
R6840 VDD.n1215 VDD.n1214 7.142
R6841 VDD.n2471 VDD.n2470 7.142
R6842 VDD.n2470 VDD.n2469 7.142
R6843 VDD.n841 VDD.n840 7.077
R6844 VDD.n373 VDD.n372 7.077
R6845 VDD.n185 VDD.n184 7.077
R6846 VDD.n184 VDD.n183 7.077
R6847 VDD.n372 VDD.n371 7.077
R6848 VDD.n840 VDD.n839 7.077
R6849 VDD.n2866 VDD.n2865 7.077
R6850 VDD.n2865 VDD.n2864 7.077
R6851 VDD.n1907 VDD.n1906 7.077
R6852 VDD.n1300 VDD.n1299 7.077
R6853 VDD.n2128 VDD.n2127 7.077
R6854 VDD.n2127 VDD.n2126 7.077
R6855 VDD.n1299 VDD.n1298 7.077
R6856 VDD.n1906 VDD.n1905 7.077
R6857 VDD.n181 VDD.n180 7.035
R6858 VDD.n1740 VDD.n1739 7.035
R6859 VDD.n2695 VDD.n2694 6.952
R6860 VDD.n1467 VDD.n1466 6.952
R6861 VDD.n2942 VDD.n2941 6.952
R6862 VDD.n138 VDD.n132 6.923
R6863 VDD.n556 VDD.n555 6.923
R6864 VDD.n1037 VDD.n1036 6.923
R6865 VDD.n1969 VDD.n1968 6.923
R6866 VDD.n1731 VDD.n1725 6.923
R6867 VDD.n539 VDD.n538 6.871
R6868 VDD.n1020 VDD.n1019 6.871
R6869 VDD.n2123 VDD.n2122 6.871
R6870 VDD.n1523 VDD.n1517 6.857
R6871 VDD.n3098 VDD.n3097 6.857
R6872 VDD.n2361 VDD.n2355 6.857
R6873 VDD.n971 VDD.n965 6.792
R6874 VDD.n503 VDD.n497 6.792
R6875 VDD.n198 VDD.n197 6.792
R6876 VDD.n1896 VDD.n1895 6.792
R6877 VDD.n1313 VDD.n1312 6.792
R6878 VDD.n2254 VDD.n2248 6.792
R6879 VDD.n2938 VDD.n2440 6.751
R6880 VDD.n2938 VDD.n2459 6.751
R6881 VDD.n2938 VDD.n2478 6.751
R6882 VDD.n2938 VDD.n2362 6.751
R6883 VDD.n2938 VDD.n2381 6.751
R6884 VDD.n2938 VDD.n2400 6.751
R6885 VDD.n2691 VDD.n2536 6.736
R6886 VDD.n2691 VDD.n2555 6.736
R6887 VDD.n2691 VDD.n2595 6.736
R6888 VDD.n2691 VDD.n2614 6.736
R6889 VDD.n2691 VDD.n2633 6.736
R6890 VDD.n2691 VDD.n2517 6.736
R6891 VDD.n81 VDD.n80 6.365
R6892 VDD.n694 VDD.n693 6.365
R6893 VDD.n1175 VDD.n1174 6.365
R6894 VDD.n2526 VDD.n2519 6.365
R6895 VDD.n2623 VDD.n2622 6.365
R6896 VDD.n2107 VDD.n2106 6.365
R6897 VDD.n1686 VDD.n1685 6.365
R6898 VDD.n1478 VDD.n1477 6.307
R6899 VDD.n2958 VDD.n2957 6.307
R6900 VDD.n2468 VDD.n2467 6.307
R6901 VDD.n914 VDD.n913 6.249
R6902 VDD.n446 VDD.n445 6.249
R6903 VDD.n336 VDD.n335 6.249
R6904 VDD.n2711 VDD.n2710 6.249
R6905 VDD.n2854 VDD.n2853 6.249
R6906 VDD.n1756 VDD.n1755 6.249
R6907 VDD.n1451 VDD.n1450 6.249
R6908 VDD.n2209 VDD.n2208 6.249
R6909 VDD.n1738 VDD.n1737 6.168
R6910 VDD.n2693 VDD.n2692 6.168
R6911 VDD.n535 VDD.n437 6.168
R6912 VDD.n1016 VDD.n905 6.168
R6913 VDD.n2260 VDD.n2259 6.168
R6914 VDD.n1469 VDD.n1468 6.168
R6915 VDD.n2938 VDD.n2343 6.154
R6916 VDD.n2940 VDD.n2939 6.154
R6917 VDD.n1529 VDD.n1528 6.154
R6918 VDD.n177 VDD.n72 6.14
R6919 VDD.n1736 VDD.n1677 6.14
R6920 VDD.n2125 VDD.n2124 6.14
R6921 VDD.n132 VDD.n131 6.136
R6922 VDD.n555 VDD.n554 6.136
R6923 VDD.n1036 VDD.n1035 6.136
R6924 VDD.n1035 VDD.n1034 6.136
R6925 VDD.n554 VDD.n553 6.136
R6926 VDD.n131 VDD.n130 6.136
R6927 VDD.n1968 VDD.n1967 6.136
R6928 VDD.n1725 VDD.n1724 6.136
R6929 VDD.n1724 VDD.n1723 6.136
R6930 VDD.n1967 VDD.n1966 6.136
R6931 VDD.n1517 VDD.n1516 6.079
R6932 VDD.n3097 VDD.n3096 6.079
R6933 VDD.n3096 VDD.n3095 6.079
R6934 VDD.n1516 VDD.n1515 6.079
R6935 VDD.n2354 VDD.n2353 6.079
R6936 VDD.n2355 VDD.n2354 6.079
R6937 VDD.n965 VDD.n964 6.024
R6938 VDD.n497 VDD.n496 6.024
R6939 VDD.n197 VDD.n196 6.024
R6940 VDD.n196 VDD.n195 6.024
R6941 VDD.n496 VDD.n495 6.024
R6942 VDD.n964 VDD.n963 6.024
R6943 VDD.n1895 VDD.n1894 6.024
R6944 VDD.n1312 VDD.n1311 6.024
R6945 VDD.n2248 VDD.n2247 6.024
R6946 VDD.n2247 VDD.n2246 6.024
R6947 VDD.n1311 VDD.n1310 6.024
R6948 VDD.n1894 VDD.n1893 6.024
R6949 VDD.n49 VDD.n48 5.769
R6950 VDD.n657 VDD.n656 5.769
R6951 VDD.n1138 VDD.n1137 5.769
R6952 VDD.n2070 VDD.n2069 5.769
R6953 VDD.n782 VDD.n781 5.769
R6954 VDD.n1269 VDD.n1268 5.714
R6955 VDD.n2993 VDD.n2992 5.714
R6956 VDD.n2383 VDD.n2382 5.714
R6957 VDD.n882 VDD.n881 5.66
R6958 VDD.n414 VDD.n413 5.66
R6959 VDD.n299 VDD.n298 5.66
R6960 VDD.n1791 VDD.n1790 5.66
R6961 VDD.n1414 VDD.n1413 5.66
R6962 VDD.n2181 VDD.n2180 5.66
R6963 VDD.n268 VDD.n267 5.463
R6964 VDD.n1825 VDD.n1824 5.463
R6965 VDD.n2415 VDD.n2414 5.463
R6966 VDD.n939 VDD.n938 5.397
R6967 VDD.n471 VDD.n470 5.397
R6968 VDD.n2784 VDD.n2783 5.397
R6969 VDD.n1381 VDD.n1380 5.397
R6970 VDD.n2159 VDD.n2158 5.397
R6971 VDD.n3027 VDD.n3026 5.397
R6972 VDD.n535 VDD.n476 5.355
R6973 VDD.n1016 VDD.n944 5.355
R6974 VDD.n2259 VDD.n2164 5.355
R6975 VDD.n1528 VDD.n1252 5.336
R6976 VDD.n2938 VDD.n2421 5.336
R6977 VDD.n106 VDD.n105 5.333
R6978 VDD.n626 VDD.n625 5.333
R6979 VDD.n1107 VDD.n1106 5.333
R6980 VDD.n2571 VDD.n2570 5.333
R6981 VDD.n2037 VDD.n2036 5.333
R6982 VDD.n760 VDD.n759 5.333
R6983 VDD.n1247 VDD.n1246 5.333
R6984 VDD.n2691 VDD.n2576 5.317
R6985 VDD.n177 VDD.n111 5.317
R6986 VDD.n1736 VDD.n765 5.317
R6987 VDD.n17 VDD.n16 5.051
R6988 VDD.n567 VDD.n566 5.051
R6989 VDD.n1048 VDD.n1047 5.051
R6990 VDD.n2528 VDD.n2527 5.051
R6991 VDD.n2607 VDD.n2606 5.051
R6992 VDD.n2529 VDD.n2528 5.051
R6993 VDD.n2606 VDD.n2605 5.051
R6994 VDD.n1047 VDD.n1046 5.051
R6995 VDD.n566 VDD.n565 5.051
R6996 VDD.n16 VDD.n15 5.051
R6997 VDD.n1980 VDD.n1979 5.051
R6998 VDD.n738 VDD.n737 5.051
R6999 VDD.n737 VDD.n736 5.051
R7000 VDD.n1979 VDD.n1978 5.051
R7001 VDD.n1225 VDD.n1224 5.004
R7002 VDD.n3085 VDD.n3084 5.004
R7003 VDD.n3084 VDD.n3083 5.004
R7004 VDD.n1224 VDD.n1223 5.004
R7005 VDD.n2452 VDD.n2451 5.004
R7006 VDD.n2451 VDD.n2450 5.004
R7007 VDD.n850 VDD.n849 4.958
R7008 VDD.n382 VDD.n381 4.958
R7009 VDD.n209 VDD.n208 4.958
R7010 VDD.n208 VDD.n207 4.958
R7011 VDD.n381 VDD.n380 4.958
R7012 VDD.n849 VDD.n848 4.958
R7013 VDD.n2722 VDD.n2721 4.958
R7014 VDD.n2841 VDD.n2840 4.958
R7015 VDD.n2723 VDD.n2722 4.958
R7016 VDD.n2840 VDD.n2839 4.958
R7017 VDD.n1883 VDD.n1882 4.958
R7018 VDD.n1324 VDD.n1323 4.958
R7019 VDD.n2137 VDD.n2136 4.958
R7020 VDD.n2136 VDD.n2135 4.958
R7021 VDD.n1323 VDD.n1322 4.958
R7022 VDD.n1882 VDD.n1881 4.958
R7023 VDD.n14 VDD.n8 4.615
R7024 VDD.n544 VDD.n543 4.615
R7025 VDD.n1025 VDD.n1024 4.615
R7026 VDD.n2516 VDD.n2510 4.615
R7027 VDD.n2632 VDD.n2626 4.615
R7028 VDD.n1957 VDD.n1956 4.615
R7029 VDD.n735 VDD.n729 4.615
R7030 VDD.n1222 VDD.n1216 4.571
R7031 VDD.n3110 VDD.n3109 4.571
R7032 VDD.n2477 VDD.n2471 4.571
R7033 VDD.n847 VDD.n841 4.528
R7034 VDD.n379 VDD.n373 4.528
R7035 VDD.n186 VDD.n185 4.528
R7036 VDD.n2700 VDD.n2698 4.528
R7037 VDD.n2868 VDD.n2866 4.528
R7038 VDD.n1908 VDD.n1907 4.528
R7039 VDD.n1301 VDD.n1300 4.528
R7040 VDD.n2134 VDD.n2128 4.528
R7041 VDD.n68 VDD.n67 4.293
R7042 VDD.n706 VDD.n705 4.293
R7043 VDD.n1187 VDD.n1186 4.293
R7044 VDD.n2118 VDD.n2117 4.293
R7045 VDD.n801 VDD.n800 4.293
R7046 VDD.n1288 VDD.n1287 4.253
R7047 VDD.n2946 VDD.n2945 4.253
R7048 VDD.n2352 VDD.n2345 4.253
R7049 VDD.n901 VDD.n900 4.214
R7050 VDD.n433 VDD.n432 4.214
R7051 VDD.n348 VDD.n347 4.214
R7052 VDD.n1744 VDD.n1743 4.214
R7053 VDD.n1462 VDD.n1461 4.214
R7054 VDD.n2200 VDD.n2199 4.214
R7055 VDD.n123 VDD.n122 3.952
R7056 VDD.n579 VDD.n578 3.952
R7057 VDD.n1060 VDD.n1059 3.952
R7058 VDD.n1059 VDD.n1058 3.952
R7059 VDD.n578 VDD.n577 3.952
R7060 VDD.n122 VDD.n121 3.952
R7061 VDD.n1992 VDD.n1991 3.952
R7062 VDD.n1716 VDD.n1715 3.952
R7063 VDD.n1715 VDD.n1714 3.952
R7064 VDD.n1991 VDD.n1990 3.952
R7065 VDD.n1508 VDD.n1507 3.916
R7066 VDD.n3073 VDD.n3072 3.916
R7067 VDD.n3072 VDD.n3071 3.916
R7068 VDD.n1507 VDD.n1506 3.916
R7069 VDD.n2373 VDD.n2372 3.916
R7070 VDD.n2374 VDD.n2373 3.916
R7071 VDD.n956 VDD.n955 3.879
R7072 VDD.n488 VDD.n487 3.879
R7073 VDD.n221 VDD.n220 3.879
R7074 VDD.n220 VDD.n219 3.879
R7075 VDD.n487 VDD.n486 3.879
R7076 VDD.n955 VDD.n954 3.879
R7077 VDD.n1871 VDD.n1870 3.879
R7078 VDD.n1336 VDD.n1335 3.879
R7079 VDD.n2239 VDD.n2238 3.879
R7080 VDD.n2238 VDD.n2237 3.879
R7081 VDD.n1335 VDD.n1334 3.879
R7082 VDD.n1870 VDD.n1869 3.879
R7083 VDD.n98 VDD.n97 3.461
R7084 VDD.n645 VDD.n644 3.461
R7085 VDD.n1126 VDD.n1125 3.461
R7086 VDD.n2557 VDD.n2556 3.461
R7087 VDD.n2584 VDD.n2583 3.461
R7088 VDD.n2058 VDD.n2057 3.461
R7089 VDD.n1703 VDD.n1702 3.461
R7090 VDD.n2576 VDD.n2574 3.449
R7091 VDD.n1099 VDD.n1098 3.449
R7092 VDD.n618 VDD.n617 3.449
R7093 VDD.n111 VDD.n109 3.449
R7094 VDD.n2031 VDD.n2030 3.449
R7095 VDD.n765 VDD.n763 3.449
R7096 VDD.n1252 VDD.n1250 3.428
R7097 VDD.n3038 VDD.n3037 3.428
R7098 VDD.n2421 VDD.n2420 3.428
R7099 VDD.n1495 VDD.n1494 3.428
R7100 VDD.n3005 VDD.n3004 3.428
R7101 VDD.n2429 VDD.n2428 3.428
R7102 VDD.n260 VDD.n259 3.408
R7103 VDD.n476 VDD.n474 3.408
R7104 VDD.n944 VDD.n942 3.408
R7105 VDD.n2776 VDD.n2775 3.408
R7106 VDD.n1836 VDD.n1835 3.408
R7107 VDD.n1375 VDD.n1374 3.408
R7108 VDD.n2164 VDD.n2162 3.408
R7109 VDD.n931 VDD.n930 3.396
R7110 VDD.n463 VDD.n462 3.396
R7111 VDD.n287 VDD.n286 3.396
R7112 VDD.n2760 VDD.n2759 3.396
R7113 VDD.n2803 VDD.n2802 3.396
R7114 VDD.n1803 VDD.n1802 3.396
R7115 VDD.n1402 VDD.n1401 3.396
R7116 VDD.n2226 VDD.n2225 3.396
R7117 VDD.n26 VDD.n25 2.841
R7118 VDD.n591 VDD.n590 2.841
R7119 VDD.n1072 VDD.n1071 2.841
R7120 VDD.n2547 VDD.n2546 2.841
R7121 VDD.n2588 VDD.n2587 2.841
R7122 VDD.n2548 VDD.n2547 2.841
R7123 VDD.n2587 VDD.n2586 2.841
R7124 VDD.n1071 VDD.n1070 2.841
R7125 VDD.n590 VDD.n589 2.841
R7126 VDD.n25 VDD.n24 2.841
R7127 VDD.n2004 VDD.n2003 2.841
R7128 VDD.n747 VDD.n746 2.841
R7129 VDD.n746 VDD.n745 2.841
R7130 VDD.n2003 VDD.n2002 2.841
R7131 VDD.n1234 VDD.n1233 2.814
R7132 VDD.n3061 VDD.n3060 2.814
R7133 VDD.n3060 VDD.n3059 2.814
R7134 VDD.n1233 VDD.n1232 2.814
R7135 VDD.n2433 VDD.n2432 2.814
R7136 VDD.n2432 VDD.n2431 2.814
R7137 VDD.n859 VDD.n858 2.788
R7138 VDD.n391 VDD.n390 2.788
R7139 VDD.n233 VDD.n232 2.788
R7140 VDD.n232 VDD.n231 2.788
R7141 VDD.n390 VDD.n389 2.788
R7142 VDD.n858 VDD.n857 2.788
R7143 VDD.n2747 VDD.n2746 2.788
R7144 VDD.n2816 VDD.n2815 2.788
R7145 VDD.n2748 VDD.n2747 2.788
R7146 VDD.n2815 VDD.n2814 2.788
R7147 VDD.n1859 VDD.n1858 2.788
R7148 VDD.n1348 VDD.n1347 2.788
R7149 VDD.n2146 VDD.n2145 2.788
R7150 VDD.n2145 VDD.n2144 2.788
R7151 VDD.n1347 VDD.n1346 2.788
R7152 VDD.n1858 VDD.n1857 2.788
R7153 VDD.n175 VDD.n174 2.721
R7154 VDD.n546 VDD.n539 2.721
R7155 VDD.n1027 VDD.n1020 2.721
R7156 VDD.n2689 VDD.n2688 2.721
R7157 VDD.n2123 VDD.n2121 2.721
R7158 VDD.n1676 VDD.n1675 2.721
R7159 VDD.n1531 VDD.n1530 2.721
R7160 VDD.n1014 VDD.n1013 2.716
R7161 VDD.n533 VDD.n532 2.716
R7162 VDD.n2702 VDD.n2695 2.716
R7163 VDD.n1467 VDD.n1465 2.716
R7164 VDD.n2262 VDD.n2261 2.716
R7165 VDD.n2949 VDD.n2942 2.716
R7166 VDD.n188 VDD.n181 2.711
R7167 VDD.n1747 VDD.n1740 2.711
R7168 VDD.n2936 VDD.n2935 2.711
R7169 VDD.n261 VDD.n254 2.497
R7170 VDD.n278 VDD.n273 2.497
R7171 VDD.n1837 VDD.n1830 2.497
R7172 VDD.n1818 VDD.n1813 2.497
R7173 VDD.n2407 VDD.n2404 2.497
R7174 VDD.n2407 VDD.n2406 2.497
R7175 VDD.n2419 VDD.n2416 2.497
R7176 VDD.n2419 VDD.n2418 2.497
R7177 VDD.n941 VDD.n937 2.467
R7178 VDD.n941 VDD.n940 2.467
R7179 VDD.n870 VDD.n867 2.467
R7180 VDD.n870 VDD.n869 2.467
R7181 VDD.n473 VDD.n469 2.467
R7182 VDD.n473 VDD.n472 2.467
R7183 VDD.n402 VDD.n399 2.467
R7184 VDD.n402 VDD.n401 2.467
R7185 VDD.n2777 VDD.n2770 2.467
R7186 VDD.n2794 VDD.n2789 2.467
R7187 VDD.n1376 VDD.n1369 2.467
R7188 VDD.n1393 VDD.n1388 2.467
R7189 VDD.n2161 VDD.n2157 2.467
R7190 VDD.n2161 VDD.n2160 2.467
R7191 VDD.n2169 VDD.n2166 2.467
R7192 VDD.n2169 VDD.n2168 2.467
R7193 VDD.n3039 VDD.n3032 2.467
R7194 VDD.n3020 VDD.n3015 2.467
R7195 VDD.n108 VDD.n104 2.438
R7196 VDD.n108 VDD.n107 2.438
R7197 VDD.n37 VDD.n34 2.438
R7198 VDD.n37 VDD.n36 2.438
R7199 VDD.n619 VDD.n612 2.438
R7200 VDD.n636 VDD.n631 2.438
R7201 VDD.n1100 VDD.n1093 2.438
R7202 VDD.n1117 VDD.n1112 2.438
R7203 VDD.n2573 VDD.n2569 2.438
R7204 VDD.n2573 VDD.n2572 2.438
R7205 VDD.n2645 VDD.n2642 2.438
R7206 VDD.n2645 VDD.n2644 2.438
R7207 VDD.n2032 VDD.n2025 2.438
R7208 VDD.n2049 VDD.n2044 2.438
R7209 VDD.n762 VDD.n758 2.438
R7210 VDD.n762 VDD.n761 2.438
R7211 VDD.n770 VDD.n767 2.438
R7212 VDD.n770 VDD.n769 2.438
R7213 VDD.n1249 VDD.n1245 2.438
R7214 VDD.n1249 VDD.n1248 2.438
R7215 VDD.n1257 VDD.n1254 2.438
R7216 VDD.n1257 VDD.n1256 2.438
R7217 VDD.n2341 VDD.n2340 2.341
R7218 VDD.n903 VDD.n902 2.313
R7219 VDD.n435 VDD.n434 2.313
R7220 VDD.n2256 VDD.n2255 2.313
R7221 VDD.n70 VDD.n69 2.285
R7222 VDD.n2635 VDD.n2634 2.285
R7223 VDD.n1733 VDD.n1732 2.285
R7224 VDD.n1525 VDD.n1524 2.285
R7225 VDD.n2517 VDD.n2516 2.227
R7226 VDD.n2536 VDD.n2535 2.227
R7227 VDD.n2555 VDD.n2554 2.227
R7228 VDD.n2595 VDD.n2594 2.227
R7229 VDD.n2614 VDD.n2613 2.227
R7230 VDD.n2633 VDD.n2632 2.227
R7231 VDD.n2362 VDD.n2361 2.211
R7232 VDD.n2381 VDD.n2380 2.211
R7233 VDD.n2400 VDD.n2399 2.211
R7234 VDD.n2440 VDD.n2439 2.211
R7235 VDD.n2459 VDD.n2458 2.211
R7236 VDD.n2478 VDD.n2477 2.211
R7237 VDD.n2700 VDD.n2699 2.195
R7238 VDD.n2725 VDD.n2724 2.195
R7239 VDD.n2750 VDD.n2749 2.195
R7240 VDD.n2818 VDD.n2817 2.195
R7241 VDD.n2843 VDD.n2842 2.195
R7242 VDD.n2868 VDD.n2867 2.195
R7243 VDD.n247 VDD.n242 2.185
R7244 VDD.n290 VDD.n285 2.185
R7245 VDD.n1849 VDD.n1844 2.185
R7246 VDD.n1806 VDD.n1801 2.185
R7247 VDD.n2398 VDD.n2395 2.185
R7248 VDD.n2398 VDD.n2397 2.185
R7249 VDD.n2426 VDD.n2423 2.185
R7250 VDD.n2426 VDD.n2425 2.185
R7251 VDD.n952 VDD.n949 2.159
R7252 VDD.n952 VDD.n951 2.159
R7253 VDD.n928 VDD.n925 2.159
R7254 VDD.n928 VDD.n927 2.159
R7255 VDD.n484 VDD.n481 2.159
R7256 VDD.n484 VDD.n483 2.159
R7257 VDD.n460 VDD.n457 2.159
R7258 VDD.n460 VDD.n459 2.159
R7259 VDD.n2763 VDD.n2758 2.159
R7260 VDD.n2806 VDD.n2801 2.159
R7261 VDD.n1362 VDD.n1357 2.159
R7262 VDD.n1405 VDD.n1400 2.159
R7263 VDD.n2235 VDD.n2232 2.159
R7264 VDD.n2235 VDD.n2234 2.159
R7265 VDD.n2223 VDD.n2220 2.159
R7266 VDD.n2223 VDD.n2222 2.159
R7267 VDD.n3051 VDD.n3046 2.159
R7268 VDD.n3008 VDD.n3003 2.159
R7269 VDD.n119 VDD.n116 2.133
R7270 VDD.n119 VDD.n118 2.133
R7271 VDD.n95 VDD.n92 2.133
R7272 VDD.n95 VDD.n94 2.133
R7273 VDD.n605 VDD.n600 2.133
R7274 VDD.n648 VDD.n643 2.133
R7275 VDD.n1086 VDD.n1081 2.133
R7276 VDD.n1129 VDD.n1124 2.133
R7277 VDD.n2562 VDD.n2559 2.133
R7278 VDD.n2562 VDD.n2561 2.133
R7279 VDD.n2581 VDD.n2578 2.133
R7280 VDD.n2581 VDD.n2580 2.133
R7281 VDD.n2018 VDD.n2013 2.133
R7282 VDD.n2061 VDD.n2056 2.133
R7283 VDD.n1712 VDD.n1709 2.133
R7284 VDD.n1712 VDD.n1711 2.133
R7285 VDD.n1700 VDD.n1697 2.133
R7286 VDD.n1700 VDD.n1699 2.133
R7287 VDD.n1504 VDD.n1501 2.133
R7288 VDD.n1504 VDD.n1503 2.133
R7289 VDD.n1492 VDD.n1489 2.133
R7290 VDD.n1492 VDD.n1491 2.133
R7291 VDD.n345 VDD.n344 2.029
R7292 VDD.n1904 VDD.n1903 2.029
R7293 VDD.n2347 VDD.n2346 2.029
R7294 VDD.n2349 VDD.n2348 2.029
R7295 VDD.n2473 VDD.n2472 2.029
R7296 VDD.n2475 VDD.n2474 2.029
R7297 VDD.n843 VDD.n842 2.004
R7298 VDD.n845 VDD.n844 2.004
R7299 VDD.n894 VDD.n893 2.004
R7300 VDD.n896 VDD.n895 2.004
R7301 VDD.n375 VDD.n374 2.004
R7302 VDD.n377 VDD.n376 2.004
R7303 VDD.n426 VDD.n425 2.004
R7304 VDD.n428 VDD.n427 2.004
R7305 VDD.n2863 VDD.n2862 2.004
R7306 VDD.n1297 VDD.n1296 2.004
R7307 VDD.n2130 VDD.n2129 2.004
R7308 VDD.n2132 VDD.n2131 2.004
R7309 VDD.n2193 VDD.n2192 2.004
R7310 VDD.n2195 VDD.n2194 2.004
R7311 VDD.n3106 VDD.n3105 2.004
R7312 VDD.n10 VDD.n9 1.98
R7313 VDD.n12 VDD.n11 1.98
R7314 VDD.n61 VDD.n60 1.98
R7315 VDD.n63 VDD.n62 1.98
R7316 VDD.n703 VDD.n702 1.98
R7317 VDD.n1184 VDD.n1183 1.98
R7318 VDD.n2512 VDD.n2511 1.98
R7319 VDD.n2514 VDD.n2513 1.98
R7320 VDD.n2628 VDD.n2627 1.98
R7321 VDD.n2630 VDD.n2629 1.98
R7322 VDD.n1953 VDD.n1952 1.98
R7323 VDD.n731 VDD.n730 1.98
R7324 VDD.n733 VDD.n732 1.98
R7325 VDD.n794 VDD.n793 1.98
R7326 VDD.n796 VDD.n795 1.98
R7327 VDD.n1218 VDD.n1217 1.98
R7328 VDD.n1220 VDD.n1219 1.98
R7329 VDD.n1281 VDD.n1280 1.98
R7330 VDD.n1283 VDD.n1282 1.98
R7331 VDD.n235 VDD.n230 1.873
R7332 VDD.n302 VDD.n297 1.873
R7333 VDD.n1861 VDD.n1856 1.873
R7334 VDD.n1794 VDD.n1789 1.873
R7335 VDD.n2388 VDD.n2385 1.873
R7336 VDD.n2388 VDD.n2387 1.873
R7337 VDD.n2438 VDD.n2435 1.873
R7338 VDD.n2438 VDD.n2437 1.873
R7339 VDD.n864 VDD.n861 1.85
R7340 VDD.n864 VDD.n863 1.85
R7341 VDD.n879 VDD.n876 1.85
R7342 VDD.n879 VDD.n878 1.85
R7343 VDD.n396 VDD.n393 1.85
R7344 VDD.n396 VDD.n395 1.85
R7345 VDD.n411 VDD.n408 1.85
R7346 VDD.n411 VDD.n410 1.85
R7347 VDD.n2751 VDD.n2745 1.85
R7348 VDD.n2819 VDD.n2813 1.85
R7349 VDD.n1350 VDD.n1345 1.85
R7350 VDD.n1417 VDD.n1412 1.85
R7351 VDD.n2151 VDD.n2148 1.85
R7352 VDD.n2151 VDD.n2150 1.85
R7353 VDD.n2178 VDD.n2175 1.85
R7354 VDD.n2178 VDD.n2177 1.85
R7355 VDD.n3063 VDD.n3058 1.85
R7356 VDD.n2996 VDD.n2991 1.85
R7357 VDD.n31 VDD.n28 1.828
R7358 VDD.n31 VDD.n30 1.828
R7359 VDD.n46 VDD.n43 1.828
R7360 VDD.n46 VDD.n45 1.828
R7361 VDD.n593 VDD.n588 1.828
R7362 VDD.n660 VDD.n655 1.828
R7363 VDD.n1074 VDD.n1069 1.828
R7364 VDD.n1141 VDD.n1136 1.828
R7365 VDD.n2553 VDD.n2550 1.828
R7366 VDD.n2553 VDD.n2552 1.828
R7367 VDD.n2593 VDD.n2590 1.828
R7368 VDD.n2593 VDD.n2592 1.828
R7369 VDD.n2006 VDD.n2001 1.828
R7370 VDD.n2073 VDD.n2068 1.828
R7371 VDD.n752 VDD.n749 1.828
R7372 VDD.n752 VDD.n751 1.828
R7373 VDD.n779 VDD.n776 1.828
R7374 VDD.n779 VDD.n778 1.828
R7375 VDD.n1239 VDD.n1236 1.828
R7376 VDD.n1239 VDD.n1238 1.828
R7377 VDD.n1266 VDD.n1263 1.828
R7378 VDD.n1266 VDD.n1265 1.828
R7379 VDD.n194 VDD.n193 1.717
R7380 VDD.n333 VDD.n332 1.717
R7381 VDD.n1892 VDD.n1891 1.717
R7382 VDD.n1753 VDD.n1752 1.717
R7383 VDD.n2357 VDD.n2356 1.717
R7384 VDD.n2359 VDD.n2358 1.717
R7385 VDD.n2461 VDD.n2460 1.717
R7386 VDD.n2463 VDD.n2462 1.717
R7387 VDD.n114 VDD.n113 1.715
R7388 VDD.n603 VDD.n602 1.715
R7389 VDD.n1084 VDD.n1083 1.715
R7390 VDD.n1083 VDD.n1082 1.715
R7391 VDD.n602 VDD.n601 1.715
R7392 VDD.n113 VDD.n112 1.715
R7393 VDD.n2016 VDD.n2015 1.715
R7394 VDD.n1707 VDD.n1706 1.715
R7395 VDD.n1706 VDD.n1705 1.715
R7396 VDD.n2015 VDD.n2014 1.715
R7397 VDD.n1499 VDD.n1498 1.699
R7398 VDD.n3049 VDD.n3048 1.699
R7399 VDD.n3048 VDD.n3047 1.699
R7400 VDD.n1498 VDD.n1497 1.699
R7401 VDD.n2392 VDD.n2391 1.699
R7402 VDD.n2393 VDD.n2392 1.699
R7403 VDD.n967 VDD.n966 1.696
R7404 VDD.n969 VDD.n968 1.696
R7405 VDD.n907 VDD.n906 1.696
R7406 VDD.n909 VDD.n908 1.696
R7407 VDD.n499 VDD.n498 1.696
R7408 VDD.n501 VDD.n500 1.696
R7409 VDD.n439 VDD.n438 1.696
R7410 VDD.n441 VDD.n440 1.696
R7411 VDD.n2708 VDD.n2707 1.696
R7412 VDD.n2851 VDD.n2850 1.696
R7413 VDD.n1309 VDD.n1308 1.696
R7414 VDD.n1448 VDD.n1447 1.696
R7415 VDD.n2250 VDD.n2249 1.696
R7416 VDD.n2252 VDD.n2251 1.696
R7417 VDD.n2202 VDD.n2201 1.696
R7418 VDD.n2204 VDD.n2203 1.696
R7419 VDD.n3094 VDD.n3093 1.696
R7420 VDD.n2955 VDD.n2954 1.696
R7421 VDD.n947 VDD.n946 1.683
R7422 VDD.n479 VDD.n478 1.683
R7423 VDD.n245 VDD.n244 1.683
R7424 VDD.n244 VDD.n243 1.683
R7425 VDD.n478 VDD.n477 1.683
R7426 VDD.n946 VDD.n945 1.683
R7427 VDD.n1847 VDD.n1846 1.683
R7428 VDD.n1360 VDD.n1359 1.683
R7429 VDD.n2230 VDD.n2229 1.683
R7430 VDD.n2229 VDD.n2228 1.683
R7431 VDD.n1359 VDD.n1358 1.683
R7432 VDD.n1846 VDD.n1845 1.683
R7433 VDD.n134 VDD.n133 1.676
R7434 VDD.n136 VDD.n135 1.676
R7435 VDD.n74 VDD.n73 1.676
R7436 VDD.n76 VDD.n75 1.676
R7437 VDD.n552 VDD.n551 1.676
R7438 VDD.n691 VDD.n690 1.676
R7439 VDD.n1033 VDD.n1032 1.676
R7440 VDD.n1172 VDD.n1171 1.676
R7441 VDD.n2521 VDD.n2520 1.676
R7442 VDD.n2523 VDD.n2522 1.676
R7443 VDD.n2616 VDD.n2615 1.676
R7444 VDD.n2618 VDD.n2617 1.676
R7445 VDD.n1965 VDD.n1964 1.676
R7446 VDD.n2104 VDD.n2103 1.676
R7447 VDD.n1727 VDD.n1726 1.676
R7448 VDD.n1729 VDD.n1728 1.676
R7449 VDD.n1679 VDD.n1678 1.676
R7450 VDD.n1681 VDD.n1680 1.676
R7451 VDD.n1519 VDD.n1518 1.676
R7452 VDD.n1521 VDD.n1520 1.676
R7453 VDD.n1471 VDD.n1470 1.676
R7454 VDD.n1473 VDD.n1472 1.676
R7455 VDD.n223 VDD.n218 1.56
R7456 VDD.n314 VDD.n309 1.56
R7457 VDD.n1873 VDD.n1868 1.56
R7458 VDD.n1782 VDD.n1777 1.56
R7459 VDD.n2379 VDD.n2376 1.56
R7460 VDD.n2379 VDD.n2378 1.56
R7461 VDD.n2445 VDD.n2442 1.56
R7462 VDD.n2445 VDD.n2444 1.56
R7463 VDD.n961 VDD.n958 1.542
R7464 VDD.n961 VDD.n960 1.542
R7465 VDD.n919 VDD.n916 1.542
R7466 VDD.n919 VDD.n918 1.542
R7467 VDD.n493 VDD.n490 1.542
R7468 VDD.n493 VDD.n492 1.542
R7469 VDD.n451 VDD.n448 1.542
R7470 VDD.n451 VDD.n450 1.542
R7471 VDD.n2738 VDD.n2733 1.542
R7472 VDD.n2831 VDD.n2826 1.542
R7473 VDD.n1338 VDD.n1333 1.542
R7474 VDD.n1429 VDD.n1424 1.542
R7475 VDD.n2244 VDD.n2241 1.542
R7476 VDD.n2244 VDD.n2243 1.542
R7477 VDD.n2214 VDD.n2211 1.542
R7478 VDD.n2214 VDD.n2213 1.542
R7479 VDD.n3075 VDD.n3070 1.542
R7480 VDD.n2984 VDD.n2979 1.542
R7481 VDD.n128 VDD.n125 1.523
R7482 VDD.n128 VDD.n127 1.523
R7483 VDD.n86 VDD.n83 1.523
R7484 VDD.n86 VDD.n85 1.523
R7485 VDD.n581 VDD.n576 1.523
R7486 VDD.n672 VDD.n667 1.523
R7487 VDD.n1062 VDD.n1057 1.523
R7488 VDD.n1153 VDD.n1148 1.523
R7489 VDD.n2543 VDD.n2540 1.523
R7490 VDD.n2543 VDD.n2542 1.523
R7491 VDD.n2600 VDD.n2597 1.523
R7492 VDD.n2600 VDD.n2599 1.523
R7493 VDD.n1994 VDD.n1989 1.523
R7494 VDD.n2085 VDD.n2080 1.523
R7495 VDD.n1721 VDD.n1718 1.523
R7496 VDD.n1721 VDD.n1720 1.523
R7497 VDD.n1691 VDD.n1688 1.523
R7498 VDD.n1691 VDD.n1690 1.523
R7499 VDD.n1513 VDD.n1510 1.523
R7500 VDD.n1513 VDD.n1512 1.523
R7501 VDD.n1483 VDD.n1480 1.523
R7502 VDD.n1483 VDD.n1482 1.523
R7503 VDD.n206 VDD.n205 1.404
R7504 VDD.n321 VDD.n320 1.404
R7505 VDD.n1880 VDD.n1879 1.404
R7506 VDD.n1765 VDD.n1764 1.404
R7507 VDD.n2366 VDD.n2365 1.404
R7508 VDD.n2368 VDD.n2367 1.404
R7509 VDD.n2454 VDD.n2453 1.404
R7510 VDD.n2456 VDD.n2455 1.404
R7511 VDD.n852 VDD.n851 1.387
R7512 VDD.n854 VDD.n853 1.387
R7513 VDD.n885 VDD.n884 1.387
R7514 VDD.n887 VDD.n886 1.387
R7515 VDD.n384 VDD.n383 1.387
R7516 VDD.n386 VDD.n385 1.387
R7517 VDD.n417 VDD.n416 1.387
R7518 VDD.n419 VDD.n418 1.387
R7519 VDD.n2720 VDD.n2719 1.387
R7520 VDD.n2838 VDD.n2837 1.387
R7521 VDD.n1321 VDD.n1320 1.387
R7522 VDD.n1436 VDD.n1435 1.387
R7523 VDD.n2139 VDD.n2138 1.387
R7524 VDD.n2141 VDD.n2140 1.387
R7525 VDD.n2184 VDD.n2183 1.387
R7526 VDD.n2186 VDD.n2185 1.387
R7527 VDD.n3082 VDD.n3081 1.387
R7528 VDD.n2967 VDD.n2966 1.387
R7529 VDD.n19 VDD.n18 1.371
R7530 VDD.n21 VDD.n20 1.371
R7531 VDD.n52 VDD.n51 1.371
R7532 VDD.n54 VDD.n53 1.371
R7533 VDD.n564 VDD.n563 1.371
R7534 VDD.n679 VDD.n678 1.371
R7535 VDD.n1045 VDD.n1044 1.371
R7536 VDD.n1160 VDD.n1159 1.371
R7537 VDD.n2531 VDD.n2530 1.371
R7538 VDD.n2533 VDD.n2532 1.371
R7539 VDD.n2609 VDD.n2608 1.371
R7540 VDD.n2611 VDD.n2610 1.371
R7541 VDD.n1977 VDD.n1976 1.371
R7542 VDD.n2092 VDD.n2091 1.371
R7543 VDD.n740 VDD.n739 1.371
R7544 VDD.n742 VDD.n741 1.371
R7545 VDD.n785 VDD.n784 1.371
R7546 VDD.n787 VDD.n786 1.371
R7547 VDD.n1227 VDD.n1226 1.371
R7548 VDD.n1229 VDD.n1228 1.371
R7549 VDD.n1272 VDD.n1271 1.371
R7550 VDD.n1274 VDD.n1273 1.371
R7551 VDD.n211 VDD.n206 1.248
R7552 VDD.n326 VDD.n321 1.248
R7553 VDD.n1885 VDD.n1880 1.248
R7554 VDD.n1770 VDD.n1765 1.248
R7555 VDD.n2369 VDD.n2366 1.248
R7556 VDD.n2369 VDD.n2368 1.248
R7557 VDD.n2457 VDD.n2454 1.248
R7558 VDD.n2457 VDD.n2456 1.248
R7559 VDD.n855 VDD.n852 1.233
R7560 VDD.n855 VDD.n854 1.233
R7561 VDD.n888 VDD.n885 1.233
R7562 VDD.n888 VDD.n887 1.233
R7563 VDD.n387 VDD.n384 1.233
R7564 VDD.n387 VDD.n386 1.233
R7565 VDD.n420 VDD.n417 1.233
R7566 VDD.n420 VDD.n419 1.233
R7567 VDD.n2726 VDD.n2720 1.233
R7568 VDD.n2844 VDD.n2838 1.233
R7569 VDD.n1326 VDD.n1321 1.233
R7570 VDD.n1441 VDD.n1436 1.233
R7571 VDD.n2142 VDD.n2139 1.233
R7572 VDD.n2142 VDD.n2141 1.233
R7573 VDD.n2187 VDD.n2184 1.233
R7574 VDD.n2187 VDD.n2186 1.233
R7575 VDD.n3087 VDD.n3082 1.233
R7576 VDD.n2972 VDD.n2967 1.233
R7577 VDD.n22 VDD.n19 1.219
R7578 VDD.n22 VDD.n21 1.219
R7579 VDD.n55 VDD.n52 1.219
R7580 VDD.n55 VDD.n54 1.219
R7581 VDD.n569 VDD.n564 1.219
R7582 VDD.n684 VDD.n679 1.219
R7583 VDD.n1050 VDD.n1045 1.219
R7584 VDD.n1165 VDD.n1160 1.219
R7585 VDD.n2534 VDD.n2531 1.219
R7586 VDD.n2534 VDD.n2533 1.219
R7587 VDD.n2612 VDD.n2609 1.219
R7588 VDD.n2612 VDD.n2611 1.219
R7589 VDD.n1982 VDD.n1977 1.219
R7590 VDD.n2097 VDD.n2092 1.219
R7591 VDD.n743 VDD.n740 1.219
R7592 VDD.n743 VDD.n742 1.219
R7593 VDD.n788 VDD.n785 1.219
R7594 VDD.n788 VDD.n787 1.219
R7595 VDD.n1230 VDD.n1227 1.219
R7596 VDD.n1230 VDD.n1229 1.219
R7597 VDD.n1275 VDD.n1272 1.219
R7598 VDD.n1275 VDD.n1274 1.219
R7599 VDD.n40 VDD.n39 1.153
R7600 VDD.n633 VDD.n632 1.153
R7601 VDD.n1114 VDD.n1113 1.153
R7602 VDD.n2046 VDD.n2045 1.153
R7603 VDD.n773 VDD.n772 1.153
R7604 VDD.n1260 VDD.n1259 1.142
R7605 VDD.n3017 VDD.n3016 1.142
R7606 VDD.n2402 VDD.n2401 1.142
R7607 VDD.n873 VDD.n872 1.132
R7608 VDD.n405 VDD.n404 1.132
R7609 VDD.n275 VDD.n274 1.132
R7610 VDD.n1815 VDD.n1814 1.132
R7611 VDD.n1390 VDD.n1389 1.132
R7612 VDD.n2172 VDD.n2171 1.132
R7613 VDD.n218 VDD.n217 1.092
R7614 VDD.n309 VDD.n308 1.092
R7615 VDD.n1868 VDD.n1867 1.092
R7616 VDD.n1777 VDD.n1776 1.092
R7617 VDD.n2376 VDD.n2375 1.092
R7618 VDD.n2378 VDD.n2377 1.092
R7619 VDD.n2442 VDD.n2441 1.092
R7620 VDD.n2444 VDD.n2443 1.092
R7621 VDD.n958 VDD.n957 1.079
R7622 VDD.n960 VDD.n959 1.079
R7623 VDD.n916 VDD.n915 1.079
R7624 VDD.n918 VDD.n917 1.079
R7625 VDD.n490 VDD.n489 1.079
R7626 VDD.n492 VDD.n491 1.079
R7627 VDD.n448 VDD.n447 1.079
R7628 VDD.n450 VDD.n449 1.079
R7629 VDD.n2733 VDD.n2732 1.079
R7630 VDD.n2826 VDD.n2825 1.079
R7631 VDD.n1333 VDD.n1332 1.079
R7632 VDD.n1424 VDD.n1423 1.079
R7633 VDD.n2241 VDD.n2240 1.079
R7634 VDD.n2243 VDD.n2242 1.079
R7635 VDD.n2211 VDD.n2210 1.079
R7636 VDD.n2213 VDD.n2212 1.079
R7637 VDD.n3070 VDD.n3069 1.079
R7638 VDD.n2979 VDD.n2978 1.079
R7639 VDD.n125 VDD.n124 1.066
R7640 VDD.n127 VDD.n126 1.066
R7641 VDD.n83 VDD.n82 1.066
R7642 VDD.n85 VDD.n84 1.066
R7643 VDD.n576 VDD.n575 1.066
R7644 VDD.n667 VDD.n666 1.066
R7645 VDD.n1057 VDD.n1056 1.066
R7646 VDD.n1148 VDD.n1147 1.066
R7647 VDD.n2540 VDD.n2539 1.066
R7648 VDD.n2542 VDD.n2541 1.066
R7649 VDD.n2597 VDD.n2596 1.066
R7650 VDD.n2599 VDD.n2598 1.066
R7651 VDD.n1989 VDD.n1988 1.066
R7652 VDD.n2080 VDD.n2079 1.066
R7653 VDD.n1718 VDD.n1717 1.066
R7654 VDD.n1720 VDD.n1719 1.066
R7655 VDD.n1688 VDD.n1687 1.066
R7656 VDD.n1690 VDD.n1689 1.066
R7657 VDD.n1510 VDD.n1509 1.066
R7658 VDD.n1512 VDD.n1511 1.066
R7659 VDD.n1480 VDD.n1479 1.066
R7660 VDD.n1482 VDD.n1481 1.066
R7661 VDD.n199 VDD.n194 0.936
R7662 VDD.n338 VDD.n333 0.936
R7663 VDD.n1897 VDD.n1892 0.936
R7664 VDD.n1758 VDD.n1753 0.936
R7665 VDD.n2360 VDD.n2357 0.936
R7666 VDD.n2360 VDD.n2359 0.936
R7667 VDD.n2464 VDD.n2461 0.936
R7668 VDD.n2464 VDD.n2463 0.936
R7669 VDD.n970 VDD.n967 0.925
R7670 VDD.n970 VDD.n969 0.925
R7671 VDD.n910 VDD.n907 0.925
R7672 VDD.n910 VDD.n909 0.925
R7673 VDD.n502 VDD.n499 0.925
R7674 VDD.n502 VDD.n501 0.925
R7675 VDD.n442 VDD.n439 0.925
R7676 VDD.n442 VDD.n441 0.925
R7677 VDD.n2713 VDD.n2708 0.925
R7678 VDD.n2856 VDD.n2851 0.925
R7679 VDD.n1314 VDD.n1309 0.925
R7680 VDD.n1453 VDD.n1448 0.925
R7681 VDD.n2253 VDD.n2250 0.925
R7682 VDD.n2253 VDD.n2252 0.925
R7683 VDD.n2205 VDD.n2202 0.925
R7684 VDD.n2205 VDD.n2204 0.925
R7685 VDD.n3099 VDD.n3094 0.925
R7686 VDD.n2960 VDD.n2955 0.925
R7687 VDD.n137 VDD.n134 0.914
R7688 VDD.n137 VDD.n136 0.914
R7689 VDD.n77 VDD.n74 0.914
R7690 VDD.n77 VDD.n76 0.914
R7691 VDD.n557 VDD.n552 0.914
R7692 VDD.n696 VDD.n691 0.914
R7693 VDD.n1038 VDD.n1033 0.914
R7694 VDD.n1177 VDD.n1172 0.914
R7695 VDD.n2524 VDD.n2521 0.914
R7696 VDD.n2524 VDD.n2523 0.914
R7697 VDD.n2619 VDD.n2616 0.914
R7698 VDD.n2619 VDD.n2618 0.914
R7699 VDD.n1970 VDD.n1965 0.914
R7700 VDD.n2109 VDD.n2104 0.914
R7701 VDD.n1730 VDD.n1727 0.914
R7702 VDD.n1730 VDD.n1729 0.914
R7703 VDD.n1682 VDD.n1679 0.914
R7704 VDD.n1682 VDD.n1681 0.914
R7705 VDD.n1522 VDD.n1519 0.914
R7706 VDD.n1522 VDD.n1521 0.914
R7707 VDD.n1474 VDD.n1471 0.914
R7708 VDD.n1474 VDD.n1473 0.914
R7709 VDD.n1116 VDD.n1115 0.807
R7710 VDD.n635 VDD.n634 0.807
R7711 VDD.n41 VDD.n38 0.807
R7712 VDD.n774 VDD.n771 0.807
R7713 VDD.n2048 VDD.n2047 0.807
R7714 VDD.n3019 VDD.n3018 0.8
R7715 VDD.n1261 VDD.n1258 0.8
R7716 VDD.n2409 VDD.n2408 0.8
R7717 VDD.n277 VDD.n276 0.794
R7718 VDD.n406 VDD.n403 0.794
R7719 VDD.n874 VDD.n871 0.794
R7720 VDD.n2173 VDD.n2170 0.794
R7721 VDD.n1392 VDD.n1391 0.794
R7722 VDD.n1817 VDD.n1816 0.794
R7723 VDD.n230 VDD.n229 0.78
R7724 VDD.n297 VDD.n296 0.78
R7725 VDD.n1856 VDD.n1855 0.78
R7726 VDD.n1789 VDD.n1788 0.78
R7727 VDD.n2385 VDD.n2384 0.78
R7728 VDD.n2387 VDD.n2386 0.78
R7729 VDD.n2435 VDD.n2434 0.78
R7730 VDD.n2437 VDD.n2436 0.78
R7731 VDD.n861 VDD.n860 0.771
R7732 VDD.n863 VDD.n862 0.771
R7733 VDD.n876 VDD.n875 0.771
R7734 VDD.n878 VDD.n877 0.771
R7735 VDD.n393 VDD.n392 0.771
R7736 VDD.n395 VDD.n394 0.771
R7737 VDD.n408 VDD.n407 0.771
R7738 VDD.n410 VDD.n409 0.771
R7739 VDD.n2745 VDD.n2744 0.771
R7740 VDD.n2813 VDD.n2812 0.771
R7741 VDD.n1345 VDD.n1344 0.771
R7742 VDD.n1412 VDD.n1411 0.771
R7743 VDD.n2148 VDD.n2147 0.771
R7744 VDD.n2150 VDD.n2149 0.771
R7745 VDD.n2175 VDD.n2174 0.771
R7746 VDD.n2177 VDD.n2176 0.771
R7747 VDD.n3058 VDD.n3057 0.771
R7748 VDD.n2991 VDD.n2990 0.771
R7749 VDD.n28 VDD.n27 0.761
R7750 VDD.n30 VDD.n29 0.761
R7751 VDD.n43 VDD.n42 0.761
R7752 VDD.n45 VDD.n44 0.761
R7753 VDD.n588 VDD.n587 0.761
R7754 VDD.n655 VDD.n654 0.761
R7755 VDD.n1069 VDD.n1068 0.761
R7756 VDD.n1136 VDD.n1135 0.761
R7757 VDD.n2550 VDD.n2549 0.761
R7758 VDD.n2552 VDD.n2551 0.761
R7759 VDD.n2590 VDD.n2589 0.761
R7760 VDD.n2592 VDD.n2591 0.761
R7761 VDD.n2001 VDD.n2000 0.761
R7762 VDD.n2068 VDD.n2067 0.761
R7763 VDD.n749 VDD.n748 0.761
R7764 VDD.n751 VDD.n750 0.761
R7765 VDD.n776 VDD.n775 0.761
R7766 VDD.n778 VDD.n777 0.761
R7767 VDD.n1236 VDD.n1235 0.761
R7768 VDD.n1238 VDD.n1237 0.761
R7769 VDD.n1263 VDD.n1262 0.761
R7770 VDD.n1265 VDD.n1264 0.761
R7771 VDD.n2585 VDD.n2582 0.714
R7772 VDD.n2564 VDD.n2563 0.714
R7773 VDD.n1128 VDD.n1127 0.714
R7774 VDD.n647 VDD.n646 0.714
R7775 VDD.n99 VDD.n96 0.714
R7776 VDD.n1704 VDD.n1701 0.714
R7777 VDD.n2060 VDD.n2059 0.714
R7778 VDD.n3007 VDD.n3006 0.708
R7779 VDD.n1496 VDD.n1493 0.708
R7780 VDD.n2430 VDD.n2427 0.708
R7781 VDD.n289 VDD.n288 0.702
R7782 VDD.n464 VDD.n461 0.702
R7783 VDD.n932 VDD.n929 0.702
R7784 VDD.n2805 VDD.n2804 0.702
R7785 VDD.n2762 VDD.n2761 0.702
R7786 VDD.n2227 VDD.n2224 0.702
R7787 VDD.n1404 VDD.n1403 0.702
R7788 VDD.n1805 VDD.n1804 0.702
R7789 VDD.n187 VDD.n182 0.624
R7790 VDD.n350 VDD.n345 0.624
R7791 VDD.n1909 VDD.n1904 0.624
R7792 VDD.n1746 VDD.n1741 0.624
R7793 VDD.n2350 VDD.n2347 0.624
R7794 VDD.n2350 VDD.n2349 0.624
R7795 VDD.n2476 VDD.n2473 0.624
R7796 VDD.n2476 VDD.n2475 0.624
R7797 VDD.n1140 VDD.n1139 0.619
R7798 VDD.n659 VDD.n658 0.619
R7799 VDD.n50 VDD.n47 0.619
R7800 VDD.n783 VDD.n780 0.619
R7801 VDD.n2072 VDD.n2071 0.619
R7802 VDD.n846 VDD.n843 0.616
R7803 VDD.n846 VDD.n845 0.616
R7804 VDD.n897 VDD.n894 0.616
R7805 VDD.n897 VDD.n896 0.616
R7806 VDD.n378 VDD.n375 0.616
R7807 VDD.n378 VDD.n377 0.616
R7808 VDD.n429 VDD.n426 0.616
R7809 VDD.n429 VDD.n428 0.616
R7810 VDD.n2701 VDD.n2696 0.616
R7811 VDD.n2869 VDD.n2863 0.616
R7812 VDD.n1302 VDD.n1297 0.616
R7813 VDD.n1464 VDD.n1459 0.616
R7814 VDD.n2133 VDD.n2130 0.616
R7815 VDD.n2133 VDD.n2132 0.616
R7816 VDD.n2196 VDD.n2193 0.616
R7817 VDD.n2196 VDD.n2195 0.616
R7818 VDD.n3111 VDD.n3106 0.616
R7819 VDD.n2948 VDD.n2943 0.616
R7820 VDD.n2995 VDD.n2994 0.614
R7821 VDD.n1270 VDD.n1267 0.614
R7822 VDD.n2390 VDD.n2389 0.614
R7823 VDD.n13 VDD.n10 0.609
R7824 VDD.n13 VDD.n12 0.609
R7825 VDD.n64 VDD.n61 0.609
R7826 VDD.n64 VDD.n63 0.609
R7827 VDD.n545 VDD.n540 0.609
R7828 VDD.n708 VDD.n703 0.609
R7829 VDD.n1026 VDD.n1021 0.609
R7830 VDD.n1189 VDD.n1184 0.609
R7831 VDD.n2515 VDD.n2512 0.609
R7832 VDD.n2515 VDD.n2514 0.609
R7833 VDD.n2631 VDD.n2628 0.609
R7834 VDD.n2631 VDD.n2630 0.609
R7835 VDD.n1958 VDD.n1953 0.609
R7836 VDD.n2120 VDD.n2115 0.609
R7837 VDD.n734 VDD.n731 0.609
R7838 VDD.n734 VDD.n733 0.609
R7839 VDD.n797 VDD.n794 0.609
R7840 VDD.n797 VDD.n796 0.609
R7841 VDD.n1221 VDD.n1218 0.609
R7842 VDD.n1221 VDD.n1220 0.609
R7843 VDD.n1284 VDD.n1281 0.609
R7844 VDD.n1284 VDD.n1283 0.609
R7845 VDD.n301 VDD.n300 0.608
R7846 VDD.n415 VDD.n412 0.608
R7847 VDD.n883 VDD.n880 0.608
R7848 VDD.n2182 VDD.n2179 0.608
R7849 VDD.n1416 VDD.n1415 0.608
R7850 VDD.n1793 VDD.n1792 0.608
R7851 VDD.n102 VDD.n101 0.575
R7852 VDD.n615 VDD.n614 0.575
R7853 VDD.n1096 VDD.n1095 0.575
R7854 VDD.n2566 VDD.n2565 0.575
R7855 VDD.n2640 VDD.n2639 0.575
R7856 VDD.n2567 VDD.n2566 0.575
R7857 VDD.n2639 VDD.n2638 0.575
R7858 VDD.n1095 VDD.n1094 0.575
R7859 VDD.n614 VDD.n613 0.575
R7860 VDD.n101 VDD.n100 0.575
R7861 VDD.n2028 VDD.n2027 0.575
R7862 VDD.n756 VDD.n755 0.575
R7863 VDD.n755 VDD.n754 0.575
R7864 VDD.n2027 VDD.n2026 0.575
R7865 VDD.n1243 VDD.n1242 0.57
R7866 VDD.n3035 VDD.n3034 0.57
R7867 VDD.n3034 VDD.n3033 0.57
R7868 VDD.n1242 VDD.n1241 0.57
R7869 VDD.n2413 VDD.n2412 0.57
R7870 VDD.n2412 VDD.n2411 0.57
R7871 VDD.n935 VDD.n934 0.565
R7872 VDD.n467 VDD.n466 0.565
R7873 VDD.n257 VDD.n256 0.565
R7874 VDD.n256 VDD.n255 0.565
R7875 VDD.n466 VDD.n465 0.565
R7876 VDD.n934 VDD.n933 0.565
R7877 VDD.n2772 VDD.n2771 0.565
R7878 VDD.n2792 VDD.n2791 0.565
R7879 VDD.n2773 VDD.n2772 0.565
R7880 VDD.n2791 VDD.n2790 0.565
R7881 VDD.n1833 VDD.n1832 0.565
R7882 VDD.n1372 VDD.n1371 0.565
R7883 VDD.n2155 VDD.n2154 0.565
R7884 VDD.n2154 VDD.n2153 0.565
R7885 VDD.n1371 VDD.n1370 0.565
R7886 VDD.n1832 VDD.n1831 0.565
R7887 VDD.n2604 VDD.n2601 0.522
R7888 VDD.n2545 VDD.n2544 0.522
R7889 VDD.n1152 VDD.n1151 0.522
R7890 VDD.n671 VDD.n670 0.522
R7891 VDD.n90 VDD.n87 0.522
R7892 VDD.n1695 VDD.n1692 0.522
R7893 VDD.n2084 VDD.n2083 0.522
R7894 VDD.n2983 VDD.n2982 0.517
R7895 VDD.n1487 VDD.n1484 0.517
R7896 VDD.n2449 VDD.n2446 0.517
R7897 VDD.n313 VDD.n312 0.512
R7898 VDD.n455 VDD.n452 0.512
R7899 VDD.n923 VDD.n920 0.512
R7900 VDD.n2830 VDD.n2829 0.512
R7901 VDD.n2737 VDD.n2736 0.512
R7902 VDD.n2218 VDD.n2215 0.512
R7903 VDD.n1428 VDD.n1427 0.512
R7904 VDD.n1781 VDD.n1780 0.512
R7905 VDD.n242 VDD.n241 0.468
R7906 VDD.n285 VDD.n284 0.468
R7907 VDD.n1844 VDD.n1843 0.468
R7908 VDD.n1801 VDD.n1800 0.468
R7909 VDD.n2395 VDD.n2394 0.468
R7910 VDD.n2397 VDD.n2396 0.468
R7911 VDD.n2423 VDD.n2422 0.468
R7912 VDD.n2425 VDD.n2424 0.468
R7913 VDD.n949 VDD.n948 0.462
R7914 VDD.n951 VDD.n950 0.462
R7915 VDD.n925 VDD.n924 0.462
R7916 VDD.n927 VDD.n926 0.462
R7917 VDD.n481 VDD.n480 0.462
R7918 VDD.n483 VDD.n482 0.462
R7919 VDD.n457 VDD.n456 0.462
R7920 VDD.n459 VDD.n458 0.462
R7921 VDD.n2758 VDD.n2757 0.462
R7922 VDD.n2801 VDD.n2800 0.462
R7923 VDD.n1357 VDD.n1356 0.462
R7924 VDD.n1400 VDD.n1399 0.462
R7925 VDD.n2232 VDD.n2231 0.462
R7926 VDD.n2234 VDD.n2233 0.462
R7927 VDD.n2220 VDD.n2219 0.462
R7928 VDD.n2222 VDD.n2221 0.462
R7929 VDD.n3046 VDD.n3045 0.462
R7930 VDD.n3003 VDD.n3002 0.462
R7931 VDD.n116 VDD.n115 0.457
R7932 VDD.n118 VDD.n117 0.457
R7933 VDD.n92 VDD.n91 0.457
R7934 VDD.n94 VDD.n93 0.457
R7935 VDD.n600 VDD.n599 0.457
R7936 VDD.n643 VDD.n642 0.457
R7937 VDD.n1081 VDD.n1080 0.457
R7938 VDD.n1124 VDD.n1123 0.457
R7939 VDD.n2559 VDD.n2558 0.457
R7940 VDD.n2561 VDD.n2560 0.457
R7941 VDD.n2578 VDD.n2577 0.457
R7942 VDD.n2580 VDD.n2579 0.457
R7943 VDD.n2013 VDD.n2012 0.457
R7944 VDD.n2056 VDD.n2055 0.457
R7945 VDD.n1709 VDD.n1708 0.457
R7946 VDD.n1711 VDD.n1710 0.457
R7947 VDD.n1697 VDD.n1696 0.457
R7948 VDD.n1699 VDD.n1698 0.457
R7949 VDD.n1501 VDD.n1500 0.457
R7950 VDD.n1503 VDD.n1502 0.457
R7951 VDD.n1489 VDD.n1488 0.457
R7952 VDD.n1491 VDD.n1490 0.457
R7953 VDD.n1164 VDD.n1163 0.422
R7954 VDD.n683 VDD.n682 0.422
R7955 VDD.n59 VDD.n56 0.422
R7956 VDD.n792 VDD.n789 0.422
R7957 VDD.n2096 VDD.n2095 0.422
R7958 VDD.n2971 VDD.n2970 0.418
R7959 VDD.n1279 VDD.n1276 0.418
R7960 VDD.n2371 VDD.n2370 0.418
R7961 VDD.n325 VDD.n324 0.415
R7962 VDD.n424 VDD.n421 0.415
R7963 VDD.n892 VDD.n889 0.415
R7964 VDD.n2191 VDD.n2188 0.415
R7965 VDD.n1440 VDD.n1439 0.415
R7966 VDD.n1769 VDD.n1768 0.415
R7967 VDD.n1918 VDD.n1917 0.38
R7968 VDD.n1291 VDD.n1207 0.38
R7969 VDD.n2885 VDD 0.38
R7970 VDD VDD.n3138 0.38
R7971 VDD VDD.n826 0.38
R7972 VDD.n1600 VDD 0.38
R7973 VDD.n1595 VDD.n1594 0.378
R7974 VDD.n818 VDD.n817 0.378
R7975 VDD.n359 VDD.n358 0.378
R7976 VDD.n2878 VDD.n2877 0.378
R7977 VDD.n2307 VDD.n2306 0.378
R7978 VDD.n2891 VDD.n2890 0.378
R7979 VDD.n2321 VDD.n2320 0.361
R7980 VDD.n1198 VDD.n1197 0.361
R7981 VDD.n1631 VDD.n1630 0.361
R7982 VDD.n1576 VDD.n1575 0.361
R7983 VDD.n3120 VDD.n3119 0.361
R7984 VDD.n717 VDD.n716 0.359
R7985 VDD.n2483 VDD.n2482 0.359
R7986 VDD.n1947 VDD.n1944 0.359
R7987 VDD.n2623 VDD.n2620 0.32
R7988 VDD.n2526 VDD.n2525 0.32
R7989 VDD.n1176 VDD.n1175 0.32
R7990 VDD.n695 VDD.n694 0.32
R7991 VDD.n81 VDD.n78 0.32
R7992 VDD.n1686 VDD.n1683 0.32
R7993 VDD.n2108 VDD.n2107 0.32
R7994 VDD.n2959 VDD.n2958 0.318
R7995 VDD.n1478 VDD.n1475 0.318
R7996 VDD.n2468 VDD.n2465 0.318
R7997 VDD.n337 VDD.n336 0.315
R7998 VDD.n446 VDD.n443 0.315
R7999 VDD.n914 VDD.n911 0.315
R8000 VDD.n2855 VDD.n2854 0.315
R8001 VDD.n2712 VDD.n2711 0.315
R8002 VDD.n2209 VDD.n2206 0.315
R8003 VDD.n1452 VDD.n1451 0.315
R8004 VDD.n1757 VDD.n1756 0.315
R8005 VDD.n2342 VDD.n2341 0.312
R8006 VDD.n904 VDD.n903 0.308
R8007 VDD.n436 VDD.n435 0.308
R8008 VDD.n2257 VDD.n2256 0.308
R8009 VDD.n71 VDD.n70 0.304
R8010 VDD.n2636 VDD.n2635 0.304
R8011 VDD.n1734 VDD.n1733 0.304
R8012 VDD.n1526 VDD.n1525 0.304
R8013 VDD.n1188 VDD.n1187 0.216
R8014 VDD.n707 VDD.n706 0.216
R8015 VDD.n68 VDD.n65 0.216
R8016 VDD.n801 VDD.n798 0.216
R8017 VDD.n2119 VDD.n2118 0.216
R8018 VDD.n2947 VDD.n2946 0.214
R8019 VDD.n1288 VDD.n1285 0.214
R8020 VDD.n2352 VDD.n2351 0.214
R8021 VDD.n349 VDD.n348 0.212
R8022 VDD.n433 VDD.n430 0.212
R8023 VDD.n901 VDD.n898 0.212
R8024 VDD.n2200 VDD.n2197 0.212
R8025 VDD.n1463 VDD.n1462 0.212
R8026 VDD.n1745 VDD.n1744 0.212
R8027 VDD.n254 VDD.n253 0.156
R8028 VDD.n273 VDD.n272 0.156
R8029 VDD.n1830 VDD.n1829 0.156
R8030 VDD.n1813 VDD.n1812 0.156
R8031 VDD.n2404 VDD.n2403 0.156
R8032 VDD.n2406 VDD.n2405 0.156
R8033 VDD.n2416 VDD.n2415 0.156
R8034 VDD.n2418 VDD.n2417 0.156
R8035 VDD.n937 VDD.n936 0.154
R8036 VDD.n940 VDD.n939 0.154
R8037 VDD.n867 VDD.n866 0.154
R8038 VDD.n869 VDD.n868 0.154
R8039 VDD.n469 VDD.n468 0.154
R8040 VDD.n472 VDD.n471 0.154
R8041 VDD.n399 VDD.n398 0.154
R8042 VDD.n401 VDD.n400 0.154
R8043 VDD.n2770 VDD.n2769 0.154
R8044 VDD.n2789 VDD.n2788 0.154
R8045 VDD.n1369 VDD.n1368 0.154
R8046 VDD.n1388 VDD.n1387 0.154
R8047 VDD.n2157 VDD.n2156 0.154
R8048 VDD.n2160 VDD.n2159 0.154
R8049 VDD.n2166 VDD.n2165 0.154
R8050 VDD.n2168 VDD.n2167 0.154
R8051 VDD.n3032 VDD.n3031 0.154
R8052 VDD.n3015 VDD.n3014 0.154
R8053 VDD.n104 VDD.n103 0.152
R8054 VDD.n107 VDD.n106 0.152
R8055 VDD.n34 VDD.n33 0.152
R8056 VDD.n36 VDD.n35 0.152
R8057 VDD.n612 VDD.n611 0.152
R8058 VDD.n631 VDD.n630 0.152
R8059 VDD.n1093 VDD.n1092 0.152
R8060 VDD.n1112 VDD.n1111 0.152
R8061 VDD.n2569 VDD.n2568 0.152
R8062 VDD.n2572 VDD.n2571 0.152
R8063 VDD.n2642 VDD.n2641 0.152
R8064 VDD.n2644 VDD.n2643 0.152
R8065 VDD.n2025 VDD.n2024 0.152
R8066 VDD.n2044 VDD.n2043 0.152
R8067 VDD.n758 VDD.n757 0.152
R8068 VDD.n761 VDD.n760 0.152
R8069 VDD.n767 VDD.n766 0.152
R8070 VDD.n769 VDD.n768 0.152
R8071 VDD.n1245 VDD.n1244 0.152
R8072 VDD.n1248 VDD.n1247 0.152
R8073 VDD.n1254 VDD.n1253 0.152
R8074 VDD.n1256 VDD.n1255 0.152
R8075 VDD.n154 VDD.n153 0.132
R8076 VDD.n627 VDD.n624 0.132
R8077 VDD.n1108 VDD.n1105 0.132
R8078 VDD.n993 VDD.n992 0.132
R8079 VDD.n512 VDD.n511 0.132
R8080 VDD.n269 VDD.n266 0.132
R8081 VDD.n2668 VDD.n2667 0.132
R8082 VDD.n2785 VDD.n2782 0.132
R8083 VDD.n1826 VDD.n1823 0.132
R8084 VDD.n1384 VDD.n1382 0.132
R8085 VDD.n2283 VDD.n2282 0.132
R8086 VDD.n2040 VDD.n2038 0.132
R8087 VDD.n1655 VDD.n1654 0.132
R8088 VDD.n1552 VDD.n1551 0.132
R8089 VDD.n3028 VDD.n3025 0.132
R8090 VDD.n2915 VDD.n2914 0.132
R8091 VDD.n1604 VDD.n1207 0.128
R8092 VDD.n2890 VDD.n2889 0.127
R8093 VDD.n2308 VDD.n2307 0.12
R8094 VDD.n1919 VDD.n1918 0.12
R8095 VDD.n2879 VDD.n2878 0.118
R8096 VDD.n819 VDD.n818 0.118
R8097 VDD.n360 VDD.n359 0.117
R8098 VDD.n1596 VDD.n1595 0.117
R8099 VDD.n172 VDD.n171 0.1
R8100 VDD.n169 VDD.n168 0.1
R8101 VDD.n166 VDD.n165 0.1
R8102 VDD.n163 VDD.n162 0.1
R8103 VDD.n160 VDD.n159 0.1
R8104 VDD.n157 VDD.n156 0.1
R8105 VDD.n151 VDD.n150 0.1
R8106 VDD.n148 VDD.n147 0.1
R8107 VDD.n145 VDD.n144 0.1
R8108 VDD.n142 VDD.n141 0.1
R8109 VDD.n2315 VDD.n2314 0.1
R8110 VDD.n2318 VDD.n2317 0.1
R8111 VDD.n558 VDD.n550 0.1
R8112 VDD.n570 VDD.n562 0.1
R8113 VDD.n582 VDD.n574 0.1
R8114 VDD.n594 VDD.n586 0.1
R8115 VDD.n606 VDD.n598 0.1
R8116 VDD.n620 VDD.n610 0.1
R8117 VDD.n639 VDD.n637 0.1
R8118 VDD.n651 VDD.n649 0.1
R8119 VDD.n663 VDD.n661 0.1
R8120 VDD.n675 VDD.n673 0.1
R8121 VDD.n687 VDD.n685 0.1
R8122 VDD.n699 VDD.n697 0.1
R8123 VDD.n711 VDD.n709 0.1
R8124 VDD.n1039 VDD.n1031 0.1
R8125 VDD.n1051 VDD.n1043 0.1
R8126 VDD.n1063 VDD.n1055 0.1
R8127 VDD.n1075 VDD.n1067 0.1
R8128 VDD.n1087 VDD.n1079 0.1
R8129 VDD.n1101 VDD.n1091 0.1
R8130 VDD.n1120 VDD.n1118 0.1
R8131 VDD.n1132 VDD.n1130 0.1
R8132 VDD.n1144 VDD.n1142 0.1
R8133 VDD.n1156 VDD.n1154 0.1
R8134 VDD.n1168 VDD.n1166 0.1
R8135 VDD.n1180 VDD.n1178 0.1
R8136 VDD.n1192 VDD.n1190 0.1
R8137 VDD.n1011 VDD.n1010 0.1
R8138 VDD.n1008 VDD.n1007 0.1
R8139 VDD.n1005 VDD.n1004 0.1
R8140 VDD.n1002 VDD.n1001 0.1
R8141 VDD.n999 VDD.n998 0.1
R8142 VDD.n996 VDD.n995 0.1
R8143 VDD.n990 VDD.n989 0.1
R8144 VDD.n987 VDD.n986 0.1
R8145 VDD.n984 VDD.n983 0.1
R8146 VDD.n981 VDD.n980 0.1
R8147 VDD.n978 VDD.n977 0.1
R8148 VDD.n975 VDD.n974 0.1
R8149 VDD.n530 VDD.n529 0.1
R8150 VDD.n527 VDD.n526 0.1
R8151 VDD.n524 VDD.n523 0.1
R8152 VDD.n521 VDD.n520 0.1
R8153 VDD.n518 VDD.n517 0.1
R8154 VDD.n515 VDD.n514 0.1
R8155 VDD.n509 VDD.n508 0.1
R8156 VDD.n506 VDD.n505 0.1
R8157 VDD.n803 VDD.n802 0.1
R8158 VDD.n806 VDD.n805 0.1
R8159 VDD.n809 VDD.n808 0.1
R8160 VDD.n812 VDD.n811 0.1
R8161 VDD.n815 VDD.n814 0.1
R8162 VDD.n200 VDD.n192 0.1
R8163 VDD.n212 VDD.n204 0.1
R8164 VDD.n224 VDD.n216 0.1
R8165 VDD.n236 VDD.n228 0.1
R8166 VDD.n248 VDD.n240 0.1
R8167 VDD.n262 VDD.n252 0.1
R8168 VDD.n281 VDD.n279 0.1
R8169 VDD.n293 VDD.n291 0.1
R8170 VDD.n305 VDD.n303 0.1
R8171 VDD.n317 VDD.n315 0.1
R8172 VDD.n329 VDD.n327 0.1
R8173 VDD.n341 VDD.n339 0.1
R8174 VDD.n353 VDD.n351 0.1
R8175 VDD.n2686 VDD.n2685 0.1
R8176 VDD.n2683 VDD.n2682 0.1
R8177 VDD.n2680 VDD.n2679 0.1
R8178 VDD.n2677 VDD.n2676 0.1
R8179 VDD.n2674 VDD.n2673 0.1
R8180 VDD.n2671 VDD.n2670 0.1
R8181 VDD.n2665 VDD.n2664 0.1
R8182 VDD.n2662 VDD.n2661 0.1
R8183 VDD.n2659 VDD.n2658 0.1
R8184 VDD.n2656 VDD.n2655 0.1
R8185 VDD.n2653 VDD.n2652 0.1
R8186 VDD.n2650 VDD.n2649 0.1
R8187 VDD.n2714 VDD.n2706 0.1
R8188 VDD.n2727 VDD.n2718 0.1
R8189 VDD.n2739 VDD.n2731 0.1
R8190 VDD.n2752 VDD.n2743 0.1
R8191 VDD.n2764 VDD.n2756 0.1
R8192 VDD.n2778 VDD.n2768 0.1
R8193 VDD.n2797 VDD.n2795 0.1
R8194 VDD.n2809 VDD.n2807 0.1
R8195 VDD.n2822 VDD.n2820 0.1
R8196 VDD.n2834 VDD.n2832 0.1
R8197 VDD.n2847 VDD.n2845 0.1
R8198 VDD.n2859 VDD.n2857 0.1
R8199 VDD.n2872 VDD.n2870 0.1
R8200 VDD.n1912 VDD.n1910 0.1
R8201 VDD.n1900 VDD.n1898 0.1
R8202 VDD.n1888 VDD.n1886 0.1
R8203 VDD.n1876 VDD.n1874 0.1
R8204 VDD.n1864 VDD.n1862 0.1
R8205 VDD.n1852 VDD.n1850 0.1
R8206 VDD.n1840 VDD.n1838 0.1
R8207 VDD.n1819 VDD.n1811 0.1
R8208 VDD.n1807 VDD.n1799 0.1
R8209 VDD.n1795 VDD.n1787 0.1
R8210 VDD.n1783 VDD.n1775 0.1
R8211 VDD.n1771 VDD.n1763 0.1
R8212 VDD.n1759 VDD.n1751 0.1
R8213 VDD.n1303 VDD.n1295 0.1
R8214 VDD.n1315 VDD.n1307 0.1
R8215 VDD.n1327 VDD.n1319 0.1
R8216 VDD.n1339 VDD.n1331 0.1
R8217 VDD.n1351 VDD.n1343 0.1
R8218 VDD.n1363 VDD.n1355 0.1
R8219 VDD.n1377 VDD.n1367 0.1
R8220 VDD.n1396 VDD.n1394 0.1
R8221 VDD.n1408 VDD.n1406 0.1
R8222 VDD.n1420 VDD.n1418 0.1
R8223 VDD.n1432 VDD.n1430 0.1
R8224 VDD.n1444 VDD.n1442 0.1
R8225 VDD.n1456 VDD.n1454 0.1
R8226 VDD.n2304 VDD.n2303 0.1
R8227 VDD.n2301 VDD.n2300 0.1
R8228 VDD.n2298 VDD.n2297 0.1
R8229 VDD.n2295 VDD.n2294 0.1
R8230 VDD.n2292 VDD.n2291 0.1
R8231 VDD.n2289 VDD.n2288 0.1
R8232 VDD.n2286 VDD.n2285 0.1
R8233 VDD.n2280 VDD.n2279 0.1
R8234 VDD.n2277 VDD.n2276 0.1
R8235 VDD.n2274 VDD.n2273 0.1
R8236 VDD.n2271 VDD.n2270 0.1
R8237 VDD.n2268 VDD.n2267 0.1
R8238 VDD.n2265 VDD.n2264 0.1
R8239 VDD.n1959 VDD.n1951 0.1
R8240 VDD.n1971 VDD.n1963 0.1
R8241 VDD.n1983 VDD.n1975 0.1
R8242 VDD.n1995 VDD.n1987 0.1
R8243 VDD.n2007 VDD.n1999 0.1
R8244 VDD.n2019 VDD.n2011 0.1
R8245 VDD.n2033 VDD.n2023 0.1
R8246 VDD.n2052 VDD.n2050 0.1
R8247 VDD.n2064 VDD.n2062 0.1
R8248 VDD.n2076 VDD.n2074 0.1
R8249 VDD.n2088 VDD.n2086 0.1
R8250 VDD.n2100 VDD.n2098 0.1
R8251 VDD.n2112 VDD.n2110 0.1
R8252 VDD.n1634 VDD.n1633 0.1
R8253 VDD.n1637 VDD.n1636 0.1
R8254 VDD.n1640 VDD.n1639 0.1
R8255 VDD.n1643 VDD.n1642 0.1
R8256 VDD.n1646 VDD.n1645 0.1
R8257 VDD.n1649 VDD.n1648 0.1
R8258 VDD.n1652 VDD.n1651 0.1
R8259 VDD.n1658 VDD.n1657 0.1
R8260 VDD.n1661 VDD.n1660 0.1
R8261 VDD.n1664 VDD.n1663 0.1
R8262 VDD.n1667 VDD.n1666 0.1
R8263 VDD.n1670 VDD.n1669 0.1
R8264 VDD.n1673 VDD.n1672 0.1
R8265 VDD.n1573 VDD.n1572 0.1
R8266 VDD.n1570 VDD.n1569 0.1
R8267 VDD.n1567 VDD.n1566 0.1
R8268 VDD.n1564 VDD.n1563 0.1
R8269 VDD.n1561 VDD.n1560 0.1
R8270 VDD.n1558 VDD.n1557 0.1
R8271 VDD.n1555 VDD.n1554 0.1
R8272 VDD.n1549 VDD.n1548 0.1
R8273 VDD.n1546 VDD.n1545 0.1
R8274 VDD.n1543 VDD.n1542 0.1
R8275 VDD.n1540 VDD.n1539 0.1
R8276 VDD.n1537 VDD.n1536 0.1
R8277 VDD.n1534 VDD.n1533 0.1
R8278 VDD.n3114 VDD.n3112 0.1
R8279 VDD.n3102 VDD.n3100 0.1
R8280 VDD.n3090 VDD.n3088 0.1
R8281 VDD.n3078 VDD.n3076 0.1
R8282 VDD.n3066 VDD.n3064 0.1
R8283 VDD.n3054 VDD.n3052 0.1
R8284 VDD.n3042 VDD.n3040 0.1
R8285 VDD.n3021 VDD.n3013 0.1
R8286 VDD.n3009 VDD.n3001 0.1
R8287 VDD.n2997 VDD.n2989 0.1
R8288 VDD.n2985 VDD.n2977 0.1
R8289 VDD.n2973 VDD.n2965 0.1
R8290 VDD.n2961 VDD.n2953 0.1
R8291 VDD.n2894 VDD.n2893 0.1
R8292 VDD.n2897 VDD.n2896 0.1
R8293 VDD.n2900 VDD.n2899 0.1
R8294 VDD.n2903 VDD.n2902 0.1
R8295 VDD.n2906 VDD.n2905 0.1
R8296 VDD.n2909 VDD.n2908 0.1
R8297 VDD.n2912 VDD.n2911 0.1
R8298 VDD.n2918 VDD.n2917 0.1
R8299 VDD.n2921 VDD.n2920 0.1
R8300 VDD.n2924 VDD.n2923 0.1
R8301 VDD.n2927 VDD.n2926 0.1
R8302 VDD.n2930 VDD.n2929 0.1
R8303 VDD.n2933 VDD.n2932 0.1
R8304 VDD.n2494 VDD.n2493 0.075
R8305 VDD.n1213 VDD.n1211 0.072
R8306 VDD.n1931 VDD.n370 0.064
R8307 VDD.n1617 VDD.n838 0.064
R8308 VDD.n3127 VDD.n2331 0.064
R8309 VDD.n3126 VDD.n2332 0.061
R8310 VDD.n1618 VDD.n837 0.061
R8311 VDD.n1932 VDD.n369 0.061
R8312 VDD.n722 VDD.n721 0.06
R8313 VDD.n2488 VDD.n2487 0.06
R8314 VDD.n1581 VDD.n1580 0.06
R8315 VDD.n2326 VDD.n2325 0.059
R8316 VDD.n1203 VDD.n1202 0.059
R8317 VDD.n1936 VDD.n1935 0.059
R8318 VDD.n1622 VDD.n1621 0.059
R8319 VDD.n2337 VDD.n2336 0.059
R8320 VDD.n2322 VDD.n2321 0.058
R8321 VDD.n718 VDD.n717 0.058
R8322 VDD.n1199 VDD.n1198 0.058
R8323 VDD.n2484 VDD.n2483 0.058
R8324 VDD.n1944 VDD.n1943 0.058
R8325 VDD.n1630 VDD.n1629 0.058
R8326 VDD.n1577 VDD.n1576 0.058
R8327 VDD.n3121 VDD.n3120 0.058
R8328 VDD.n2328 VDD.n2327 0.051
R8329 VDD.n1624 VDD.n1623 0.051
R8330 VDD.n1583 VDD.n1582 0.051
R8331 VDD.n2339 VDD.n2338 0.051
R8332 VDD.n724 VDD.n723 0.05
R8333 VDD.n1205 VDD.n1204 0.05
R8334 VDD.n2490 VDD.n2489 0.05
R8335 VDD.n1938 VDD.n1937 0.05
R8336 VDD.n2327 VDD.n2326 0.043
R8337 VDD.n723 VDD.n722 0.043
R8338 VDD.n1204 VDD.n1203 0.043
R8339 VDD.n2489 VDD.n2488 0.043
R8340 VDD.n1937 VDD.n1936 0.043
R8341 VDD.n1623 VDD.n1622 0.043
R8342 VDD.n1582 VDD.n1581 0.043
R8343 VDD.n2338 VDD.n2337 0.043
R8344 VDD.n2324 VDD.n2323 0.039
R8345 VDD.n2323 VDD.n2322 0.039
R8346 VDD.n720 VDD.n719 0.039
R8347 VDD.n719 VDD.n718 0.039
R8348 VDD.n1201 VDD.n1200 0.039
R8349 VDD.n1200 VDD.n1199 0.039
R8350 VDD.n2486 VDD.n2485 0.039
R8351 VDD.n2485 VDD.n2484 0.039
R8352 VDD.n1943 VDD.n1942 0.039
R8353 VDD.n1942 VDD.n1941 0.039
R8354 VDD.n1629 VDD.n1628 0.039
R8355 VDD.n1628 VDD.n1627 0.039
R8356 VDD.n1578 VDD.n1577 0.039
R8357 VDD.n1579 VDD.n1578 0.039
R8358 VDD.n3122 VDD.n3121 0.039
R8359 VDD.n3123 VDD.n3122 0.039
R8360 VDD.n3129 VDD.n2324 0.03
R8361 VDD.n156 VDD.n155 0.03
R8362 VDD.n152 VDD.n151 0.03
R8363 VDD.n1928 VDD.n720 0.03
R8364 VDD.n622 VDD.n620 0.03
R8365 VDD.n637 VDD.n629 0.03
R8366 VDD.n1206 VDD.n1201 0.03
R8367 VDD.n1103 VDD.n1101 0.03
R8368 VDD.n1118 VDD.n1110 0.03
R8369 VDD.n995 VDD.n994 0.03
R8370 VDD.n991 VDD.n990 0.03
R8371 VDD.n514 VDD.n513 0.03
R8372 VDD.n510 VDD.n509 0.03
R8373 VDD.n264 VDD.n262 0.03
R8374 VDD.n279 VDD.n271 0.03
R8375 VDD.n2495 VDD.n2486 0.03
R8376 VDD.n2670 VDD.n2669 0.03
R8377 VDD.n2666 VDD.n2665 0.03
R8378 VDD.n2780 VDD.n2778 0.03
R8379 VDD.n2795 VDD.n2787 0.03
R8380 VDD.n1838 VDD.n1828 0.03
R8381 VDD.n1821 VDD.n1819 0.03
R8382 VDD.n1379 VDD.n1377 0.03
R8383 VDD.n1394 VDD.n1386 0.03
R8384 VDD.n2285 VDD.n2284 0.03
R8385 VDD.n2281 VDD.n2280 0.03
R8386 VDD.n1941 VDD.n1940 0.03
R8387 VDD.n2035 VDD.n2033 0.03
R8388 VDD.n2050 VDD.n2042 0.03
R8389 VDD.n1627 VDD.n1626 0.03
R8390 VDD.n1653 VDD.n1652 0.03
R8391 VDD.n1657 VDD.n1656 0.03
R8392 VDD.n1585 VDD.n1579 0.03
R8393 VDD.n1554 VDD.n1553 0.03
R8394 VDD.n1550 VDD.n1549 0.03
R8395 VDD.n3124 VDD.n3123 0.03
R8396 VDD.n3040 VDD.n3030 0.03
R8397 VDD.n3023 VDD.n3021 0.03
R8398 VDD.n2913 VDD.n2912 0.03
R8399 VDD.n2917 VDD.n2916 0.03
R8400 VDD.n2319 VDD.n2318 0.028
R8401 VDD.n713 VDD.n711 0.028
R8402 VDD.n1194 VDD.n1192 0.028
R8403 VDD.n1593 VDD.n1592 0.028
R8404 VDD.n816 VDD.n815 0.028
R8405 VDD.n355 VDD.n353 0.028
R8406 VDD.n2481 VDD.n2480 0.028
R8407 VDD.n2874 VDD.n2872 0.028
R8408 VDD.n1914 VDD.n1912 0.028
R8409 VDD.n1295 VDD.n1293 0.028
R8410 VDD.n2305 VDD.n2304 0.028
R8411 VDD.n1951 VDD.n1949 0.028
R8412 VDD.n1633 VDD.n1632 0.028
R8413 VDD.n1574 VDD.n1573 0.028
R8414 VDD.n3116 VDD.n3114 0.028
R8415 VDD.n2893 VDD.n2892 0.028
R8416 VDD.n159 VDD.n158 0.026
R8417 VDD.n149 VDD.n148 0.026
R8418 VDD.n608 VDD.n606 0.026
R8419 VDD.n649 VDD.n641 0.026
R8420 VDD.n1089 VDD.n1087 0.026
R8421 VDD.n1130 VDD.n1122 0.026
R8422 VDD.n998 VDD.n997 0.026
R8423 VDD.n988 VDD.n987 0.026
R8424 VDD.n517 VDD.n516 0.026
R8425 VDD.n507 VDD.n506 0.026
R8426 VDD.n250 VDD.n248 0.026
R8427 VDD.n291 VDD.n283 0.026
R8428 VDD.n2673 VDD.n2672 0.026
R8429 VDD.n2663 VDD.n2662 0.026
R8430 VDD.n2766 VDD.n2764 0.026
R8431 VDD.n2807 VDD.n2799 0.026
R8432 VDD.n1850 VDD.n1842 0.026
R8433 VDD.n1809 VDD.n1807 0.026
R8434 VDD.n1365 VDD.n1363 0.026
R8435 VDD.n1406 VDD.n1398 0.026
R8436 VDD.n2288 VDD.n2287 0.026
R8437 VDD.n2278 VDD.n2277 0.026
R8438 VDD.n2021 VDD.n2019 0.026
R8439 VDD.n2062 VDD.n2054 0.026
R8440 VDD.n1650 VDD.n1649 0.026
R8441 VDD.n1660 VDD.n1659 0.026
R8442 VDD.n1557 VDD.n1556 0.026
R8443 VDD.n1547 VDD.n1546 0.026
R8444 VDD.n3052 VDD.n3044 0.026
R8445 VDD.n3011 VDD.n3009 0.026
R8446 VDD.n2910 VDD.n2909 0.026
R8447 VDD.n2920 VDD.n2919 0.026
R8448 VDD.n173 VDD.n172 0.024
R8449 VDD.n2316 VDD.n2315 0.024
R8450 VDD.n550 VDD.n548 0.024
R8451 VDD.n701 VDD.n699 0.024
R8452 VDD.n1031 VDD.n1029 0.024
R8453 VDD.n1182 VDD.n1180 0.024
R8454 VDD.n1012 VDD.n1011 0.024
R8455 VDD.n974 VDD.n973 0.024
R8456 VDD.n531 VDD.n530 0.024
R8457 VDD.n813 VDD.n812 0.024
R8458 VDD.n192 VDD.n190 0.024
R8459 VDD.n343 VDD.n341 0.024
R8460 VDD.n2687 VDD.n2686 0.024
R8461 VDD.n2649 VDD.n2648 0.024
R8462 VDD.n2706 VDD.n2704 0.024
R8463 VDD.n2861 VDD.n2859 0.024
R8464 VDD.n1902 VDD.n1900 0.024
R8465 VDD.n1751 VDD.n1749 0.024
R8466 VDD.n1307 VDD.n1305 0.024
R8467 VDD.n1458 VDD.n1456 0.024
R8468 VDD.n2302 VDD.n2301 0.024
R8469 VDD.n2264 VDD.n2263 0.024
R8470 VDD.n1963 VDD.n1961 0.024
R8471 VDD.n2114 VDD.n2112 0.024
R8472 VDD.n1636 VDD.n1635 0.024
R8473 VDD.n1674 VDD.n1673 0.024
R8474 VDD.n1571 VDD.n1570 0.024
R8475 VDD.n1533 VDD.n1532 0.024
R8476 VDD.n3104 VDD.n3102 0.024
R8477 VDD.n2953 VDD.n2951 0.024
R8478 VDD.n2896 VDD.n2895 0.024
R8479 VDD.n2934 VDD.n2933 0.024
R8480 VDD.n162 VDD.n161 0.022
R8481 VDD.n146 VDD.n145 0.022
R8482 VDD.n596 VDD.n594 0.022
R8483 VDD.n661 VDD.n653 0.022
R8484 VDD.n1077 VDD.n1075 0.022
R8485 VDD.n1142 VDD.n1134 0.022
R8486 VDD.n1001 VDD.n1000 0.022
R8487 VDD.n985 VDD.n984 0.022
R8488 VDD.n520 VDD.n519 0.022
R8489 VDD.n238 VDD.n236 0.022
R8490 VDD.n303 VDD.n295 0.022
R8491 VDD.n2676 VDD.n2675 0.022
R8492 VDD.n2660 VDD.n2659 0.022
R8493 VDD.n2754 VDD.n2752 0.022
R8494 VDD.n2820 VDD.n2811 0.022
R8495 VDD.n1862 VDD.n1854 0.022
R8496 VDD.n1797 VDD.n1795 0.022
R8497 VDD.n1353 VDD.n1351 0.022
R8498 VDD.n1418 VDD.n1410 0.022
R8499 VDD.n2291 VDD.n2290 0.022
R8500 VDD.n2275 VDD.n2274 0.022
R8501 VDD.n2009 VDD.n2007 0.022
R8502 VDD.n2074 VDD.n2066 0.022
R8503 VDD.n1647 VDD.n1646 0.022
R8504 VDD.n1663 VDD.n1662 0.022
R8505 VDD.n1560 VDD.n1559 0.022
R8506 VDD.n1544 VDD.n1543 0.022
R8507 VDD.n3064 VDD.n3056 0.022
R8508 VDD.n2999 VDD.n2997 0.022
R8509 VDD.n2907 VDD.n2906 0.022
R8510 VDD.n2923 VDD.n2922 0.022
R8511 VDD.n170 VDD.n169 0.02
R8512 VDD.n2313 VDD.n2312 0.02
R8513 VDD.n562 VDD.n560 0.02
R8514 VDD.n689 VDD.n687 0.02
R8515 VDD.n1043 VDD.n1041 0.02
R8516 VDD.n1170 VDD.n1168 0.02
R8517 VDD.n1009 VDD.n1008 0.02
R8518 VDD.n977 VDD.n976 0.02
R8519 VDD.n528 VDD.n527 0.02
R8520 VDD.n810 VDD.n809 0.02
R8521 VDD.n204 VDD.n202 0.02
R8522 VDD.n331 VDD.n329 0.02
R8523 VDD.n2684 VDD.n2683 0.02
R8524 VDD.n2652 VDD.n2651 0.02
R8525 VDD.n2718 VDD.n2716 0.02
R8526 VDD.n2849 VDD.n2847 0.02
R8527 VDD.n1890 VDD.n1888 0.02
R8528 VDD.n1763 VDD.n1761 0.02
R8529 VDD.n1319 VDD.n1317 0.02
R8530 VDD.n1446 VDD.n1444 0.02
R8531 VDD.n2299 VDD.n2298 0.02
R8532 VDD.n2267 VDD.n2266 0.02
R8533 VDD.n1975 VDD.n1973 0.02
R8534 VDD.n2102 VDD.n2100 0.02
R8535 VDD.n1639 VDD.n1638 0.02
R8536 VDD.n1671 VDD.n1670 0.02
R8537 VDD.n1568 VDD.n1567 0.02
R8538 VDD.n1536 VDD.n1535 0.02
R8539 VDD.n3092 VDD.n3090 0.02
R8540 VDD.n2965 VDD.n2963 0.02
R8541 VDD.n2899 VDD.n2898 0.02
R8542 VDD.n2931 VDD.n2930 0.02
R8543 VDD.n165 VDD.n164 0.018
R8544 VDD.n143 VDD.n142 0.018
R8545 VDD.n584 VDD.n582 0.018
R8546 VDD.n673 VDD.n665 0.018
R8547 VDD.n1065 VDD.n1063 0.018
R8548 VDD.n1154 VDD.n1146 0.018
R8549 VDD.n1004 VDD.n1003 0.018
R8550 VDD.n982 VDD.n981 0.018
R8551 VDD.n523 VDD.n522 0.018
R8552 VDD.n805 VDD.n804 0.018
R8553 VDD.n226 VDD.n224 0.018
R8554 VDD.n315 VDD.n307 0.018
R8555 VDD.n2679 VDD.n2678 0.018
R8556 VDD.n2657 VDD.n2656 0.018
R8557 VDD.n2741 VDD.n2739 0.018
R8558 VDD.n2832 VDD.n2824 0.018
R8559 VDD.n1874 VDD.n1866 0.018
R8560 VDD.n1785 VDD.n1783 0.018
R8561 VDD.n1341 VDD.n1339 0.018
R8562 VDD.n1430 VDD.n1422 0.018
R8563 VDD.n2294 VDD.n2293 0.018
R8564 VDD.n2272 VDD.n2271 0.018
R8565 VDD.n1997 VDD.n1995 0.018
R8566 VDD.n2086 VDD.n2078 0.018
R8567 VDD.n1644 VDD.n1643 0.018
R8568 VDD.n1666 VDD.n1665 0.018
R8569 VDD.n1563 VDD.n1562 0.018
R8570 VDD.n1541 VDD.n1540 0.018
R8571 VDD.n3076 VDD.n3068 0.018
R8572 VDD.n2987 VDD.n2985 0.018
R8573 VDD.n2904 VDD.n2903 0.018
R8574 VDD.n2926 VDD.n2925 0.018
R8575 VDD.n167 VDD.n166 0.017
R8576 VDD.n141 VDD.n140 0.017
R8577 VDD.n574 VDD.n572 0.017
R8578 VDD.n677 VDD.n675 0.017
R8579 VDD.n1055 VDD.n1053 0.017
R8580 VDD.n1158 VDD.n1156 0.017
R8581 VDD.n1006 VDD.n1005 0.017
R8582 VDD.n980 VDD.n979 0.017
R8583 VDD.n525 VDD.n524 0.017
R8584 VDD.n807 VDD.n806 0.017
R8585 VDD.n216 VDD.n214 0.017
R8586 VDD.n319 VDD.n317 0.017
R8587 VDD.n2681 VDD.n2680 0.017
R8588 VDD.n2655 VDD.n2654 0.017
R8589 VDD.n2731 VDD.n2729 0.017
R8590 VDD.n2836 VDD.n2834 0.017
R8591 VDD.n1878 VDD.n1876 0.017
R8592 VDD.n1775 VDD.n1773 0.017
R8593 VDD.n1331 VDD.n1329 0.017
R8594 VDD.n1434 VDD.n1432 0.017
R8595 VDD.n2296 VDD.n2295 0.017
R8596 VDD.n2270 VDD.n2269 0.017
R8597 VDD.n1987 VDD.n1985 0.017
R8598 VDD.n2090 VDD.n2088 0.017
R8599 VDD.n1642 VDD.n1641 0.017
R8600 VDD.n1668 VDD.n1667 0.017
R8601 VDD.n1565 VDD.n1564 0.017
R8602 VDD.n1539 VDD.n1538 0.017
R8603 VDD.n3080 VDD.n3078 0.017
R8604 VDD.n2977 VDD.n2975 0.017
R8605 VDD.n2902 VDD.n2901 0.017
R8606 VDD.n2928 VDD.n2927 0.017
R8607 VDD.n1618 VDD.n1617 0.017
R8608 VDD.n1932 VDD.n1931 0.017
R8609 VDD.n3129 VDD.n2328 0.016
R8610 VDD.n1928 VDD.n724 0.016
R8611 VDD.n1206 VDD.n1205 0.016
R8612 VDD.n2495 VDD.n2490 0.016
R8613 VDD.n1940 VDD.n1938 0.016
R8614 VDD.n1626 VDD.n1624 0.016
R8615 VDD.n1585 VDD.n1583 0.016
R8616 VDD.n3124 VDD.n2339 0.016
R8617 VDD.n1603 VDD.n1602 0.015
R8618 VDD.n2888 VDD.n2887 0.015
R8619 VDD.n168 VDD.n167 0.015
R8620 VDD.n140 VDD.n139 0.015
R8621 VDD.n572 VDD.n570 0.015
R8622 VDD.n685 VDD.n677 0.015
R8623 VDD.n1053 VDD.n1051 0.015
R8624 VDD.n1166 VDD.n1158 0.015
R8625 VDD.n1007 VDD.n1006 0.015
R8626 VDD.n979 VDD.n978 0.015
R8627 VDD.n526 VDD.n525 0.015
R8628 VDD.n808 VDD.n807 0.015
R8629 VDD.n214 VDD.n212 0.015
R8630 VDD.n327 VDD.n319 0.015
R8631 VDD.n2682 VDD.n2681 0.015
R8632 VDD.n2654 VDD.n2653 0.015
R8633 VDD.n2729 VDD.n2727 0.015
R8634 VDD.n2845 VDD.n2836 0.015
R8635 VDD.n1886 VDD.n1878 0.015
R8636 VDD.n1773 VDD.n1771 0.015
R8637 VDD.n1329 VDD.n1327 0.015
R8638 VDD.n1442 VDD.n1434 0.015
R8639 VDD.n2297 VDD.n2296 0.015
R8640 VDD.n2269 VDD.n2268 0.015
R8641 VDD.n1985 VDD.n1983 0.015
R8642 VDD.n2098 VDD.n2090 0.015
R8643 VDD.n1641 VDD.n1640 0.015
R8644 VDD.n1669 VDD.n1668 0.015
R8645 VDD.n1566 VDD.n1565 0.015
R8646 VDD.n1538 VDD.n1537 0.015
R8647 VDD.n3088 VDD.n3080 0.015
R8648 VDD.n2975 VDD.n2973 0.015
R8649 VDD.n2901 VDD.n2900 0.015
R8650 VDD.n2929 VDD.n2928 0.015
R8651 VDD.n3127 VDD.n3126 0.015
R8652 VDD.n1923 VDD.n1921 0.015
R8653 VDD.n2501 VDD.n2500 0.015
R8654 VDD.n3134 VDD.n3133 0.014
R8655 VDD.n1607 VDD.n1605 0.014
R8656 VDD.n834 VDD.n833 0.014
R8657 VDD.n1210 VDD.n1209 0.014
R8658 VDD.n826 VDD.n825 0.014
R8659 VDD.n366 VDD.n365 0.014
R8660 VDD.n3138 VDD.n3137 0.014
R8661 VDD.n1 VDD.n0 0.014
R8662 VDD.n1920 VDD.n1919 0.014
R8663 VDD.n2504 VDD.n2503 0.014
R8664 VDD.n2881 VDD.n2507 0.013
R8665 VDD.n363 VDD.n362 0.013
R8666 VDD.n831 VDD.n830 0.013
R8667 VDD.n164 VDD.n163 0.013
R8668 VDD.n144 VDD.n143 0.013
R8669 VDD.n586 VDD.n584 0.013
R8670 VDD.n665 VDD.n663 0.013
R8671 VDD.n1067 VDD.n1065 0.013
R8672 VDD.n1146 VDD.n1144 0.013
R8673 VDD.n1003 VDD.n1002 0.013
R8674 VDD.n983 VDD.n982 0.013
R8675 VDD.n522 VDD.n521 0.013
R8676 VDD.n804 VDD.n803 0.013
R8677 VDD.n228 VDD.n226 0.013
R8678 VDD.n307 VDD.n305 0.013
R8679 VDD.n2678 VDD.n2677 0.013
R8680 VDD.n2658 VDD.n2657 0.013
R8681 VDD.n2743 VDD.n2741 0.013
R8682 VDD.n2824 VDD.n2822 0.013
R8683 VDD.n1866 VDD.n1864 0.013
R8684 VDD.n1787 VDD.n1785 0.013
R8685 VDD.n1343 VDD.n1341 0.013
R8686 VDD.n1422 VDD.n1420 0.013
R8687 VDD.n2293 VDD.n2292 0.013
R8688 VDD.n2273 VDD.n2272 0.013
R8689 VDD.n1999 VDD.n1997 0.013
R8690 VDD.n2078 VDD.n2076 0.013
R8691 VDD.n1645 VDD.n1644 0.013
R8692 VDD.n1665 VDD.n1664 0.013
R8693 VDD.n1562 VDD.n1561 0.013
R8694 VDD.n1542 VDD.n1541 0.013
R8695 VDD.n3068 VDD.n3066 0.013
R8696 VDD.n2989 VDD.n2987 0.013
R8697 VDD.n2905 VDD.n2904 0.013
R8698 VDD.n2925 VDD.n2924 0.013
R8699 VDD.n1612 VDD.n1610 0.013
R8700 VDD.n820 VDD.n819 0.013
R8701 VDD.n2311 VDD.n2310 0.013
R8702 VDD.n2334 VDD.n2333 0.013
R8703 VDD.n2880 VDD.n2879 0.013
R8704 VDD.n2309 VDD.n2308 0.013
R8705 VDD.n1591 VDD.n1589 0.012
R8706 VDD.n1587 VDD.n1586 0.012
R8707 VDD.n836 VDD.n835 0.012
R8708 VDD.n368 VDD.n367 0.012
R8709 VDD.n2505 VDD.n2335 0.012
R8710 VDD.n1620 VDD.n1618 0.012
R8711 VDD.n1934 VDD.n1932 0.012
R8712 VDD.n3126 VDD.n3125 0.012
R8713 VDD.n3129 VDD.n2329 0.012
R8714 VDD.n1928 VDD.n725 0.012
R8715 VDD.n1925 VDD.n1924 0.012
R8716 VDD.n1609 VDD.n1608 0.012
R8717 VDD.n1614 VDD.n1613 0.012
R8718 VDD.n828 VDD.n821 0.012
R8719 VDD.n2499 VDD.n2498 0.012
R8720 VDD.n2495 VDD.n2491 0.012
R8721 VDD.n1626 VDD.n1625 0.012
R8722 VDD.n1585 VDD.n1584 0.012
R8723 VDD.n1597 VDD.n1596 0.012
R8724 VDD.n1940 VDD.n1939 0.012
R8725 VDD.n361 VDD.n360 0.012
R8726 VDD.n3128 VDD.n3127 0.011
R8727 VDD.n1931 VDD.n1930 0.011
R8728 VDD.n171 VDD.n170 0.011
R8729 VDD.n2314 VDD.n2313 0.011
R8730 VDD.n560 VDD.n558 0.011
R8731 VDD.n697 VDD.n689 0.011
R8732 VDD.n1041 VDD.n1039 0.011
R8733 VDD.n1178 VDD.n1170 0.011
R8734 VDD.n1010 VDD.n1009 0.011
R8735 VDD.n976 VDD.n975 0.011
R8736 VDD.n529 VDD.n528 0.011
R8737 VDD.n811 VDD.n810 0.011
R8738 VDD.n202 VDD.n200 0.011
R8739 VDD.n339 VDD.n331 0.011
R8740 VDD.n2685 VDD.n2684 0.011
R8741 VDD.n2651 VDD.n2650 0.011
R8742 VDD.n2716 VDD.n2714 0.011
R8743 VDD.n2857 VDD.n2849 0.011
R8744 VDD.n1898 VDD.n1890 0.011
R8745 VDD.n1761 VDD.n1759 0.011
R8746 VDD.n1317 VDD.n1315 0.011
R8747 VDD.n1454 VDD.n1446 0.011
R8748 VDD.n2300 VDD.n2299 0.011
R8749 VDD.n2266 VDD.n2265 0.011
R8750 VDD.n1973 VDD.n1971 0.011
R8751 VDD.n2110 VDD.n2102 0.011
R8752 VDD.n1638 VDD.n1637 0.011
R8753 VDD.n1672 VDD.n1671 0.011
R8754 VDD.n1569 VDD.n1568 0.011
R8755 VDD.n1535 VDD.n1534 0.011
R8756 VDD.n3100 VDD.n3092 0.011
R8757 VDD.n2963 VDD.n2961 0.011
R8758 VDD.n2898 VDD.n2897 0.011
R8759 VDD.n2932 VDD.n2931 0.011
R8760 VDD.n1927 VDD.n1926 0.01
R8761 VDD.n3131 VDD.n3130 0.01
R8762 VDD.n2497 VDD.n2496 0.01
R8763 VDD.n161 VDD.n160 0.009
R8764 VDD.n147 VDD.n146 0.009
R8765 VDD.n598 VDD.n596 0.009
R8766 VDD.n653 VDD.n651 0.009
R8767 VDD.n1079 VDD.n1077 0.009
R8768 VDD.n1134 VDD.n1132 0.009
R8769 VDD.n1000 VDD.n999 0.009
R8770 VDD.n986 VDD.n985 0.009
R8771 VDD.n519 VDD.n518 0.009
R8772 VDD.n505 VDD.n504 0.009
R8773 VDD.n240 VDD.n238 0.009
R8774 VDD.n295 VDD.n293 0.009
R8775 VDD.n2675 VDD.n2674 0.009
R8776 VDD.n2661 VDD.n2660 0.009
R8777 VDD.n2756 VDD.n2754 0.009
R8778 VDD.n2811 VDD.n2809 0.009
R8779 VDD.n1854 VDD.n1852 0.009
R8780 VDD.n1799 VDD.n1797 0.009
R8781 VDD.n1355 VDD.n1353 0.009
R8782 VDD.n1410 VDD.n1408 0.009
R8783 VDD.n2290 VDD.n2289 0.009
R8784 VDD.n2276 VDD.n2275 0.009
R8785 VDD.n2011 VDD.n2009 0.009
R8786 VDD.n2066 VDD.n2064 0.009
R8787 VDD.n1648 VDD.n1647 0.009
R8788 VDD.n1662 VDD.n1661 0.009
R8789 VDD.n1559 VDD.n1558 0.009
R8790 VDD.n1545 VDD.n1544 0.009
R8791 VDD.n3056 VDD.n3054 0.009
R8792 VDD.n3001 VDD.n2999 0.009
R8793 VDD.n2908 VDD.n2907 0.009
R8794 VDD.n2922 VDD.n2921 0.009
R8795 VDD.n1617 VDD.n1616 0.009
R8796 VDD VDD.n2884 0.009
R8797 VDD VDD.n1599 0.008
R8798 VDD VDD.n2 0.008
R8799 VDD.n827 VDD 0.007
R8800 VDD.n174 VDD.n173 0.007
R8801 VDD.n2317 VDD.n2316 0.007
R8802 VDD.n548 VDD.n546 0.007
R8803 VDD.n709 VDD.n701 0.007
R8804 VDD.n1029 VDD.n1027 0.007
R8805 VDD.n1190 VDD.n1182 0.007
R8806 VDD.n1013 VDD.n1012 0.007
R8807 VDD.n973 VDD.n972 0.007
R8808 VDD.n532 VDD.n531 0.007
R8809 VDD.n814 VDD.n813 0.007
R8810 VDD.n190 VDD.n188 0.007
R8811 VDD.n351 VDD.n343 0.007
R8812 VDD.n2688 VDD.n2687 0.007
R8813 VDD.n2648 VDD.n2647 0.007
R8814 VDD.n2704 VDD.n2702 0.007
R8815 VDD.n2870 VDD.n2861 0.007
R8816 VDD.n1910 VDD.n1902 0.007
R8817 VDD.n1749 VDD.n1747 0.007
R8818 VDD.n1305 VDD.n1303 0.007
R8819 VDD.n1465 VDD.n1458 0.007
R8820 VDD.n2303 VDD.n2302 0.007
R8821 VDD.n2263 VDD.n2262 0.007
R8822 VDD.n1961 VDD.n1959 0.007
R8823 VDD.n2121 VDD.n2114 0.007
R8824 VDD.n1635 VDD.n1634 0.007
R8825 VDD.n1675 VDD.n1674 0.007
R8826 VDD.n1572 VDD.n1571 0.007
R8827 VDD.n1532 VDD.n1531 0.007
R8828 VDD.n3112 VDD.n3104 0.007
R8829 VDD.n2951 VDD.n2949 0.007
R8830 VDD.n2895 VDD.n2894 0.007
R8831 VDD.n2935 VDD.n2934 0.007
R8832 VDD.n158 VDD.n157 0.005
R8833 VDD.n150 VDD.n149 0.005
R8834 VDD.n610 VDD.n608 0.005
R8835 VDD.n641 VDD.n639 0.005
R8836 VDD.n1091 VDD.n1089 0.005
R8837 VDD.n1122 VDD.n1120 0.005
R8838 VDD.n997 VDD.n996 0.005
R8839 VDD.n989 VDD.n988 0.005
R8840 VDD.n516 VDD.n515 0.005
R8841 VDD.n508 VDD.n507 0.005
R8842 VDD.n252 VDD.n250 0.005
R8843 VDD.n283 VDD.n281 0.005
R8844 VDD.n2672 VDD.n2671 0.005
R8845 VDD.n2664 VDD.n2663 0.005
R8846 VDD.n2768 VDD.n2766 0.005
R8847 VDD.n2799 VDD.n2797 0.005
R8848 VDD.n1842 VDD.n1840 0.005
R8849 VDD.n1811 VDD.n1809 0.005
R8850 VDD.n1367 VDD.n1365 0.005
R8851 VDD.n1398 VDD.n1396 0.005
R8852 VDD.n2287 VDD.n2286 0.005
R8853 VDD.n2279 VDD.n2278 0.005
R8854 VDD.n2023 VDD.n2021 0.005
R8855 VDD.n2054 VDD.n2052 0.005
R8856 VDD.n1651 VDD.n1650 0.005
R8857 VDD.n1659 VDD.n1658 0.005
R8858 VDD.n1556 VDD.n1555 0.005
R8859 VDD.n1548 VDD.n1547 0.005
R8860 VDD.n3044 VDD.n3042 0.005
R8861 VDD.n3013 VDD.n3011 0.005
R8862 VDD.n2911 VDD.n2910 0.005
R8863 VDD.n2919 VDD.n2918 0.005
R8864 VDD.n2320 VDD.n2319 0.003
R8865 VDD.n716 VDD.n713 0.003
R8866 VDD.n1197 VDD.n1194 0.003
R8867 VDD.n1594 VDD.n1593 0.003
R8868 VDD.n817 VDD.n816 0.003
R8869 VDD.n358 VDD.n355 0.003
R8870 VDD.n2482 VDD.n2481 0.003
R8871 VDD.n2877 VDD.n2874 0.003
R8872 VDD.n1917 VDD.n1914 0.003
R8873 VDD.n1293 VDD.n1291 0.003
R8874 VDD.n2306 VDD.n2305 0.003
R8875 VDD.n1949 VDD.n1947 0.003
R8876 VDD.n1632 VDD.n1631 0.003
R8877 VDD.n1575 VDD.n1574 0.003
R8878 VDD.n3119 VDD.n3116 0.003
R8879 VDD.n2892 VDD.n2891 0.003
R8880 VDD.n3136 VDD.n3135 0.002
R8881 VDD.n824 VDD.n726 0.002
R8882 VDD VDD.n823 0.002
R8883 VDD VDD.n3 0.002
R8884 VDD.n2888 VDD 0.002
R8885 VDD.n2496 VDD.n2495 0.002
R8886 VDD.n3132 VDD.n3131 0.002
R8887 VDD.n1926 VDD.n1925 0.002
R8888 VDD.n1610 VDD.n1609 0.002
R8889 VDD.n2499 VDD.n2497 0.002
R8890 VDD.n3124 VDD.n2335 0.002
R8891 VDD.n1586 VDD.n1585 0.002
R8892 VDD.n2883 VDD.n2882 0.002
R8893 VDD.n2889 VDD.n2888 0.002
R8894 VDD.n1616 VDD.n1615 0.001
R8895 VDD.n2507 VDD.n2506 0.001
R8896 VDD.n832 VDD.n831 0.001
R8897 VDD.n1589 VDD.n1588 0.001
R8898 VDD.n364 VDD.n363 0.001
R8899 VDD.n2884 VDD.n2502 0.001
R8900 VDD.n3133 VDD.n2311 0.001
R8901 VDD.n1923 VDD.n1922 0.001
R8902 VDD.n1607 VDD.n1606 0.001
R8903 VDD.n1612 VDD.n1611 0.001
R8904 VDD.n2500 VDD.n2479 0.001
R8905 VDD.n3125 VDD.n2334 0.001
R8906 VDD.n1620 VDD.n1619 0.001
R8907 VDD.n830 VDD.n820 0.001
R8908 VDD.n1934 VDD.n1933 0.001
R8909 VDD.n362 VDD.n4 0.001
R8910 VDD.n2881 VDD.n2880 0.001
R8911 VDD.n1599 VDD.n1208 0.001
R8912 VDD.n1213 VDD.n1212 0.001
R8913 VDD.n1591 VDD.n1590 0.001
R8914 VDD.n155 VDD.n154 0.001
R8915 VDD.n153 VDD.n152 0.001
R8916 VDD.n624 VDD.n622 0.001
R8917 VDD.n629 VDD.n627 0.001
R8918 VDD.n1105 VDD.n1103 0.001
R8919 VDD.n1110 VDD.n1108 0.001
R8920 VDD.n994 VDD.n993 0.001
R8921 VDD.n992 VDD.n991 0.001
R8922 VDD.n513 VDD.n512 0.001
R8923 VDD.n511 VDD.n510 0.001
R8924 VDD.n266 VDD.n264 0.001
R8925 VDD.n271 VDD.n269 0.001
R8926 VDD.n2669 VDD.n2668 0.001
R8927 VDD.n2667 VDD.n2666 0.001
R8928 VDD.n2782 VDD.n2780 0.001
R8929 VDD.n2787 VDD.n2785 0.001
R8930 VDD.n1828 VDD.n1826 0.001
R8931 VDD.n1823 VDD.n1821 0.001
R8932 VDD.n1382 VDD.n1379 0.001
R8933 VDD.n1386 VDD.n1384 0.001
R8934 VDD.n2284 VDD.n2283 0.001
R8935 VDD.n2282 VDD.n2281 0.001
R8936 VDD.n2038 VDD.n2035 0.001
R8937 VDD.n2042 VDD.n2040 0.001
R8938 VDD.n1654 VDD.n1653 0.001
R8939 VDD.n1656 VDD.n1655 0.001
R8940 VDD.n1553 VDD.n1552 0.001
R8941 VDD.n1551 VDD.n1550 0.001
R8942 VDD.n3030 VDD.n3028 0.001
R8943 VDD.n3025 VDD.n3023 0.001
R8944 VDD.n2914 VDD.n2913 0.001
R8945 VDD.n2916 VDD.n2915 0.001
R8946 VDD.n2 VDD.n1 0.001
R8947 VDD.n1921 VDD.n1920 0.001
R8948 VDD.n1921 VDD.n726 0.001
R8949 VDD.n5 VDD.n2 0.001
R8950 VDD.n2886 VDD.n2885 0.001
R8951 VDD.n3138 VDD.n3136 0.001
R8952 VDD.n826 VDD.n824 0.001
R8953 VDD.n1601 VDD.n1600 0.001
R8954 VDD.n1603 VDD.n1601 0.001
R8955 VDD.n824 VDD.n823 0.001
R8956 VDD.n3136 VDD.n3 0.001
R8957 VDD.n2888 VDD.n2886 0.001
R8958 VDD.n1599 VDD.n1598 0.001
R8959 VDD.n1605 VDD.n1604 0.001
R8960 VDD.n1597 VDD.n1591 0.001
R8961 VDD.n1585 VDD.n1213 0.001
R8962 VDD.n1603 VDD 0.001
R8963 VDD.n1928 VDD.n1927 0.001
R8964 VDD.n3130 VDD.n3129 0.001
R8965 VDD.n1626 VDD.n836 0.001
R8966 VDD.n1940 VDD.n368 0.001
R8967 VDD.n3133 VDD.n3132 0.001
R8968 VDD.n1925 VDD.n1923 0.001
R8969 VDD.n1609 VDD.n1607 0.001
R8970 VDD.n1614 VDD.n1612 0.001
R8971 VDD.n2500 VDD.n2499 0.001
R8972 VDD.n2884 VDD.n2883 0.001
R8973 VDD.n2889 VDD.n2501 0.001
R8974 VDD.n2882 VDD.n2881 0.001
R8975 VDD.n3125 VDD.n3124 0.001
R8976 VDD.n362 VDD.n361 0.001
R8977 VDD.n830 VDD.n829 0.001
R8978 VDD.n1626 VDD.n1620 0.001
R8979 VDD.n1940 VDD.n1934 0.001
R8980 VDD.n1598 VDD.n1597 0.001
R8981 VDD.n1604 VDD.n1603 0.001
R8982 VDD.n361 VDD.n5 0.001
R8983 VDD.n829 VDD.n828 0.001
R8984 VDD.n1615 VDD.n1206 0.001
R8985 VDD.n3129 VDD.n3128 0.001
R8986 VDD.n3128 VDD.n2330 0.001
R8987 VDD.n1930 VDD.n1928 0.001
R8988 VDD.n1930 VDD.n1929 0.001
R8989 VDD.n1615 VDD.n1614 0.001
R8990 VDD.n828 VDD.n827 0.001
R8991 VDD.n827 VDD.n822 0.001
R8992 VDD.n3135 VDD.n3134 0.001
R8993 VDD.n3134 VDD.n2309 0.001
R8994 VDD.n2495 VDD.n2494 0.001
R8995 VDD.n2494 VDD.n2492 0.001
R8996 VDD.n2505 VDD.n2504 0.001
R8997 VDD.n2506 VDD.n2505 0.001
R8998 VDD.n367 VDD.n366 0.001
R8999 VDD.n367 VDD.n364 0.001
R9000 VDD.n1587 VDD.n1210 0.001
R9001 VDD.n1588 VDD.n1587 0.001
R9002 VDD.n835 VDD.n834 0.001
R9003 VDD.n835 VDD.n832 0.001
R9004 a_n18753_11548.n97 a_n18753_11548.t4 1040.33
R9005 a_n18753_11548.n97 a_n18753_11548.t5 794.533
R9006 a_n18753_11548.n46 a_n18753_11548.n45 13.176
R9007 a_n18753_11548.n98 a_n18753_11548.t2 11.611
R9008 a_n18753_11548.n98 a_n18753_11548.t1 11.295
R9009 a_n18753_11548.n142 a_n18753_11548.n39 9.3
R9010 a_n18753_11548.n142 a_n18753_11548.n138 9.3
R9011 a_n18753_11548.n142 a_n18753_11548.n132 9.3
R9012 a_n18753_11548.n142 a_n18753_11548.n58 9.3
R9013 a_n18753_11548.n142 a_n18753_11548.n66 9.3
R9014 a_n18753_11548.n142 a_n18753_11548.n127 9.3
R9015 a_n18753_11548.n101 a_n18753_11548.t0 9.017
R9016 a_n18753_11548.n142 a_n18753_11548.n122 8.47
R9017 a_n18753_11548.n142 a_n18753_11548.n141 8.469
R9018 a_n18753_11548.n142 a_n18753_11548.n119 8.124
R9019 a_n18753_11548.n142 a_n18753_11548.n29 8.124
R9020 a_n18753_11548.n142 a_n18753_11548.n34 8.097
R9021 a_n18753_11548.n142 a_n18753_11548.n114 8.097
R9022 a_n18753_11548.n142 a_n18753_11548.n61 8.016
R9023 a_n18753_11548.n142 a_n18753_11548.n44 8.016
R9024 a_n18753_11548.n142 a_n18753_11548.n53 7.964
R9025 a_n18753_11548.n142 a_n18753_11548.n49 7.964
R9026 a_n18753_11548.n60 a_n18753_11548.n59 6.4
R9027 a_n18753_11548.n113 a_n18753_11548.n67 6.4
R9028 a_n18753_11548.n32 a_n18753_11548.n31 6.023
R9029 a_n18753_11548.n42 a_n18753_11548.n41 6.023
R9030 a_n18753_11548.n132 a_n18753_11548.n131 6.023
R9031 a_n18753_11548.n48 a_n18753_11548.n47 6.023
R9032 a_n18753_11548.n52 a_n18753_11548.n51 6.023
R9033 a_n18753_11548.n140 a_n18753_11548.n139 5.647
R9034 a_n18753_11548.n58 a_n18753_11548.n55 5.647
R9035 a_n18753_11548.n117 a_n18753_11548.n116 5.647
R9036 a_n18753_11548.n121 a_n18753_11548.n120 5.647
R9037 a_n18753_11548.n129 a_n18753_11548.n128 5.457
R9038 a_n18753_11548.n27 a_n18753_11548.n26 5.27
R9039 a_n18753_11548.n57 a_n18753_11548.n56 5.08
R9040 a_n18753_11548.n39 a_n18753_11548.n38 4.517
R9041 a_n18753_11548.n127 a_n18753_11548.n124 4.517
R9042 a_n18753_11548.n75 a_n18753_11548.n74 4.5
R9043 a_n18753_11548.n2 a_n18753_11548.n1 4.5
R9044 a_n18753_11548.n36 a_n18753_11548.n35 4.314
R9045 a_n18753_11548.n137 a_n18753_11548.n136 4.141
R9046 a_n18753_11548.n63 a_n18753_11548.n62 4.141
R9047 a_n18753_11548.n134 a_n18753_11548.n133 3.944
R9048 a_n18753_11548.n126 a_n18753_11548.n125 3.937
R9049 a_n18753_11548.n65 a_n18753_11548.n64 3.567
R9050 a_n18753_11548.n104 a_n18753_11548.n97 3.396
R9051 a_n18753_11548.n113 a_n18753_11548.n112 3.033
R9052 a_n18753_11548.t3 a_n18753_11548.n142 2.9
R9053 a_n18753_11548.n105 a_n18753_11548.n104 2.397
R9054 a_n18753_11548.n138 a_n18753_11548.n137 2.258
R9055 a_n18753_11548.n66 a_n18753_11548.n63 2.258
R9056 a_n18753_11548.n102 a_n18753_11548.n101 2.237
R9057 a_n18753_11548.n38 a_n18753_11548.n37 1.882
R9058 a_n18753_11548.n124 a_n18753_11548.n123 1.882
R9059 a_n18753_11548.n66 a_n18753_11548.n65 1.505
R9060 a_n18753_11548.n94 a_n18753_11548.n106 1.5
R9061 a_n18753_11548.n76 a_n18753_11548.n78 1.5
R9062 a_n18753_11548.n75 a_n18753_11548.n73 1.5
R9063 a_n18753_11548.n21 a_n18753_11548.n24 1.5
R9064 a_n18753_11548.n12 a_n18753_11548.n11 1.5
R9065 a_n18753_11548.n112 a_n18753_11548.n92 1.5
R9066 a_n18753_11548.n28 a_n18753_11548.n27 1.129
R9067 a_n18753_11548.n26 a_n18753_11548.n25 1.129
R9068 a_n18753_11548.n138 a_n18753_11548.n134 1.129
R9069 a_n18753_11548.n136 a_n18753_11548.n135 1.129
R9070 a_n18753_11548.n104 a_n18753_11548.n103 1.022
R9071 a_n18753_11548.n141 a_n18753_11548.n140 0.752
R9072 a_n18753_11548.n55 a_n18753_11548.n54 0.752
R9073 a_n18753_11548.n58 a_n18753_11548.n57 0.752
R9074 a_n18753_11548.n127 a_n18753_11548.n126 0.752
R9075 a_n18753_11548.n116 a_n18753_11548.n115 0.752
R9076 a_n18753_11548.n118 a_n18753_11548.n117 0.752
R9077 a_n18753_11548.n122 a_n18753_11548.n121 0.752
R9078 a_n18753_11548.n53 a_n18753_11548.n52 0.536
R9079 a_n18753_11548.n49 a_n18753_11548.n48 0.536
R9080 a_n18753_11548.n61 a_n18753_11548.n60 0.475
R9081 a_n18753_11548.n44 a_n18753_11548.n43 0.475
R9082 a_n18753_11548.n34 a_n18753_11548.n33 0.382
R9083 a_n18753_11548.n114 a_n18753_11548.n113 0.382
R9084 a_n18753_11548.n33 a_n18753_11548.n32 0.376
R9085 a_n18753_11548.n31 a_n18753_11548.n30 0.376
R9086 a_n18753_11548.n39 a_n18753_11548.n36 0.376
R9087 a_n18753_11548.n43 a_n18753_11548.n42 0.376
R9088 a_n18753_11548.n41 a_n18753_11548.n40 0.376
R9089 a_n18753_11548.n132 a_n18753_11548.n129 0.376
R9090 a_n18753_11548.n131 a_n18753_11548.n130 0.376
R9091 a_n18753_11548.n47 a_n18753_11548.n46 0.376
R9092 a_n18753_11548.n51 a_n18753_11548.n50 0.376
R9093 a_n18753_11548.n29 a_n18753_11548.n28 0.349
R9094 a_n18753_11548.n119 a_n18753_11548.n118 0.349
R9095 a_n18753_11548.n99 a_n18753_11548.n98 0.276
R9096 a_n18753_11548.n94 a_n18753_11548.n93 0.15
R9097 a_n18753_11548.n105 a_n18753_11548.n95 0.148
R9098 a_n18753_11548.n2 a_n18753_11548.n0 0.066
R9099 a_n18753_11548.n84 a_n18753_11548.n83 0.043
R9100 a_n18753_11548.n80 a_n18753_11548.n79 0.043
R9101 a_n18753_11548.n76 a_n18753_11548.n75 0.041
R9102 a_n18753_11548.n102 a_n18753_11548.n99 0.039
R9103 a_n18753_11548.n91 a_n18753_11548.n90 0.035
R9104 a_n18753_11548.n111 a_n18753_11548.n110 0.035
R9105 a_n18753_11548.n19 a_n18753_11548.n18 0.034
R9106 a_n18753_11548.n23 a_n18753_11548.n22 0.034
R9107 a_n18753_11548.n8 a_n18753_11548.n7 0.034
R9108 a_n18753_11548.n89 a_n18753_11548.n88 0.034
R9109 a_n18753_11548.n109 a_n18753_11548.n108 0.034
R9110 a_n18753_11548.n12 a_n18753_11548.n6 0.032
R9111 a_n18753_11548.n112 a_n18753_11548.n82 0.032
R9112 a_n18753_11548.n101 a_n18753_11548.n100 0.032
R9113 a_n18753_11548.n9 a_n18753_11548.n8 0.03
R9114 a_n18753_11548.n87 a_n18753_11548.n86 0.03
R9115 a_n18753_11548.n11 a_n18753_11548.n10 0.028
R9116 a_n18753_11548.n72 a_n18753_11548.n70 0.028
R9117 a_n18753_11548.n85 a_n18753_11548.n84 0.028
R9118 a_n18753_11548.n13 a_n18753_11548.n12 0.028
R9119 a_n18753_11548.n69 a_n18753_11548.n68 0.028
R9120 a_n18753_11548.n81 a_n18753_11548.n80 0.028
R9121 a_n18753_11548.n107 a_n18753_11548.n94 0.028
R9122 a_n18753_11548.n17 a_n18753_11548.n15 0.026
R9123 a_n18753_11548.n78 a_n18753_11548.n77 0.026
R9124 a_n18753_11548.n4 a_n18753_11548.n3 0.026
R9125 a_n18753_11548.n18 a_n18753_11548.n17 0.024
R9126 a_n18753_11548.n6 a_n18753_11548.n5 0.024
R9127 a_n18753_11548.n15 a_n18753_11548.n16 0.022
R9128 a_n18753_11548.n5 a_n18753_11548.n4 0.022
R9129 a_n18753_11548.n3 a_n18753_11548.n2 0.022
R9130 a_n18753_11548.n20 a_n18753_11548.n19 0.02
R9131 a_n18753_11548.n10 a_n18753_11548.n9 0.02
R9132 a_n18753_11548.n14 a_n18753_11548.n13 0.02
R9133 a_n18753_11548.n106 a_n18753_11548.n105 0.018
R9134 a_n18753_11548.n82 a_n18753_11548.n81 0.018
R9135 a_n18753_11548.n24 a_n18753_11548.n23 0.017
R9136 a_n18753_11548.n86 a_n18753_11548.n85 0.017
R9137 a_n18753_11548.n70 a_n18753_11548.n71 0.015
R9138 a_n18753_11548.n73 a_n18753_11548.n72 0.015
R9139 a_n18753_11548.n68 a_n18753_11548.n0 0.015
R9140 a_n18753_11548.n75 a_n18753_11548.n69 0.015
R9141 a_n18753_11548.n92 a_n18753_11548.n91 0.013
R9142 a_n18753_11548.n90 a_n18753_11548.n89 0.013
R9143 a_n18753_11548.n112 a_n18753_11548.n111 0.013
R9144 a_n18753_11548.n110 a_n18753_11548.n109 0.013
R9145 a_n18753_11548.n95 a_n18753_11548.n96 0.007
R9146 a_n18753_11548.n21 a_n18753_11548.n20 1.424
R9147 a_n18753_11548.n79 a_n18753_11548.n76 0.005
R9148 a_n18753_11548.n92 a_n18753_11548.n87 0.003
R9149 a_n18753_11548.n108 a_n18753_11548.n107 0.003
R9150 a_n18753_11548.n103 a_n18753_11548.n102 0.001
R9151 a_n18753_11548.n14 a_n18753_11548.n21 0.47
R9152 fout1.n118 fout1.t14 1038.95
R9153 fout1.n139 fout1.t4 1037.29
R9154 fout1.n140 fout1.t12 797.185
R9155 fout1.n110 fout1.t9 795.565
R9156 fout1.n509 fout1.t6 732.331
R9157 fout1.n80 fout1.t10 731.671
R9158 fout1.n23 fout1.t13 731.671
R9159 fout1.n0 fout1.t11 730.672
R9160 fout1.n43 fout1.t5 400.618
R9161 fout1.n86 fout1.t3 400.616
R9162 fout1.n524 fout1.t8 397.315
R9163 fout1.n0 fout1.t7 395.84
R9164 fout1.n349 fout1.n348 13.176
R9165 fout1.n161 fout1.t0 11.724
R9166 fout1.n161 fout1.t2 10.994
R9167 fout1.n169 fout1.n167 9.3
R9168 fout1.n471 fout1.n470 9.3
R9169 fout1.n217 fout1.n216 9.3
R9170 fout1.n219 fout1.n218 9.3
R9171 fout1.n277 fout1.n276 9.3
R9172 fout1.n274 fout1.n273 9.3
R9173 fout1.n231 fout1.n230 9.3
R9174 fout1.n229 fout1.n228 9.3
R9175 fout1.n355 fout1.n354 9.3
R9176 fout1.n255 fout1.n254 9.3
R9177 fout1.n263 fout1.n262 9.3
R9178 fout1.n266 fout1.n265 9.3
R9179 fout1.n385 fout1.n384 9.3
R9180 fout1.n382 fout1.n381 9.3
R9181 fout1.n466 fout1.n465 9.3
R9182 fout1.n464 fout1.n463 9.3
R9183 fout1.n457 fout1.n456 8.097
R9184 fout1.n265 fout1.n264 5.457
R9185 fout1.n384 fout1.n383 5.08
R9186 fout1.n455 fout1.n454 4.65
R9187 fout1.n394 fout1.n393 4.65
R9188 fout1.n476 fout1.n469 4.5
R9189 fout1.n450 fout1.n449 4.5
R9190 fout1.n443 fout1.n442 4.5
R9191 fout1.n374 fout1.n373 4.5
R9192 fout1.n364 fout1.n363 4.5
R9193 fout1.n351 fout1.n350 4.5
R9194 fout1.n327 fout1.n326 4.5
R9195 fout1.n260 fout1.n251 4.5
R9196 fout1.n283 fout1.n282 4.5
R9197 fout1.n227 fout1.n226 4.5
R9198 fout1.n239 fout1.n238 4.5
R9199 fout1.n246 fout1.n245 4.5
R9200 fout1.n291 fout1.n290 4.5
R9201 fout1.n271 fout1.n270 4.5
R9202 fout1.n436 fout1.n435 4.5
R9203 fout1.n215 fout1.n214 4.5
R9204 fout1.n485 fout1.n482 4.5
R9205 fout1.n172 fout1.n171 4.5
R9206 fout1.n238 fout1.n236 4.314
R9207 fout1.n290 fout1.n287 3.944
R9208 fout1.n449 fout1.n448 3.937
R9209 fout1.n435 fout1.n434 3.567
R9210 fout1.n395 fout1.n388 3.033
R9211 fout1.n459 fout1.n458 3.033
R9212 fout1.n456 fout1.t1 2.9
R9213 fout1.n289 fout1.n288 2.258
R9214 fout1.n433 fout1.n432 2.258
R9215 fout1.n244 fout1.n243 1.882
R9216 fout1.n245 fout1.n244 1.882
R9217 fout1.n441 fout1.n440 1.882
R9218 fout1.n497 fout1.n161 1.517
R9219 fout1.n435 fout1.n433 1.505
R9220 fout1.n442 fout1.n441 1.505
R9221 fout1.n477 fout1.n476 1.5
R9222 fout1.n328 fout1.n327 1.5
R9223 fout1.n365 fout1.n364 1.5
R9224 fout1.n396 fout1.n395 1.5
R9225 fout1.n375 fout1.n374 1.5
R9226 fout1.n486 fout1.n485 1.5
R9227 fout1.n173 fout1.n172 1.5
R9228 fout1.n66 fout1.n64 1.435
R9229 fout1.n32 fout1.n31 1.435
R9230 fout1.n153 fout1.n139 1.388
R9231 fout1.n141 fout1.n140 1.355
R9232 fout1.n120 fout1.n118 1.354
R9233 fout1.n111 fout1.n110 1.354
R9234 fout1.n526 fout1.n524 1.354
R9235 fout1.n510 fout1.n509 1.354
R9236 fout1.n81 fout1.n80 1.354
R9237 fout1.n24 fout1.n23 1.354
R9238 fout1.n527 fout1.n526 1.142
R9239 fout1.n112 fout1.n111 1.142
R9240 fout1.n67 fout1.n66 1.142
R9241 fout1.n25 fout1.n24 1.142
R9242 fout1.n528 fout1.n527 1.138
R9243 fout1.n113 fout1.n112 1.138
R9244 fout1.n26 fout1.n25 1.138
R9245 fout1.n68 fout1.n67 1.138
R9246 fout1.n511 fout1.n510 1.137
R9247 fout1.n537 fout1.n536 1.137
R9248 fout1.n502 fout1.n501 1.137
R9249 fout1.n532 fout1.n531 1.137
R9250 fout1.n517 fout1.n516 1.137
R9251 fout1.n96 fout1.n95 1.137
R9252 fout1.n126 fout1.n125 1.137
R9253 fout1.n92 fout1.n91 1.137
R9254 fout1.n102 fout1.n101 1.137
R9255 fout1.n121 fout1.n120 1.137
R9256 fout1.n82 fout1.n81 1.137
R9257 fout1.n52 fout1.n51 1.137
R9258 fout1.n73 fout1.n72 1.137
R9259 fout1.n49 fout1.n48 1.137
R9260 fout1.n58 fout1.n57 1.137
R9261 fout1.n9 fout1.n8 1.137
R9262 fout1.n38 fout1.n37 1.137
R9263 fout1.n4 fout1.n3 1.137
R9264 fout1.n15 fout1.n14 1.137
R9265 fout1.n33 fout1.n32 1.137
R9266 fout1.n539 fout1.n538 1.136
R9267 fout1.n11 fout1.n10 1.136
R9268 fout1.n54 fout1.n53 1.136
R9269 fout1.n513 fout1.n512 1.136
R9270 fout1.n84 fout1.n83 1.136
R9271 fout1.n129 fout1.n128 1.136
R9272 fout1.n98 fout1.n97 1.136
R9273 fout1.n41 fout1.n40 1.136
R9274 fout1.n214 fout1.n213 1.129
R9275 fout1.n290 fout1.n289 1.129
R9276 fout1.n282 fout1.n281 1.129
R9277 fout1.n292 fout1.n291 1.042
R9278 fout1.n185 fout1.n184 0.853
R9279 fout1.n309 fout1.n308 0.853
R9280 fout1.n398 fout1.n397 0.853
R9281 fout1.n492 fout1.n491 0.853
R9282 fout1.n541 fout1.n160 0.823
R9283 fout1.n171 fout1.n170 0.752
R9284 fout1.n363 fout1.n362 0.752
R9285 fout1.n373 fout1.n372 0.752
R9286 fout1.n449 fout1.n447 0.752
R9287 fout1.n469 fout1.n468 0.752
R9288 fout1.n482 fout1.n481 0.752
R9289 fout1.n175 fout1.n174 0.717
R9290 fout1.n497 fout1.n496 0.69
R9291 fout1.n498 fout1.n497 0.68
R9292 fout1.n354 fout1.n353 0.536
R9293 fout1.n254 fout1.n253 0.536
R9294 fout1.n276 fout1.n275 0.475
R9295 fout1.n393 fout1.n392 0.475
R9296 fout1.n541 fout1.n540 0.471
R9297 fout1.n154 fout1.n153 0.44
R9298 fout1.n458 fout1.n457 0.382
R9299 fout1.n225 fout1.n224 0.382
R9300 fout1.n226 fout1.n225 0.376
R9301 fout1.n238 fout1.n237 0.376
R9302 fout1.n270 fout1.n269 0.376
R9303 fout1.n251 fout1.n250 0.376
R9304 fout1.n326 fout1.n325 0.376
R9305 fout1.n350 fout1.n349 0.376
R9306 fout1.n213 fout1.n212 0.349
R9307 fout1.n468 fout1.n467 0.349
R9308 fout1 fout1.n541 0.243
R9309 fout1.n88 fout1.n87 0.152
R9310 fout1.n43 fout1.n42 0.123
R9311 fout1.n86 fout1.n85 0.123
R9312 fout1.n44 fout1.n43 0.091
R9313 fout1.n524 fout1.n523 0.083
R9314 fout1.n509 fout1.n508 0.083
R9315 fout1.n80 fout1.n79 0.083
R9316 fout1.n23 fout1.n22 0.083
R9317 fout1.n118 fout1.n117 0.076
R9318 fout1.n110 fout1.n109 0.076
R9319 fout1.n139 fout1.n138 0.075
R9320 fout1 fout1.n130 0.073
R9321 fout1.n87 fout1.n86 0.07
R9322 fout1.n135 fout1.n134 0.058
R9323 fout1.n267 fout1.n266 0.047
R9324 fout1.n257 fout1.n256 0.047
R9325 fout1.n345 fout1.n344 0.047
R9326 fout1.n358 fout1.n357 0.047
R9327 fout1.n386 fout1.n385 0.047
R9328 fout1.n473 fout1.n472 0.047
R9329 fout1.n452 fout1.n451 0.043
R9330 fout1.n421 fout1.n420 0.043
R9331 fout1.n235 fout1.n234 0.041
R9332 fout1.n202 fout1.n201 0.041
R9333 fout1.n461 fout1.n460 0.035
R9334 fout1.n329 fout1.n328 0.035
R9335 fout1.n334 fout1.n333 0.035
R9336 fout1.n427 fout1.n426 0.035
R9337 fout1.n222 fout1.n221 0.034
R9338 fout1.n343 fout1.n342 0.034
R9339 fout1.n347 fout1.n346 0.034
R9340 fout1.n464 fout1.n462 0.034
R9341 fout1.n182 fout1.n181 0.034
R9342 fout1.n180 fout1.n179 0.034
R9343 fout1.n299 fout1.n298 0.034
R9344 fout1.n306 fout1.n305 0.034
R9345 fout1.n365 fout1.n341 0.034
R9346 fout1.n367 fout1.n366 0.034
R9347 fout1.n380 fout1.n379 0.034
R9348 fout1.n429 fout1.n428 0.034
R9349 fout1.n536 fout1.n534 0.032
R9350 fout1.n149 fout1.n148 0.032
R9351 fout1.n148 fout1.n147 0.032
R9352 fout1.n220 fout1.n219 0.032
R9353 fout1.n395 fout1.n394 0.032
R9354 fout1.n459 fout1.n455 0.032
R9355 fout1.n304 fout1.n303 0.032
R9356 fout1.n477 fout1.n429 0.032
R9357 fout1.n91 fout1.n90 0.032
R9358 fout1.n48 fout1.n47 0.032
R9359 fout1.n8 fout1.n6 0.032
R9360 fout1.n153 fout1.n152 0.032
R9361 fout1.n187 fout1.n186 0.031
R9362 fout1.n198 fout1.n197 0.031
R9363 fout1.n411 fout1.n410 0.031
R9364 fout1.n494 fout1.n493 0.031
R9365 fout1.n143 fout1.n142 0.03
R9366 fout1.n229 fout1.n227 0.03
R9367 fout1.n274 fout1.n272 0.03
R9368 fout1.n259 fout1.n258 0.03
R9369 fout1.n360 fout1.n359 0.03
R9370 fout1.n474 fout1.n473 0.03
R9371 fout1.n183 fout1.n182 0.03
R9372 fout1.n177 fout1.n176 0.03
R9373 fout1.n302 fout1.n301 0.03
R9374 fout1.n339 fout1.n338 0.03
R9375 fout1.n368 fout1.n367 0.03
R9376 fout1.n424 fout1.n423 0.03
R9377 fout1.n491 fout1.n490 0.03
R9378 fout1.n311 fout1.n310 0.03
R9379 fout1.n322 fout1.n321 0.03
R9380 fout1.n400 fout1.n399 0.03
R9381 fout1.n523 fout1.n522 0.028
R9382 fout1.n521 fout1.n520 0.028
R9383 fout1.n506 fout1.n505 0.028
R9384 fout1.n508 fout1.n507 0.028
R9385 fout1.n516 fout1.n515 0.028
R9386 fout1.n531 fout1.n530 0.028
R9387 fout1.n536 fout1.n535 0.028
R9388 fout1.n501 fout1.n499 0.028
R9389 fout1.n152 fout1.n151 0.028
R9390 fout1.n150 fout1.n149 0.028
R9391 fout1.n147 fout1.n146 0.028
R9392 fout1.n145 fout1.n144 0.028
R9393 fout1.n172 fout1.n169 0.028
R9394 fout1.n210 fout1.n209 0.028
R9395 fout1.n233 fout1.n232 0.028
R9396 fout1.n248 fout1.n247 0.028
R9397 fout1.n291 fout1.n249 0.028
R9398 fout1.n280 fout1.n279 0.028
R9399 fout1.n395 fout1.n387 0.028
R9400 fout1.n439 fout1.n438 0.028
R9401 fout1.n453 fout1.n452 0.028
R9402 fout1.n476 fout1.n466 0.028
R9403 fout1.n173 fout1.n165 0.028
R9404 fout1.n200 fout1.n199 0.028
R9405 fout1.n207 fout1.n206 0.028
R9406 fout1.n292 fout1.n208 0.028
R9407 fout1.n297 fout1.n296 0.028
R9408 fout1.n307 fout1.n306 0.028
R9409 fout1.n324 fout1.n323 0.028
R9410 fout1.n336 fout1.n335 0.028
R9411 fout1.n397 fout1.n396 0.028
R9412 fout1.n416 fout1.n415 0.028
R9413 fout1.n422 fout1.n421 0.028
R9414 fout1.n487 fout1.n486 0.028
R9415 fout1.n125 fout1.n124 0.028
R9416 fout1.n91 fout1.n89 0.028
R9417 fout1.n95 fout1.n94 0.028
R9418 fout1.n101 fout1.n99 0.028
R9419 fout1.n64 fout1.n63 0.028
R9420 fout1.n62 fout1.n61 0.028
R9421 fout1.n77 fout1.n76 0.028
R9422 fout1.n79 fout1.n78 0.028
R9423 fout1.n57 fout1.n56 0.028
R9424 fout1.n48 fout1.n46 0.028
R9425 fout1.n51 fout1.n50 0.028
R9426 fout1.n72 fout1.n70 0.028
R9427 fout1.n31 fout1.n30 0.028
R9428 fout1.n29 fout1.n28 0.028
R9429 fout1.n20 fout1.n19 0.028
R9430 fout1.n22 fout1.n21 0.028
R9431 fout1.n37 fout1.n36 0.028
R9432 fout1.n3 fout1.n2 0.028
R9433 fout1.n8 fout1.n7 0.028
R9434 fout1.n14 fout1.n12 0.028
R9435 fout1.n191 fout1.n190 0.027
R9436 fout1.n194 fout1.n193 0.027
R9437 fout1.n217 fout1.n215 0.026
R9438 fout1.n271 fout1.n268 0.026
R9439 fout1.n390 fout1.n389 0.026
R9440 fout1.n437 fout1.n436 0.026
R9441 fout1.n294 fout1.n293 0.026
R9442 fout1.n308 fout1.n300 0.026
R9443 fout1.n378 fout1.n377 0.026
R9444 fout1.n414 fout1.n413 0.026
R9445 fout1.n419 fout1.n418 0.026
R9446 fout1.n489 fout1.n488 0.026
R9447 fout1.n315 fout1.n314 0.026
R9448 fout1.n318 fout1.n317 0.026
R9449 fout1.n404 fout1.n403 0.026
R9450 fout1.n407 fout1.n406 0.026
R9451 fout1.n117 fout1.n116 0.026
R9452 fout1.n115 fout1.n114 0.026
R9453 fout1.n107 fout1.n106 0.026
R9454 fout1.n109 fout1.n108 0.026
R9455 fout1.n138 fout1.n137 0.025
R9456 fout1.n136 fout1.n135 0.025
R9457 fout1.n134 fout1.n133 0.025
R9458 fout1.n132 fout1.n131 0.025
R9459 fout1.n174 fout1.n173 0.024
R9460 fout1.n278 fout1.n277 0.024
R9461 fout1.n394 fout1.n391 0.024
R9462 fout1.n164 fout1.n163 0.024
R9463 fout1.n204 fout1.n203 0.024
R9464 fout1.n300 fout1.n299 0.024
R9465 fout1.n332 fout1.n331 0.024
R9466 fout1.n375 fout1.n369 0.024
R9467 fout1.n157 fout1.n156 0.023
R9468 fout1.n241 fout1.n240 0.022
R9469 fout1.n268 fout1.n267 0.022
R9470 fout1.n255 fout1.n252 0.022
R9471 fout1.n355 fout1.n352 0.022
R9472 fout1.n391 fout1.n390 0.022
R9473 fout1.n446 fout1.n445 0.022
R9474 fout1.n163 fout1.n162 0.022
R9475 fout1.n308 fout1.n307 0.022
R9476 fout1.n331 fout1.n330 0.022
R9477 fout1.n396 fout1.n380 0.022
R9478 fout1.n379 fout1.n378 0.022
R9479 fout1.n285 fout1.n284 0.02
R9480 fout1.n283 fout1.n280 0.02
R9481 fout1.n279 fout1.n278 0.02
R9482 fout1.n387 fout1.n386 0.02
R9483 fout1.n371 fout1.n370 0.02
R9484 fout1.n184 fout1.n183 0.02
R9485 fout1.n298 fout1.n297 0.02
R9486 fout1.n397 fout1.n368 0.02
R9487 fout1.n490 fout1.n489 0.02
R9488 fout1.n486 fout1.n480 0.02
R9489 fout1.n185 fout1.n175 0.019
R9490 fout1.n186 fout1.n185 0.019
R9491 fout1.n492 fout1.n411 0.019
R9492 fout1.n493 fout1.n492 0.019
R9493 fout1.n455 fout1.n453 0.018
R9494 fout1.n205 fout1.n204 0.018
R9495 fout1.n491 fout1.n477 0.018
R9496 fout1.n309 fout1.n198 0.018
R9497 fout1.n310 fout1.n309 0.018
R9498 fout1.n398 fout1.n322 0.018
R9499 fout1.n399 fout1.n398 0.018
R9500 fout1.n526 fout1.n525 0.017
R9501 fout1.n516 fout1.n514 0.017
R9502 fout1.n501 fout1.n500 0.017
R9503 fout1.n510 fout1.n504 0.017
R9504 fout1.n144 fout1.n143 0.017
R9505 fout1.n142 fout1.n141 0.017
R9506 fout1.n232 fout1.n231 0.017
R9507 fout1.n261 fout1.n260 0.017
R9508 fout1.n258 fout1.n257 0.017
R9509 fout1.n484 fout1.n483 0.017
R9510 fout1.n293 fout1.n292 0.017
R9511 fout1.n296 fout1.n295 0.017
R9512 fout1.n305 fout1.n304 0.017
R9513 fout1.n303 fout1.n302 0.017
R9514 fout1.n377 fout1.n376 0.017
R9515 fout1.n418 fout1.n417 0.017
R9516 fout1.n423 fout1.n422 0.017
R9517 fout1.n480 fout1.n479 0.017
R9518 fout1.n120 fout1.n119 0.017
R9519 fout1.n125 fout1.n123 0.017
R9520 fout1.n101 fout1.n100 0.017
R9521 fout1.n111 fout1.n105 0.017
R9522 fout1.n66 fout1.n65 0.017
R9523 fout1.n57 fout1.n55 0.017
R9524 fout1.n72 fout1.n71 0.017
R9525 fout1.n81 fout1.n75 0.017
R9526 fout1.n32 fout1.n27 0.017
R9527 fout1.n37 fout1.n35 0.017
R9528 fout1.n14 fout1.n13 0.017
R9529 fout1.n24 fout1.n18 0.017
R9530 fout1.n532 fout1.n529 0.016
R9531 fout1.n537 fout1.n533 0.016
R9532 fout1.n96 fout1.n93 0.016
R9533 fout1.n49 fout1.n45 0.016
R9534 fout1.n9 fout1.n5 0.016
R9535 fout1.n522 fout1.n521 0.015
R9536 fout1.n507 fout1.n506 0.015
R9537 fout1.n151 fout1.n150 0.015
R9538 fout1.n146 fout1.n145 0.015
R9539 fout1.n211 fout1.n210 0.015
R9540 fout1.n221 fout1.n220 0.015
R9541 fout1.n249 fout1.n248 0.015
R9542 fout1.n359 fout1.n358 0.015
R9543 fout1.n364 fout1.n361 0.015
R9544 fout1.n438 fout1.n437 0.015
R9545 fout1.n443 fout1.n439 0.015
R9546 fout1.n475 fout1.n474 0.015
R9547 fout1.n181 fout1.n180 0.015
R9548 fout1.n179 fout1.n178 0.015
R9549 fout1.n208 fout1.n207 0.015
R9550 fout1.n338 fout1.n337 0.015
R9551 fout1.n341 fout1.n340 0.015
R9552 fout1.n366 fout1.n365 0.015
R9553 fout1.n415 fout1.n414 0.015
R9554 fout1.n417 fout1.n416 0.015
R9555 fout1.n63 fout1.n62 0.015
R9556 fout1.n78 fout1.n77 0.015
R9557 fout1.n30 fout1.n29 0.015
R9558 fout1.n21 fout1.n20 0.015
R9559 fout1.n137 fout1.n136 0.013
R9560 fout1.n133 fout1.n132 0.013
R9561 fout1.n223 fout1.n222 0.013
R9562 fout1.n247 fout1.n246 0.013
R9563 fout1.n263 fout1.n261 0.013
R9564 fout1.n460 fout1.n459 0.013
R9565 fout1.n462 fout1.n461 0.013
R9566 fout1.n206 fout1.n205 0.013
R9567 fout1.n426 fout1.n425 0.013
R9568 fout1.n428 fout1.n427 0.013
R9569 fout1.n496 fout1.n495 0.013
R9570 fout1.n116 fout1.n115 0.013
R9571 fout1.n108 fout1.n107 0.013
R9572 fout1.n538 fout1.n532 0.012
R9573 fout1.n538 fout1.n537 0.012
R9574 fout1.n192 fout1.n191 0.012
R9575 fout1.n193 fout1.n192 0.012
R9576 fout1.n97 fout1.n92 0.012
R9577 fout1.n97 fout1.n96 0.012
R9578 fout1.n53 fout1.n49 0.012
R9579 fout1.n53 fout1.n52 0.012
R9580 fout1.n10 fout1.n4 0.012
R9581 fout1.n10 fout1.n9 0.012
R9582 fout1.n519 fout1.n518 0.011
R9583 fout1.n512 fout1.n503 0.011
R9584 fout1.n286 fout1.n285 0.011
R9585 fout1.n189 fout1.n188 0.011
R9586 fout1.n196 fout1.n195 0.011
R9587 fout1.n313 fout1.n312 0.011
R9588 fout1.n316 fout1.n315 0.011
R9589 fout1.n317 fout1.n316 0.011
R9590 fout1.n320 fout1.n319 0.011
R9591 fout1.n402 fout1.n401 0.011
R9592 fout1.n405 fout1.n404 0.011
R9593 fout1.n406 fout1.n405 0.011
R9594 fout1.n409 fout1.n408 0.011
R9595 fout1.n128 fout1.n127 0.011
R9596 fout1.n104 fout1.n103 0.011
R9597 fout1.n60 fout1.n59 0.011
R9598 fout1.n83 fout1.n74 0.011
R9599 fout1.n40 fout1.n39 0.011
R9600 fout1.n17 fout1.n16 0.011
R9601 fout1.n126 fout1.n122 0.01
R9602 fout1.n73 fout1.n69 0.01
R9603 fout1.n38 fout1.n34 0.01
R9604 fout1.n155 fout1.n154 0.01
R9605 fout1.n156 fout1.n155 0.01
R9606 fout1.n159 fout1.n158 0.009
R9607 fout1.n169 fout1.n168 0.009
R9608 fout1.n242 fout1.n241 0.009
R9609 fout1.n246 fout1.n242 0.009
R9610 fout1.n344 fout1.n343 0.009
R9611 fout1.n445 fout1.n444 0.009
R9612 fout1.n165 fout1.n164 0.009
R9613 fout1.n330 fout1.n329 0.009
R9614 fout1.n239 fout1.n235 0.007
R9615 fout1.n346 fout1.n345 0.007
R9616 fout1.n352 fout1.n351 0.007
R9617 fout1.n444 fout1.n443 0.007
R9618 fout1.n472 fout1.n471 0.007
R9619 fout1.n203 fout1.n202 0.007
R9620 fout1.n328 fout1.n324 0.007
R9621 fout1.n333 fout1.n332 0.007
R9622 fout1.n335 fout1.n334 0.007
R9623 fout1.n488 fout1.n487 0.007
R9624 fout1.n479 fout1.n478 0.007
R9625 fout1.n518 fout1.n517 0.006
R9626 fout1.n503 fout1.n502 0.006
R9627 fout1.n512 fout1.n511 0.006
R9628 fout1.n188 fout1.n187 0.006
R9629 fout1.n190 fout1.n189 0.006
R9630 fout1.n195 fout1.n194 0.006
R9631 fout1.n197 fout1.n196 0.006
R9632 fout1.n312 fout1.n311 0.006
R9633 fout1.n314 fout1.n313 0.006
R9634 fout1.n319 fout1.n318 0.006
R9635 fout1.n321 fout1.n320 0.006
R9636 fout1.n401 fout1.n400 0.006
R9637 fout1.n403 fout1.n402 0.006
R9638 fout1.n408 fout1.n407 0.006
R9639 fout1.n410 fout1.n409 0.006
R9640 fout1.n495 fout1.n494 0.006
R9641 fout1.n128 fout1.n121 0.006
R9642 fout1.n127 fout1.n126 0.006
R9643 fout1.n103 fout1.n102 0.006
R9644 fout1.n59 fout1.n58 0.006
R9645 fout1.n74 fout1.n73 0.006
R9646 fout1.n83 fout1.n82 0.006
R9647 fout1.n40 fout1.n33 0.006
R9648 fout1.n39 fout1.n38 0.006
R9649 fout1.n16 fout1.n15 0.006
R9650 fout1.n158 fout1.n157 0.005
R9651 fout1.n160 fout1.n159 0.005
R9652 fout1.n215 fout1.n211 0.005
R9653 fout1.n219 fout1.n217 0.005
R9654 fout1.n291 fout1.n286 0.005
R9655 fout1.n284 fout1.n283 0.005
R9656 fout1.n256 fout1.n255 0.005
R9657 fout1.n356 fout1.n355 0.005
R9658 fout1.n431 fout1.n430 0.005
R9659 fout1.n451 fout1.n450 0.005
R9660 fout1.n376 fout1.n375 0.005
R9661 fout1.n420 fout1.n419 0.005
R9662 fout1.n540 fout1.n539 0.004
R9663 fout1.n11 fout1.n1 0.004
R9664 fout1.n54 fout1.n44 0.004
R9665 fout1.n513 fout1.n498 0.003
R9666 fout1.n42 fout1.n41 0.003
R9667 fout1.n85 fout1.n84 0.003
R9668 fout1.n98 fout1.n88 0.003
R9669 fout1.n130 fout1.n129 0.003
R9670 fout1.n172 fout1.n166 0.003
R9671 fout1.n364 fout1.n360 0.003
R9672 fout1.n385 fout1.n382 0.003
R9673 fout1.n374 fout1.n371 0.003
R9674 fout1.n450 fout1.n446 0.003
R9675 fout1.n466 fout1.n464 0.003
R9676 fout1.n476 fout1.n475 0.003
R9677 fout1.n485 fout1.n484 0.003
R9678 fout1.n295 fout1.n294 0.003
R9679 fout1.n425 fout1.n424 0.003
R9680 fout1.n527 fout1.n519 0.003
R9681 fout1.n67 fout1.n60 0.003
R9682 fout1.n112 fout1.n104 0.003
R9683 fout1.n25 fout1.n17 0.003
R9684 fout1.n539 fout1.n528 0.002
R9685 fout1.n68 fout1.n54 0.002
R9686 fout1.n26 fout1.n11 0.002
R9687 fout1.n528 fout1.n513 0.002
R9688 fout1.n84 fout1.n68 0.002
R9689 fout1.n129 fout1.n113 0.002
R9690 fout1.n113 fout1.n98 0.002
R9691 fout1.n41 fout1.n26 0.002
R9692 fout1.n227 fout1.n223 0.001
R9693 fout1.n231 fout1.n229 0.001
R9694 fout1.n234 fout1.n233 0.001
R9695 fout1.n240 fout1.n239 0.001
R9696 fout1.n277 fout1.n274 0.001
R9697 fout1.n272 fout1.n271 0.001
R9698 fout1.n266 fout1.n263 0.001
R9699 fout1.n260 fout1.n259 0.001
R9700 fout1.n351 fout1.n347 0.001
R9701 fout1.n357 fout1.n356 0.001
R9702 fout1.n436 fout1.n431 0.001
R9703 fout1.n178 fout1.n177 0.001
R9704 fout1.n201 fout1.n200 0.001
R9705 fout1.n337 fout1.n336 0.001
R9706 fout1.n340 fout1.n339 0.001
R9707 fout1.n413 fout1.n412 0.001
R9708 fout1.n87 fout1.n0 0.001
R9709 a_n6002_2899.n33 a_n6002_2899.t2 733.436
R9710 a_n6002_2899.n53 a_n6002_2899.t5 733.436
R9711 a_n6002_2899.n24 a_n6002_2899.t4 399.248
R9712 a_n6002_2899.n44 a_n6002_2899.t3 399.248
R9713 a_n6002_2899.n95 a_n6002_2899.n94 92.5
R9714 a_n6002_2899.n12 a_n6002_2899.n11 92.5
R9715 a_n6002_2899.n94 a_n6002_2899.t0 70.344
R9716 a_n6002_2899.n89 a_n6002_2899.n88 31.034
R9717 a_n6002_2899.n68 a_n6002_2899.n67 31.034
R9718 a_n6002_2899.n71 a_n6002_2899.n72 9.3
R9719 a_n6002_2899.n82 a_n6002_2899.n83 9.3
R9720 a_n6002_2899.n90 a_n6002_2899.n89 9.3
R9721 a_n6002_2899.n69 a_n6002_2899.n68 9.3
R9722 a_n6002_2899.n162 a_n6002_2899.n155 9.154
R9723 a_n6002_2899.n162 a_n6002_2899.n113 9.143
R9724 a_n6002_2899.n162 a_n6002_2899.n120 9.143
R9725 a_n6002_2899.n162 a_n6002_2899.n126 9.132
R9726 a_n6002_2899.n162 a_n6002_2899.n106 9.132
R9727 a_n6002_2899.n162 a_n6002_2899.n159 8.885
R9728 a_n6002_2899.n162 a_n6002_2899.n130 8.885
R9729 a_n6002_2899.n162 a_n6002_2899.n134 8.875
R9730 a_n6002_2899.n162 a_n6002_2899.n100 8.875
R9731 a_n6002_2899.n162 a_n6002_2899.n161 8.864
R9732 a_n6002_2899.n162 a_n6002_2899.n136 8.864
R9733 a_n6002_2899.n96 a_n6002_2899.n95 8.282
R9734 a_n6002_2899.n13 a_n6002_2899.n12 8.282
R9735 a_n6002_2899.t1 a_n6002_2899.n162 7.141
R9736 a_n6002_2899.n59 a_n6002_2899.n58 6.379
R9737 a_n6002_2899.n90 a_n6002_2899.n86 5.647
R9738 a_n6002_2899.n69 a_n6002_2899.n65 5.647
R9739 a_n6002_2899.n16 a_n6002_2899.n15 4.65
R9740 a_n6002_2899.n155 a_n6002_2899.n5 4.65
R9741 a_n6002_2899.n155 a_n6002_2899.n138 4.517
R9742 a_n6002_2899.n14 a_n6002_2899.n13 4.5
R9743 a_n6002_2899.n17 a_n6002_2899.n10 4.5
R9744 a_n6002_2899.n9 a_n6002_2899.n96 4.5
R9745 a_n6002_2899.n84 a_n6002_2899.n92 4.5
R9746 a_n6002_2899.n18 a_n6002_2899.n81 4.5
R9747 a_n6002_2899.n61 a_n6002_2899.n76 4.5
R9748 a_n6002_2899.n157 a_n6002_2899.n156 4.141
R9749 a_n6002_2899.n155 a_n6002_2899.n137 4.141
R9750 a_n6002_2899.n128 a_n6002_2899.n127 4.141
R9751 a_n6002_2899.n88 a_n6002_2899.n87 4.137
R9752 a_n6002_2899.n67 a_n6002_2899.n66 4.137
R9753 a_n6002_2899.n81 a_n6002_2899.n79 3.764
R9754 a_n6002_2899.n70 a_n6002_2899.n63 3.764
R9755 a_n6002_2899.n102 a_n6002_2899.n101 3.764
R9756 a_n6002_2899.n116 a_n6002_2899.n115 3.764
R9757 a_n6002_2899.n106 a_n6002_2899.n105 3.736
R9758 a_n6002_2899.n92 a_n6002_2899.n91 3.388
R9759 a_n6002_2899.n76 a_n6002_2899.n75 3.388
R9760 a_n6002_2899.n98 a_n6002_2899.n97 3.388
R9761 a_n6002_2899.n112 a_n6002_2899.n111 3.388
R9762 a_n6002_2899.n124 a_n6002_2899.n123 3.388
R9763 a_n6002_2899.n132 a_n6002_2899.n131 3.388
R9764 a_n6002_2899.n126 a_n6002_2899.n122 3.36
R9765 a_n6002_2899.n92 a_n6002_2899.n90 3.011
R9766 a_n6002_2899.n96 a_n6002_2899.n93 3.011
R9767 a_n6002_2899.n76 a_n6002_2899.n74 3.011
R9768 a_n6002_2899.n99 a_n6002_2899.n98 3.011
R9769 a_n6002_2899.n111 a_n6002_2899.n110 3.011
R9770 a_n6002_2899.n109 a_n6002_2899.n108 3.011
R9771 a_n6002_2899.n122 a_n6002_2899.n121 3.011
R9772 a_n6002_2899.n125 a_n6002_2899.n124 3.011
R9773 a_n6002_2899.n133 a_n6002_2899.n132 3.011
R9774 a_n6002_2899.n139 a_n6002_2899.n58 2.921
R9775 a_n6002_2899.n81 a_n6002_2899.n80 2.635
R9776 a_n6002_2899.n70 a_n6002_2899.n69 2.635
R9777 a_n6002_2899.n103 a_n6002_2899.n102 2.635
R9778 a_n6002_2899.n105 a_n6002_2899.n104 2.635
R9779 a_n6002_2899.n119 a_n6002_2899.n118 2.635
R9780 a_n6002_2899.n115 a_n6002_2899.n114 2.635
R9781 a_n6002_2899.n60 a_n6002_2899.n59 2.632
R9782 a_n6002_2899.n158 a_n6002_2899.n157 2.258
R9783 a_n6002_2899.n129 a_n6002_2899.n128 2.258
R9784 a_n6002_2899.n113 a_n6002_2899.n109 2.245
R9785 a_n6002_2899.n120 a_n6002_2899.n119 2.245
R9786 a_n6002_2899.n151 a_n6002_2899.n150 1.633
R9787 a_n6002_2899.n147 a_n6002_2899.n146 1.619
R9788 a_n6002_2899.n149 a_n6002_2899.n164 1.594
R9789 a_n6002_2899.n140 a_n6002_2899.n143 1.588
R9790 a_n6002_2899.n151 a_n6002_2899.n163 1.587
R9791 a_n6002_2899.n118 a_n6002_2899.n117 1.505
R9792 a_n6002_2899.n18 a_n6002_2899.n78 1.5
R9793 a_n6002_2899.n4 a_n6002_2899.n6 1.5
R9794 a_n6002_2899.n141 a_n6002_2899.n153 1.5
R9795 a_n6002_2899.n34 a_n6002_2899.n33 2.49
R9796 a_n6002_2899.n54 a_n6002_2899.n53 2.49
R9797 a_n6002_2899.n22 a_n6002_2899.n28 1.137
R9798 a_n6002_2899.n25 a_n6002_2899.n26 1.137
R9799 a_n6002_2899.n41 a_n6002_2899.n48 1.137
R9800 a_n6002_2899.n45 a_n6002_2899.n46 1.137
R9801 a_n6002_2899.n3 a_n6002_2899.n36 1.136
R9802 a_n6002_2899.n0 a_n6002_2899.n42 1.136
R9803 a_n6002_2899.n1 a_n6002_2899.n56 1.136
R9804 a_n6002_2899.n108 a_n6002_2899.n107 1.129
R9805 a_n6002_2899.n86 a_n6002_2899.n85 0.752
R9806 a_n6002_2899.n65 a_n6002_2899.n64 0.752
R9807 a_n6002_2899.n161 a_n6002_2899.n160 0.155
R9808 a_n6002_2899.n136 a_n6002_2899.n135 0.155
R9809 a_n6002_2899.n100 a_n6002_2899.n99 0.144
R9810 a_n6002_2899.n134 a_n6002_2899.n133 0.144
R9811 a_n6002_2899.n159 a_n6002_2899.n158 0.132
R9812 a_n6002_2899.n130 a_n6002_2899.n129 0.132
R9813 a_n6002_2899.n149 a_n6002_2899.n148 0.127
R9814 a_n6002_2899.n147 a_n6002_2899.n145 0.119
R9815 a_n6002_2899.n140 a_n6002_2899.n142 0.111
R9816 a_n6002_2899.n4 a_n6002_2899.n5 0.103
R9817 a_n6002_2899.n33 a_n6002_2899.n32 0.126
R9818 a_n6002_2899.n53 a_n6002_2899.n52 0.126
R9819 a_n6002_2899.n20 a_n6002_2899.n19 0.064
R9820 a_n6002_2899.n31 a_n6002_2899.n30 0.064
R9821 a_n6002_2899.n39 a_n6002_2899.n38 0.064
R9822 a_n6002_2899.n51 a_n6002_2899.n50 0.064
R9823 a_n6002_2899.n139 a_n6002_2899.n141 0.083
R9824 a_n6002_2899.n141 a_n6002_2899.n140 0.042
R9825 a_n6002_2899.n163 a_n6002_2899.n168 0.037
R9826 a_n6002_2899.n150 a_n6002_2899.n152 0.034
R9827 a_n6002_2899.n28 a_n6002_2899.n29 0.032
R9828 a_n6002_2899.n35 a_n6002_2899.n37 0.032
R9829 a_n6002_2899.n48 a_n6002_2899.n49 0.032
R9830 a_n6002_2899.n55 a_n6002_2899.n57 0.032
R9831 a_n6002_2899.n84 a_n6002_2899.n82 0.094
R9832 a_n6002_2899.n21 a_n6002_2899.n20 0.028
R9833 a_n6002_2899.n32 a_n6002_2899.n31 0.028
R9834 a_n6002_2899.n40 a_n6002_2899.n39 0.028
R9835 a_n6002_2899.n52 a_n6002_2899.n51 0.028
R9836 a_n6002_2899.n78 a_n6002_2899.n77 0.293
R9837 a_n6002_2899.n78 a_n6002_2899.n62 0.877
R9838 a_n6002_2899.n143 a_n6002_2899.n144 0.024
R9839 a_n6002_2899.n164 a_n6002_2899.n169 0.024
R9840 a_n6002_2899.n106 a_n6002_2899.n103 0.024
R9841 a_n6002_2899.n126 a_n6002_2899.n125 0.024
R9842 a_n6002_2899.n5 a_n6002_2899.n139 0.022
R9843 a_n6002_2899.n16 a_n6002_2899.n14 0.022
R9844 a_n6002_2899.n17 a_n6002_2899.n16 0.02
R9845 a_n6002_2899.n62 a_n6002_2899.n60 0.019
R9846 a_n6002_2899.n62 a_n6002_2899.n61 2.433
R9847 a_n6002_2899.n9 a_n6002_2899.n84 0.044
R9848 a_n6002_2899.n61 a_n6002_2899.n71 0.032
R9849 a_n6002_2899.n82 a_n6002_2899.n18 0.031
R9850 a_n6002_2899.n61 a_n6002_2899.n73 0.017
R9851 a_n6002_2899.n26 a_n6002_2899.n27 0.017
R9852 a_n6002_2899.n46 a_n6002_2899.n47 0.017
R9853 a_n6002_2899.n166 a_n6002_2899.n165 0.016
R9854 a_n6002_2899.n71 a_n6002_2899.n70 4.595
R9855 a_n6002_2899.n56 a_n6002_2899.n55 1.181
R9856 a_n6002_2899.n42 a_n6002_2899.n41 0.044
R9857 a_n6002_2899.n41 a_n6002_2899.n43 0.04
R9858 a_n6002_2899.n45 a_n6002_2899.n44 0.02
R9859 a_n6002_2899.n6 a_n6002_2899.n7 0.013
R9860 a_n6002_2899.n142 a_n6002_2899.n147 0.013
R9861 a_n6002_2899.n120 a_n6002_2899.n116 0.012
R9862 a_n6002_2899.n113 a_n6002_2899.n112 0.012
R9863 a_n6002_2899.n8 a_n6002_2899.n17 0.011
R9864 a_n6002_2899.n153 a_n6002_2899.n154 0.011
R9865 a_n6002_2899.n23 a_n6002_2899.n25 0.01
R9866 a_n6002_2899.n43 a_n6002_2899.n45 0.01
R9867 a_n6002_2899.n169 a_n6002_2899.n167 0.009
R9868 a_n6002_2899.n2 a_n6002_2899.n21 2.621
R9869 a_n6002_2899.n36 a_n6002_2899.n34 0.006
R9870 a_n6002_2899.n42 a_n6002_2899.n40 2.621
R9871 a_n6002_2899.n36 a_n6002_2899.n35 1.181
R9872 a_n6002_2899.n2 a_n6002_2899.n22 0.044
R9873 a_n6002_2899.n22 a_n6002_2899.n23 0.04
R9874 a_n6002_2899.n25 a_n6002_2899.n24 0.02
R9875 a_n6002_2899.n56 a_n6002_2899.n54 0.006
R9876 a_n6002_2899.n145 a_n6002_2899.n149 0.005
R9877 a_n6002_2899.n148 a_n6002_2899.n151 0.005
R9878 a_n6002_2899.n3 a_n6002_2899.n2 1.245
R9879 a_n6002_2899.n4 a_n6002_2899.n166 2.057
R9880 a_n6002_2899.n0 a_n6002_2899.n3 0.11
R9881 a_n6002_2899.n1 a_n6002_2899.n0 0.109
R9882 a_n6002_2899.n59 a_n6002_2899.n1 0.072
R9883 a_n6002_2899.n9 a_n6002_2899.n8 0.07
R9884 fout4.n510 fout4.t10 1038.92
R9885 fout4.n388 fout4.t5 1037.29
R9886 fout4.n389 fout4.t4 797.225
R9887 fout4.n525 fout4.t6 795.549
R9888 fout4.n367 fout4.t11 732.331
R9889 fout4.n479 fout4.t13 731.671
R9890 fout4.n417 fout4.t14 731.671
R9891 fout4.n497 fout4.t8 730.671
R9892 fout4.n453 fout4.t3 400.618
R9893 fout4.n496 fout4.t7 400.599
R9894 fout4.n11 fout4.t12 397.315
R9895 fout4.n497 fout4.t9 395.839
R9896 fout4.n244 fout4.n243 13.176
R9897 fout4.n14 fout4.t0 11.722
R9898 fout4.n14 fout4.t2 10.994
R9899 fout4.n23 fout4.n22 9.3
R9900 fout4.n322 fout4.n321 9.3
R9901 fout4.n288 fout4.n287 9.3
R9902 fout4.n285 fout4.n284 9.3
R9903 fout4.n222 fout4.n221 9.3
R9904 fout4.n336 fout4.n335 9.3
R9905 fout4.n338 fout4.n337 9.3
R9906 fout4.n220 fout4.n219 9.3
R9907 fout4.n253 fout4.n252 9.3
R9908 fout4.n266 fout4.n265 9.3
R9909 fout4.n274 fout4.n273 9.3
R9910 fout4.n277 fout4.n276 9.3
R9911 fout4.n137 fout4.n136 9.3
R9912 fout4.n134 fout4.n133 9.3
R9913 fout4.n50 fout4.n49 9.3
R9914 fout4.n48 fout4.n47 9.3
R9915 fout4.n41 fout4.n40 8.097
R9916 fout4.n276 fout4.n275 5.457
R9917 fout4.n136 fout4.n135 5.08
R9918 fout4.n39 fout4.n38 4.65
R9919 fout4.n146 fout4.n145 4.65
R9920 fout4.n55 fout4.n53 4.5
R9921 fout4.n107 fout4.n103 4.5
R9922 fout4.n111 fout4.n100 4.5
R9923 fout4.n126 fout4.n125 4.5
R9924 fout4.n81 fout4.n80 4.5
R9925 fout4.n255 fout4.n247 4.5
R9926 fout4.n262 fout4.n245 4.5
R9927 fout4.n271 fout4.n242 4.5
R9928 fout4.n294 fout4.n293 4.5
R9929 fout4.n342 fout4.n341 4.5
R9930 fout4.n330 fout4.n329 4.5
R9931 fout4.n230 fout4.n229 4.5
R9932 fout4.n237 fout4.n236 4.5
R9933 fout4.n302 fout4.n301 4.5
R9934 fout4.n282 fout4.n281 4.5
R9935 fout4.n119 fout4.n118 4.5
R9936 fout4.n213 fout4.n212 4.5
R9937 fout4.n27 fout4.n25 4.5
R9938 fout4.n229 fout4.n227 4.314
R9939 fout4.n301 fout4.n298 3.944
R9940 fout4.n103 fout4.n102 3.937
R9941 fout4.n118 fout4.n117 3.567
R9942 fout4.n147 fout4.n140 3.033
R9943 fout4.n43 fout4.n42 3.033
R9944 fout4.n40 fout4.t1 2.9
R9945 fout4.n300 fout4.n299 2.258
R9946 fout4.n116 fout4.n115 2.258
R9947 fout4.n235 fout4.n234 1.882
R9948 fout4.n236 fout4.n235 1.882
R9949 fout4.n99 fout4.n98 1.882
R9950 fout4.n350 fout4.n14 1.519
R9951 fout4.n118 fout4.n116 1.505
R9952 fout4.n100 fout4.n99 1.505
R9953 fout4.n56 fout4.n55 1.5
R9954 fout4.n343 fout4.n342 1.5
R9955 fout4.n82 fout4.n81 1.5
R9956 fout4.n148 fout4.n147 1.5
R9957 fout4.n127 fout4.n126 1.5
R9958 fout4.n214 fout4.n213 1.5
R9959 fout4.n28 fout4.n27 1.5
R9960 fout4.n465 fout4.n464 1.435
R9961 fout4.n448 fout4.n447 1.435
R9962 fout4.n402 fout4.n388 1.388
R9963 fout4.n527 fout4.n525 1.355
R9964 fout4.n511 fout4.n510 1.355
R9965 fout4.n390 fout4.n389 1.354
R9966 fout4.n419 fout4.n417 1.354
R9967 fout4.n369 fout4.n367 1.354
R9968 fout4.n481 fout4.n479 1.354
R9969 fout4.n12 fout4.n11 1.354
R9970 fout4.n528 fout4.n527 1.142
R9971 fout4.n482 fout4.n481 1.142
R9972 fout4.n13 fout4.n12 1.142
R9973 fout4.n420 fout4.n419 1.14
R9974 fout4.n529 fout4.n528 1.138
R9975 fout4.n483 fout4.n482 1.138
R9976 fout4.n362 fout4.n13 1.138
R9977 fout4.n512 fout4.n511 1.137
R9978 fout4.n538 fout4.n537 1.137
R9979 fout4.n503 fout4.n502 1.137
R9980 fout4.n534 fout4.n533 1.137
R9981 fout4.n518 fout4.n517 1.137
R9982 fout4.n466 fout4.n465 1.137
R9983 fout4.n492 fout4.n491 1.137
R9984 fout4.n458 fout4.n457 1.137
R9985 fout4.n488 fout4.n487 1.137
R9986 fout4.n472 fout4.n471 1.137
R9987 fout4.n449 fout4.n448 1.137
R9988 fout4.n440 fout4.n439 1.137
R9989 fout4.n425 fout4.n424 1.137
R9990 fout4.n430 fout4.n429 1.137
R9991 fout4.n434 fout4.n433 1.137
R9992 fout4.n359 fout4.n358 1.137
R9993 fout4.n375 fout4.n374 1.137
R9994 fout4.n354 fout4.n353 1.137
R9995 fout4.n3 fout4.n2 1.137
R9996 fout4.n370 fout4.n369 1.137
R9997 fout4.n540 fout4.n539 1.136
R9998 fout4.n494 fout4.n493 1.136
R9999 fout4.n468 fout4.n467 1.136
R10000 fout4.n514 fout4.n513 1.136
R10001 fout4.n451 fout4.n450 1.136
R10002 fout4.n378 fout4.n377 1.136
R10003 fout4.n361 fout4.n360 1.136
R10004 fout4.n341 fout4.n340 1.129
R10005 fout4.n301 fout4.n300 1.129
R10006 fout4.n293 fout4.n292 1.129
R10007 fout4.n303 fout4.n302 1.042
R10008 fout4.n345 fout4.n344 0.853
R10009 fout4.n192 fout4.n191 0.853
R10010 fout4.n150 fout4.n149 0.853
R10011 fout4.n58 fout4.n57 0.853
R10012 fout4.n410 fout4.n409 0.826
R10013 fout4.n212 fout4.n211 0.752
R10014 fout4.n80 fout4.n79 0.752
R10015 fout4.n125 fout4.n124 0.752
R10016 fout4.n103 fout4.n101 0.752
R10017 fout4.n53 fout4.n52 0.752
R10018 fout4.n25 fout4.n24 0.752
R10019 fout4.n30 fout4.n29 0.716
R10020 fout4.n350 fout4.n349 0.689
R10021 fout4.n351 fout4.n350 0.68
R10022 fout4.n252 fout4.n251 0.536
R10023 fout4.n265 fout4.n264 0.536
R10024 fout4.n145 fout4.n144 0.476
R10025 fout4.n287 fout4.n286 0.475
R10026 fout4.n410 fout4.n379 0.471
R10027 fout4.n403 fout4.n402 0.44
R10028 fout4.n42 fout4.n41 0.382
R10029 fout4.n328 fout4.n327 0.382
R10030 fout4.n329 fout4.n328 0.376
R10031 fout4.n229 fout4.n228 0.376
R10032 fout4.n281 fout4.n280 0.376
R10033 fout4.n242 fout4.n241 0.376
R10034 fout4.n245 fout4.n244 0.376
R10035 fout4.n247 fout4.n246 0.376
R10036 fout4.n52 fout4.n51 0.35
R10037 fout4.n340 fout4.n339 0.349
R10038 fout4 fout4.n541 0.165
R10039 fout4.n499 fout4.n498 0.152
R10040 fout4.n496 fout4.n495 0.123
R10041 fout4.n453 fout4.n452 0.123
R10042 fout4 fout4.n410 0.107
R10043 fout4.n454 fout4.n453 0.091
R10044 fout4.n479 fout4.n478 0.083
R10045 fout4.n417 fout4.n416 0.083
R10046 fout4.n367 fout4.n366 0.083
R10047 fout4.n11 fout4.n10 0.083
R10048 fout4.n388 fout4.n387 0.076
R10049 fout4.n525 fout4.n524 0.075
R10050 fout4.n510 fout4.n509 0.075
R10051 fout4.n498 fout4.n496 0.07
R10052 fout4.n444 fout4.n443 0.064
R10053 fout4.n384 fout4.n383 0.059
R10054 fout4.n324 fout4.n323 0.047
R10055 fout4.n278 fout4.n277 0.047
R10056 fout4.n268 fout4.n267 0.047
R10057 fout4.n259 fout4.n258 0.047
R10058 fout4.n249 fout4.n248 0.047
R10059 fout4.n138 fout4.n137 0.047
R10060 fout4.n21 fout4.n20 0.047
R10061 fout4.n106 fout4.n105 0.043
R10062 fout4.n88 fout4.n87 0.043
R10063 fout4.n226 fout4.n225 0.041
R10064 fout4.n311 fout4.n310 0.041
R10065 fout4.n45 fout4.n44 0.035
R10066 fout4.n181 fout4.n180 0.035
R10067 fout4.n176 fout4.n175 0.035
R10068 fout4.n35 fout4.n34 0.035
R10069 fout4.n333 fout4.n332 0.034
R10070 fout4.n261 fout4.n260 0.034
R10071 fout4.n257 fout4.n256 0.034
R10072 fout4.n48 fout4.n46 0.034
R10073 fout4.n320 fout4.n319 0.034
R10074 fout4.n318 fout4.n317 0.034
R10075 fout4.n170 fout4.n169 0.034
R10076 fout4.n189 fout4.n188 0.034
R10077 fout4.n82 fout4.n75 0.034
R10078 fout4.n84 fout4.n83 0.034
R10079 fout4.n132 fout4.n131 0.034
R10080 fout4.n37 fout4.n36 0.034
R10081 fout4.n533 fout4.n532 0.032
R10082 fout4.n487 fout4.n486 0.032
R10083 fout4.n433 fout4.n432 0.032
R10084 fout4.n336 fout4.n334 0.032
R10085 fout4.n147 fout4.n146 0.032
R10086 fout4.n43 fout4.n39 0.032
R10087 fout4.n187 fout4.n186 0.032
R10088 fout4.n56 fout4.n37 0.032
R10089 fout4.n358 fout4.n356 0.032
R10090 fout4.n397 fout4.n396 0.032
R10091 fout4.n398 fout4.n397 0.032
R10092 fout4.n402 fout4.n401 0.032
R10093 fout4.n347 fout4.n346 0.031
R10094 fout4.n205 fout4.n204 0.031
R10095 fout4.n194 fout4.n193 0.031
R10096 fout4.n163 fout4.n162 0.031
R10097 fout4.n152 fout4.n151 0.031
R10098 fout4.n71 fout4.n70 0.031
R10099 fout4.n60 fout4.n59 0.031
R10100 fout4.n285 fout4.n283 0.03
R10101 fout4.n270 fout4.n269 0.03
R10102 fout4.n77 fout4.n76 0.03
R10103 fout4.n20 fout4.n19 0.03
R10104 fout4.n343 fout4.n320 0.03
R10105 fout4.n315 fout4.n314 0.03
R10106 fout4.n185 fout4.n184 0.03
R10107 fout4.n73 fout4.n72 0.03
R10108 fout4.n85 fout4.n84 0.03
R10109 fout4.n32 fout4.n31 0.03
R10110 fout4.n392 fout4.n391 0.03
R10111 fout4.n517 fout4.n516 0.028
R10112 fout4.n533 fout4.n531 0.028
R10113 fout4.n537 fout4.n536 0.028
R10114 fout4.n502 fout4.n500 0.028
R10115 fout4.n478 fout4.n477 0.028
R10116 fout4.n476 fout4.n475 0.028
R10117 fout4.n462 fout4.n461 0.028
R10118 fout4.n464 fout4.n463 0.028
R10119 fout4.n471 fout4.n470 0.028
R10120 fout4.n487 fout4.n485 0.028
R10121 fout4.n491 fout4.n490 0.028
R10122 fout4.n457 fout4.n455 0.028
R10123 fout4.n416 fout4.n415 0.028
R10124 fout4.n445 fout4.n444 0.028
R10125 fout4.n447 fout4.n446 0.028
R10126 fout4.n429 fout4.n428 0.028
R10127 fout4.n439 fout4.n437 0.028
R10128 fout4.n325 fout4.n324 0.028
R10129 fout4.n224 fout4.n223 0.028
R10130 fout4.n239 fout4.n238 0.028
R10131 fout4.n302 fout4.n240 0.028
R10132 fout4.n291 fout4.n290 0.028
R10133 fout4.n147 fout4.n139 0.028
R10134 fout4.n113 fout4.n112 0.028
R10135 fout4.n105 fout4.n104 0.028
R10136 fout4.n55 fout4.n50 0.028
R10137 fout4.n27 fout4.n23 0.028
R10138 fout4.n215 fout4.n214 0.028
R10139 fout4.n344 fout4.n218 0.028
R10140 fout4.n313 fout4.n312 0.028
R10141 fout4.n306 fout4.n305 0.028
R10142 fout4.n304 fout4.n303 0.028
R10143 fout4.n168 fout4.n167 0.028
R10144 fout4.n190 fout4.n189 0.028
R10145 fout4.n183 fout4.n182 0.028
R10146 fout4.n174 fout4.n173 0.028
R10147 fout4.n149 fout4.n148 0.028
R10148 fout4.n93 fout4.n92 0.028
R10149 fout4.n87 fout4.n86 0.028
R10150 fout4.n28 fout4.n18 0.028
R10151 fout4.n366 fout4.n365 0.028
R10152 fout4.n364 fout4.n363 0.028
R10153 fout4.n8 fout4.n7 0.028
R10154 fout4.n10 fout4.n9 0.028
R10155 fout4.n374 fout4.n373 0.028
R10156 fout4.n353 fout4.n352 0.028
R10157 fout4.n358 fout4.n357 0.028
R10158 fout4.n2 fout4.n0 0.028
R10159 fout4.n394 fout4.n393 0.028
R10160 fout4.n396 fout4.n395 0.028
R10161 fout4.n399 fout4.n398 0.028
R10162 fout4.n401 fout4.n400 0.028
R10163 fout4.n201 fout4.n200 0.027
R10164 fout4.n198 fout4.n197 0.027
R10165 fout4.n159 fout4.n158 0.027
R10166 fout4.n156 fout4.n155 0.027
R10167 fout4.n67 fout4.n66 0.027
R10168 fout4.n64 fout4.n63 0.027
R10169 fout4.n342 fout4.n338 0.026
R10170 fout4.n282 fout4.n279 0.026
R10171 fout4.n142 fout4.n141 0.026
R10172 fout4.n119 fout4.n114 0.026
R10173 fout4.n165 fout4.n164 0.026
R10174 fout4.n191 fout4.n171 0.026
R10175 fout4.n130 fout4.n129 0.026
R10176 fout4.n95 fout4.n94 0.026
R10177 fout4.n90 fout4.n89 0.026
R10178 fout4.n17 fout4.n16 0.026
R10179 fout4.n381 fout4.n380 0.026
R10180 fout4.n383 fout4.n382 0.026
R10181 fout4.n385 fout4.n384 0.026
R10182 fout4.n387 fout4.n386 0.026
R10183 fout4.n524 fout4.n523 0.025
R10184 fout4.n522 fout4.n521 0.025
R10185 fout4.n507 fout4.n506 0.025
R10186 fout4.n509 fout4.n508 0.025
R10187 fout4.n29 fout4.n28 0.024
R10188 fout4.n289 fout4.n288 0.024
R10189 fout4.n146 fout4.n143 0.024
R10190 fout4.n217 fout4.n216 0.024
R10191 fout4.n309 fout4.n308 0.024
R10192 fout4.n171 fout4.n170 0.024
R10193 fout4.n178 fout4.n177 0.024
R10194 fout4.n127 fout4.n97 0.024
R10195 fout4.n406 fout4.n405 0.023
R10196 fout4.n232 fout4.n231 0.022
R10197 fout4.n279 fout4.n278 0.022
R10198 fout4.n266 fout4.n263 0.022
R10199 fout4.n254 fout4.n253 0.022
R10200 fout4.n143 fout4.n142 0.022
R10201 fout4.n109 fout4.n108 0.022
R10202 fout4.n218 fout4.n217 0.022
R10203 fout4.n191 fout4.n190 0.022
R10204 fout4.n179 fout4.n178 0.022
R10205 fout4.n148 fout4.n132 0.022
R10206 fout4.n131 fout4.n130 0.022
R10207 fout4.n296 fout4.n295 0.02
R10208 fout4.n294 fout4.n291 0.02
R10209 fout4.n290 fout4.n289 0.02
R10210 fout4.n139 fout4.n138 0.02
R10211 fout4.n123 fout4.n122 0.02
R10212 fout4.n214 fout4.n208 0.02
R10213 fout4.n344 fout4.n343 0.02
R10214 fout4.n169 fout4.n168 0.02
R10215 fout4.n149 fout4.n85 0.02
R10216 fout4.n16 fout4.n15 0.02
R10217 fout4.n346 fout4.n345 0.019
R10218 fout4.n345 fout4.n205 0.019
R10219 fout4.n193 fout4.n192 0.019
R10220 fout4.n192 fout4.n163 0.019
R10221 fout4.n151 fout4.n150 0.019
R10222 fout4.n150 fout4.n71 0.019
R10223 fout4.n59 fout4.n58 0.019
R10224 fout4.n58 fout4.n30 0.019
R10225 fout4.n308 fout4.n307 0.018
R10226 fout4.n57 fout4.n56 0.018
R10227 fout4.n527 fout4.n526 0.017
R10228 fout4.n517 fout4.n515 0.017
R10229 fout4.n502 fout4.n501 0.017
R10230 fout4.n511 fout4.n505 0.017
R10231 fout4.n481 fout4.n480 0.017
R10232 fout4.n471 fout4.n469 0.017
R10233 fout4.n457 fout4.n456 0.017
R10234 fout4.n465 fout4.n460 0.017
R10235 fout4.n419 fout4.n418 0.017
R10236 fout4.n424 fout4.n423 0.017
R10237 fout4.n439 fout4.n438 0.017
R10238 fout4.n448 fout4.n442 0.017
R10239 fout4.n210 fout4.n209 0.017
R10240 fout4.n223 fout4.n222 0.017
R10241 fout4.n272 fout4.n271 0.017
R10242 fout4.n269 fout4.n268 0.017
R10243 fout4.n208 fout4.n207 0.017
R10244 fout4.n314 fout4.n313 0.017
R10245 fout4.n167 fout4.n166 0.017
R10246 fout4.n188 fout4.n187 0.017
R10247 fout4.n186 fout4.n185 0.017
R10248 fout4.n184 fout4.n183 0.017
R10249 fout4.n129 fout4.n128 0.017
R10250 fout4.n97 fout4.n96 0.017
R10251 fout4.n91 fout4.n90 0.017
R10252 fout4.n369 fout4.n368 0.017
R10253 fout4.n374 fout4.n372 0.017
R10254 fout4.n2 fout4.n1 0.017
R10255 fout4.n12 fout4.n6 0.017
R10256 fout4.n391 fout4.n390 0.017
R10257 fout4.n393 fout4.n392 0.017
R10258 fout4.n534 fout4.n530 0.016
R10259 fout4.n538 fout4.n535 0.016
R10260 fout4.n488 fout4.n484 0.016
R10261 fout4.n492 fout4.n489 0.016
R10262 fout4.n430 fout4.n426 0.016
R10263 fout4.n435 fout4.n434 0.016
R10264 fout4.n359 fout4.n355 0.016
R10265 fout4.n477 fout4.n476 0.015
R10266 fout4.n463 fout4.n462 0.015
R10267 fout4.n415 fout4.n414 0.015
R10268 fout4.n446 fout4.n445 0.015
R10269 fout4.n428 fout4.n427 0.015
R10270 fout4.n437 fout4.n436 0.015
R10271 fout4.n326 fout4.n325 0.015
R10272 fout4.n334 fout4.n333 0.015
R10273 fout4.n240 fout4.n239 0.015
R10274 fout4.n81 fout4.n78 0.015
R10275 fout4.n114 fout4.n113 0.015
R10276 fout4.n112 fout4.n111 0.015
R10277 fout4.n319 fout4.n318 0.015
R10278 fout4.n317 fout4.n316 0.015
R10279 fout4.n305 fout4.n304 0.015
R10280 fout4.n75 fout4.n74 0.015
R10281 fout4.n83 fout4.n82 0.015
R10282 fout4.n94 fout4.n93 0.015
R10283 fout4.n92 fout4.n91 0.015
R10284 fout4.n365 fout4.n364 0.015
R10285 fout4.n9 fout4.n8 0.015
R10286 fout4.n395 fout4.n394 0.015
R10287 fout4.n400 fout4.n399 0.015
R10288 fout4.n523 fout4.n522 0.013
R10289 fout4.n508 fout4.n507 0.013
R10290 fout4.n332 fout4.n331 0.013
R10291 fout4.n238 fout4.n237 0.013
R10292 fout4.n274 fout4.n272 0.013
R10293 fout4.n44 fout4.n43 0.013
R10294 fout4.n46 fout4.n45 0.013
R10295 fout4.n307 fout4.n306 0.013
R10296 fout4.n34 fout4.n33 0.013
R10297 fout4.n36 fout4.n35 0.013
R10298 fout4.n349 fout4.n348 0.013
R10299 fout4.n382 fout4.n381 0.013
R10300 fout4.n386 fout4.n385 0.013
R10301 fout4.n539 fout4.n534 0.012
R10302 fout4.n539 fout4.n538 0.012
R10303 fout4.n493 fout4.n488 0.012
R10304 fout4.n493 fout4.n492 0.012
R10305 fout4.n431 fout4.n430 0.012
R10306 fout4.n434 fout4.n431 0.012
R10307 fout4.n200 fout4.n199 0.012
R10308 fout4.n199 fout4.n198 0.012
R10309 fout4.n158 fout4.n157 0.012
R10310 fout4.n157 fout4.n156 0.012
R10311 fout4.n66 fout4.n65 0.012
R10312 fout4.n65 fout4.n64 0.012
R10313 fout4.n360 fout4.n354 0.012
R10314 fout4.n360 fout4.n359 0.012
R10315 fout4.n520 fout4.n519 0.011
R10316 fout4.n513 fout4.n504 0.011
R10317 fout4.n474 fout4.n473 0.011
R10318 fout4.n467 fout4.n459 0.011
R10319 fout4.n422 fout4.n421 0.011
R10320 fout4.n450 fout4.n441 0.011
R10321 fout4.n297 fout4.n296 0.011
R10322 fout4.n122 fout4.n121 0.011
R10323 fout4.n203 fout4.n202 0.011
R10324 fout4.n196 fout4.n195 0.011
R10325 fout4.n161 fout4.n160 0.011
R10326 fout4.n154 fout4.n153 0.011
R10327 fout4.n69 fout4.n68 0.011
R10328 fout4.n62 fout4.n61 0.011
R10329 fout4.n377 fout4.n376 0.011
R10330 fout4.n5 fout4.n4 0.011
R10331 fout4.n426 fout4.n425 0.01
R10332 fout4.n440 fout4.n435 0.01
R10333 fout4.n375 fout4.n371 0.01
R10334 fout4.n405 fout4.n404 0.01
R10335 fout4.n404 fout4.n403 0.01
R10336 fout4.n323 fout4.n322 0.009
R10337 fout4.n233 fout4.n232 0.009
R10338 fout4.n237 fout4.n233 0.009
R10339 fout4.n260 fout4.n259 0.009
R10340 fout4.n110 fout4.n109 0.009
R10341 fout4.n216 fout4.n215 0.009
R10342 fout4.n180 fout4.n179 0.009
R10343 fout4.n408 fout4.n407 0.009
R10344 fout4.n230 fout4.n226 0.007
R10345 fout4.n263 fout4.n262 0.007
R10346 fout4.n258 fout4.n257 0.007
R10347 fout4.n255 fout4.n254 0.007
R10348 fout4.n111 fout4.n110 0.007
R10349 fout4.n23 fout4.n21 0.007
R10350 fout4.n310 fout4.n309 0.007
R10351 fout4.n182 fout4.n181 0.007
R10352 fout4.n177 fout4.n176 0.007
R10353 fout4.n175 fout4.n174 0.007
R10354 fout4.n18 fout4.n17 0.007
R10355 fout4.n519 fout4.n518 0.006
R10356 fout4.n504 fout4.n503 0.006
R10357 fout4.n513 fout4.n512 0.006
R10358 fout4.n473 fout4.n472 0.006
R10359 fout4.n459 fout4.n458 0.006
R10360 fout4.n467 fout4.n466 0.006
R10361 fout4.n425 fout4.n422 0.006
R10362 fout4.n441 fout4.n440 0.006
R10363 fout4.n450 fout4.n449 0.006
R10364 fout4.n348 fout4.n347 0.006
R10365 fout4.n204 fout4.n203 0.006
R10366 fout4.n202 fout4.n201 0.006
R10367 fout4.n197 fout4.n196 0.006
R10368 fout4.n195 fout4.n194 0.006
R10369 fout4.n162 fout4.n161 0.006
R10370 fout4.n160 fout4.n159 0.006
R10371 fout4.n155 fout4.n154 0.006
R10372 fout4.n153 fout4.n152 0.006
R10373 fout4.n70 fout4.n69 0.006
R10374 fout4.n68 fout4.n67 0.006
R10375 fout4.n63 fout4.n62 0.006
R10376 fout4.n61 fout4.n60 0.006
R10377 fout4.n377 fout4.n370 0.006
R10378 fout4.n376 fout4.n375 0.006
R10379 fout4.n4 fout4.n3 0.006
R10380 fout4.n342 fout4.n326 0.005
R10381 fout4.n338 fout4.n336 0.005
R10382 fout4.n302 fout4.n297 0.005
R10383 fout4.n295 fout4.n294 0.005
R10384 fout4.n267 fout4.n266 0.005
R10385 fout4.n253 fout4.n250 0.005
R10386 fout4.n121 fout4.n120 0.005
R10387 fout4.n107 fout4.n106 0.005
R10388 fout4.n207 fout4.n206 0.005
R10389 fout4.n128 fout4.n127 0.005
R10390 fout4.n89 fout4.n88 0.005
R10391 fout4.n409 fout4.n408 0.005
R10392 fout4.n407 fout4.n406 0.005
R10393 fout4.n541 fout4.n540 0.004
R10394 fout4.n495 fout4.n494 0.004
R10395 fout4.n421 fout4.n420 0.003
R10396 fout4.n514 fout4.n499 0.003
R10397 fout4.n468 fout4.n454 0.003
R10398 fout4.n452 fout4.n451 0.003
R10399 fout4.n361 fout4.n351 0.003
R10400 fout4.n379 fout4.n378 0.003
R10401 fout4.n213 fout4.n210 0.003
R10402 fout4.n81 fout4.n77 0.003
R10403 fout4.n137 fout4.n134 0.003
R10404 fout4.n126 fout4.n123 0.003
R10405 fout4.n108 fout4.n107 0.003
R10406 fout4.n50 fout4.n48 0.003
R10407 fout4.n55 fout4.n54 0.003
R10408 fout4.n27 fout4.n26 0.003
R10409 fout4.n166 fout4.n165 0.003
R10410 fout4.n33 fout4.n32 0.003
R10411 fout4.n528 fout4.n520 0.003
R10412 fout4.n482 fout4.n474 0.003
R10413 fout4.n13 fout4.n5 0.003
R10414 fout4.n412 fout4.n411 0.003
R10415 fout4.n413 fout4.n412 0.002
R10416 fout4.n494 fout4.n483 0.002
R10417 fout4.n540 fout4.n529 0.002
R10418 fout4.n451 fout4.n413 0.002
R10419 fout4.n483 fout4.n468 0.002
R10420 fout4.n529 fout4.n514 0.002
R10421 fout4.n378 fout4.n362 0.002
R10422 fout4.n362 fout4.n361 0.002
R10423 fout4.n331 fout4.n330 0.001
R10424 fout4.n222 fout4.n220 0.001
R10425 fout4.n225 fout4.n224 0.001
R10426 fout4.n231 fout4.n230 0.001
R10427 fout4.n288 fout4.n285 0.001
R10428 fout4.n283 fout4.n282 0.001
R10429 fout4.n277 fout4.n274 0.001
R10430 fout4.n271 fout4.n270 0.001
R10431 fout4.n262 fout4.n261 0.001
R10432 fout4.n256 fout4.n255 0.001
R10433 fout4.n250 fout4.n249 0.001
R10434 fout4.n120 fout4.n119 0.001
R10435 fout4.n316 fout4.n315 0.001
R10436 fout4.n312 fout4.n311 0.001
R10437 fout4.n173 fout4.n172 0.001
R10438 fout4.n74 fout4.n73 0.001
R10439 fout4.n96 fout4.n95 0.001
R10440 fout4.n498 fout4.n497 0.001
R10441 a_n20158_11542.n97 a_n20158_11542.t4 730.676
R10442 a_n20158_11542.n97 a_n20158_11542.t3 395.824
R10443 a_n20158_11542.n50 a_n20158_11542.n49 13.176
R10444 a_n20158_11542.n98 a_n20158_11542.t2 11.731
R10445 a_n20158_11542.n98 a_n20158_11542.t1 10.988
R10446 a_n20158_11542.n137 a_n20158_11542.n39 9.3
R10447 a_n20158_11542.n137 a_n20158_11542.n133 9.3
R10448 a_n20158_11542.n137 a_n20158_11542.n127 9.3
R10449 a_n20158_11542.n137 a_n20158_11542.n58 9.3
R10450 a_n20158_11542.n137 a_n20158_11542.n66 9.3
R10451 a_n20158_11542.n137 a_n20158_11542.n122 9.3
R10452 a_n20158_11542.n137 a_n20158_11542.n117 8.47
R10453 a_n20158_11542.n137 a_n20158_11542.n136 8.469
R10454 a_n20158_11542.n137 a_n20158_11542.n114 8.124
R10455 a_n20158_11542.n137 a_n20158_11542.n29 8.124
R10456 a_n20158_11542.n137 a_n20158_11542.n34 8.097
R10457 a_n20158_11542.n137 a_n20158_11542.n109 8.097
R10458 a_n20158_11542.n137 a_n20158_11542.n61 8.016
R10459 a_n20158_11542.n137 a_n20158_11542.n44 8.016
R10460 a_n20158_11542.n137 a_n20158_11542.n53 7.964
R10461 a_n20158_11542.n137 a_n20158_11542.n48 7.964
R10462 a_n20158_11542.n60 a_n20158_11542.n59 6.4
R10463 a_n20158_11542.n108 a_n20158_11542.n67 6.4
R10464 a_n20158_11542.n32 a_n20158_11542.n31 6.023
R10465 a_n20158_11542.n42 a_n20158_11542.n41 6.023
R10466 a_n20158_11542.n127 a_n20158_11542.n126 6.023
R10467 a_n20158_11542.n47 a_n20158_11542.n46 6.023
R10468 a_n20158_11542.n52 a_n20158_11542.n51 6.023
R10469 a_n20158_11542.n135 a_n20158_11542.n134 5.647
R10470 a_n20158_11542.n58 a_n20158_11542.n55 5.647
R10471 a_n20158_11542.n112 a_n20158_11542.n111 5.647
R10472 a_n20158_11542.n116 a_n20158_11542.n115 5.647
R10473 a_n20158_11542.n124 a_n20158_11542.n123 5.457
R10474 a_n20158_11542.n27 a_n20158_11542.n26 5.27
R10475 a_n20158_11542.n57 a_n20158_11542.n56 5.08
R10476 a_n20158_11542.n39 a_n20158_11542.n38 4.517
R10477 a_n20158_11542.n122 a_n20158_11542.n119 4.517
R10478 a_n20158_11542.n75 a_n20158_11542.n74 4.5
R10479 a_n20158_11542.n2 a_n20158_11542.n1 4.5
R10480 a_n20158_11542.n36 a_n20158_11542.n35 4.314
R10481 a_n20158_11542.n132 a_n20158_11542.n131 4.141
R10482 a_n20158_11542.n63 a_n20158_11542.n62 4.141
R10483 a_n20158_11542.n129 a_n20158_11542.n128 3.944
R10484 a_n20158_11542.n121 a_n20158_11542.n120 3.937
R10485 a_n20158_11542.n65 a_n20158_11542.n64 3.567
R10486 a_n20158_11542.n108 a_n20158_11542.n107 3.033
R10487 a_n20158_11542.t0 a_n20158_11542.n137 2.9
R10488 a_n20158_11542.n133 a_n20158_11542.n132 2.258
R10489 a_n20158_11542.n66 a_n20158_11542.n63 2.258
R10490 a_n20158_11542.n100 a_n20158_11542.n99 1.903
R10491 a_n20158_11542.n38 a_n20158_11542.n37 1.882
R10492 a_n20158_11542.n119 a_n20158_11542.n118 1.882
R10493 a_n20158_11542.n66 a_n20158_11542.n65 1.505
R10494 a_n20158_11542.n94 a_n20158_11542.n101 1.5
R10495 a_n20158_11542.n76 a_n20158_11542.n78 1.5
R10496 a_n20158_11542.n75 a_n20158_11542.n73 1.5
R10497 a_n20158_11542.n21 a_n20158_11542.n24 1.5
R10498 a_n20158_11542.n12 a_n20158_11542.n11 1.5
R10499 a_n20158_11542.n107 a_n20158_11542.n92 1.5
R10500 a_n20158_11542.n99 a_n20158_11542.n98 1.345
R10501 a_n20158_11542.n28 a_n20158_11542.n27 1.129
R10502 a_n20158_11542.n26 a_n20158_11542.n25 1.129
R10503 a_n20158_11542.n133 a_n20158_11542.n129 1.129
R10504 a_n20158_11542.n131 a_n20158_11542.n130 1.129
R10505 a_n20158_11542.n136 a_n20158_11542.n135 0.752
R10506 a_n20158_11542.n55 a_n20158_11542.n54 0.752
R10507 a_n20158_11542.n58 a_n20158_11542.n57 0.752
R10508 a_n20158_11542.n122 a_n20158_11542.n121 0.752
R10509 a_n20158_11542.n111 a_n20158_11542.n110 0.752
R10510 a_n20158_11542.n113 a_n20158_11542.n112 0.752
R10511 a_n20158_11542.n117 a_n20158_11542.n116 0.752
R10512 a_n20158_11542.n99 a_n20158_11542.n97 0.637
R10513 a_n20158_11542.n53 a_n20158_11542.n52 0.536
R10514 a_n20158_11542.n48 a_n20158_11542.n47 0.536
R10515 a_n20158_11542.n61 a_n20158_11542.n60 0.475
R10516 a_n20158_11542.n44 a_n20158_11542.n43 0.475
R10517 a_n20158_11542.n34 a_n20158_11542.n33 0.382
R10518 a_n20158_11542.n109 a_n20158_11542.n108 0.382
R10519 a_n20158_11542.n33 a_n20158_11542.n32 0.376
R10520 a_n20158_11542.n31 a_n20158_11542.n30 0.376
R10521 a_n20158_11542.n39 a_n20158_11542.n36 0.376
R10522 a_n20158_11542.n43 a_n20158_11542.n42 0.376
R10523 a_n20158_11542.n41 a_n20158_11542.n40 0.376
R10524 a_n20158_11542.n127 a_n20158_11542.n124 0.376
R10525 a_n20158_11542.n126 a_n20158_11542.n125 0.376
R10526 a_n20158_11542.n46 a_n20158_11542.n45 0.376
R10527 a_n20158_11542.n51 a_n20158_11542.n50 0.376
R10528 a_n20158_11542.n29 a_n20158_11542.n28 0.349
R10529 a_n20158_11542.n114 a_n20158_11542.n113 0.349
R10530 a_n20158_11542.n94 a_n20158_11542.n93 0.15
R10531 a_n20158_11542.n100 a_n20158_11542.n95 0.148
R10532 a_n20158_11542.n2 a_n20158_11542.n0 0.066
R10533 a_n20158_11542.n84 a_n20158_11542.n83 0.043
R10534 a_n20158_11542.n80 a_n20158_11542.n79 0.043
R10535 a_n20158_11542.n76 a_n20158_11542.n75 0.041
R10536 a_n20158_11542.n91 a_n20158_11542.n90 0.035
R10537 a_n20158_11542.n106 a_n20158_11542.n105 0.035
R10538 a_n20158_11542.n19 a_n20158_11542.n18 0.034
R10539 a_n20158_11542.n23 a_n20158_11542.n22 0.034
R10540 a_n20158_11542.n8 a_n20158_11542.n7 0.034
R10541 a_n20158_11542.n89 a_n20158_11542.n88 0.034
R10542 a_n20158_11542.n104 a_n20158_11542.n103 0.034
R10543 a_n20158_11542.n12 a_n20158_11542.n6 0.032
R10544 a_n20158_11542.n107 a_n20158_11542.n82 0.032
R10545 a_n20158_11542.n9 a_n20158_11542.n8 0.03
R10546 a_n20158_11542.n87 a_n20158_11542.n86 0.03
R10547 a_n20158_11542.n11 a_n20158_11542.n10 0.028
R10548 a_n20158_11542.n72 a_n20158_11542.n70 0.028
R10549 a_n20158_11542.n85 a_n20158_11542.n84 0.028
R10550 a_n20158_11542.n13 a_n20158_11542.n12 0.028
R10551 a_n20158_11542.n69 a_n20158_11542.n68 0.028
R10552 a_n20158_11542.n81 a_n20158_11542.n80 0.028
R10553 a_n20158_11542.n102 a_n20158_11542.n94 0.028
R10554 a_n20158_11542.n17 a_n20158_11542.n15 0.026
R10555 a_n20158_11542.n78 a_n20158_11542.n77 0.026
R10556 a_n20158_11542.n4 a_n20158_11542.n3 0.026
R10557 a_n20158_11542.n18 a_n20158_11542.n17 0.024
R10558 a_n20158_11542.n6 a_n20158_11542.n5 0.024
R10559 a_n20158_11542.n15 a_n20158_11542.n16 0.022
R10560 a_n20158_11542.n5 a_n20158_11542.n4 0.022
R10561 a_n20158_11542.n3 a_n20158_11542.n2 0.022
R10562 a_n20158_11542.n20 a_n20158_11542.n19 0.02
R10563 a_n20158_11542.n10 a_n20158_11542.n9 0.02
R10564 a_n20158_11542.n14 a_n20158_11542.n13 0.02
R10565 a_n20158_11542.n101 a_n20158_11542.n100 0.018
R10566 a_n20158_11542.n82 a_n20158_11542.n81 0.018
R10567 a_n20158_11542.n24 a_n20158_11542.n23 0.017
R10568 a_n20158_11542.n86 a_n20158_11542.n85 0.017
R10569 a_n20158_11542.n70 a_n20158_11542.n71 0.015
R10570 a_n20158_11542.n73 a_n20158_11542.n72 0.015
R10571 a_n20158_11542.n68 a_n20158_11542.n0 0.015
R10572 a_n20158_11542.n75 a_n20158_11542.n69 0.015
R10573 a_n20158_11542.n92 a_n20158_11542.n91 0.013
R10574 a_n20158_11542.n90 a_n20158_11542.n89 0.013
R10575 a_n20158_11542.n107 a_n20158_11542.n106 0.013
R10576 a_n20158_11542.n105 a_n20158_11542.n104 0.013
R10577 a_n20158_11542.n95 a_n20158_11542.n96 0.007
R10578 a_n20158_11542.n21 a_n20158_11542.n20 1.424
R10579 a_n20158_11542.n79 a_n20158_11542.n76 0.005
R10580 a_n20158_11542.n92 a_n20158_11542.n87 0.003
R10581 a_n20158_11542.n103 a_n20158_11542.n102 0.003
R10582 a_n20158_11542.n14 a_n20158_11542.n21 0.47
R10583 a_n21540_12270.n40 a_n21540_12270.t2 732.452
R10584 a_n21540_12270.n40 a_n21540_12270.t3 397.573
R10585 a_n21540_12270.n46 a_n21540_12270.n45 92.5
R10586 a_n21540_12270.n64 a_n21540_12270.n63 92.5
R10587 a_n21540_12270.n45 a_n21540_12270.t1 70.344
R10588 a_n21540_12270.n53 a_n21540_12270.n52 31.034
R10589 a_n21540_12270.n76 a_n21540_12270.n75 31.034
R10590 a_n21540_12270.n1 a_n21540_12270.n57 9.3
R10591 a_n21540_12270.n0 a_n21540_12270.n79 9.3
R10592 a_n21540_12270.n77 a_n21540_12270.n76 9.3
R10593 a_n21540_12270.n54 a_n21540_12270.n53 9.3
R10594 a_n21540_12270.n103 a_n21540_12270.n90 9.154
R10595 a_n21540_12270.n103 a_n21540_12270.n7 9.143
R10596 a_n21540_12270.n103 a_n21540_12270.n6 9.143
R10597 a_n21540_12270.n103 a_n21540_12270.n22 9.132
R10598 a_n21540_12270.n103 a_n21540_12270.n96 9.132
R10599 a_n21540_12270.n103 a_n21540_12270.n100 8.886
R10600 a_n21540_12270.n103 a_n21540_12270.n26 8.885
R10601 a_n21540_12270.n103 a_n21540_12270.n11 8.875
R10602 a_n21540_12270.n103 a_n21540_12270.n32 8.875
R10603 a_n21540_12270.n103 a_n21540_12270.n102 8.864
R10604 a_n21540_12270.n103 a_n21540_12270.n28 8.864
R10605 a_n21540_12270.n47 a_n21540_12270.n46 8.282
R10606 a_n21540_12270.n65 a_n21540_12270.n64 8.282
R10607 a_n21540_12270.t0 a_n21540_12270.n103 7.141
R10608 a_n21540_12270.n54 a_n21540_12270.n50 5.647
R10609 a_n21540_12270.n77 a_n21540_12270.n73 5.647
R10610 a_n21540_12270.n84 a_n21540_12270.n83 4.723
R10611 a_n21540_12270.n2 a_n21540_12270.n62 4.65
R10612 a_n21540_12270.n90 a_n21540_12270.n85 4.65
R10613 a_n21540_12270.n83 a_n21540_12270.n3 4.566
R10614 a_n21540_12270.n90 a_n21540_12270.n39 4.517
R10615 a_n21540_12270.n66 a_n21540_12270.n65 4.5
R10616 a_n21540_12270.n67 a_n21540_12270.n69 4.5
R10617 a_n21540_12270.n43 a_n21540_12270.n47 4.5
R10618 a_n21540_12270.n70 a_n21540_12270.n78 4.5
R10619 a_n21540_12270.n2 a_n21540_12270.n61 4.5
R10620 a_n21540_12270.n4 a_n21540_12270.n56 4.5
R10621 a_n21540_12270.n0 a_n21540_12270.n82 4.5
R10622 a_n21540_12270.n1 a_n21540_12270.n60 4.5
R10623 a_n21540_12270.n98 a_n21540_12270.n97 4.141
R10624 a_n21540_12270.n90 a_n21540_12270.n38 4.141
R10625 a_n21540_12270.n24 a_n21540_12270.n23 4.141
R10626 a_n21540_12270.n52 a_n21540_12270.n51 4.137
R10627 a_n21540_12270.n75 a_n21540_12270.n74 4.137
R10628 a_n21540_12270.n60 a_n21540_12270.n58 3.764
R10629 a_n21540_12270.n78 a_n21540_12270.n71 3.764
R10630 a_n21540_12270.n92 a_n21540_12270.n91 3.764
R10631 a_n21540_12270.n7 a_n21540_12270.n34 3.764
R10632 a_n21540_12270.n96 a_n21540_12270.n95 3.736
R10633 a_n21540_12270.n56 a_n21540_12270.n55 3.388
R10634 a_n21540_12270.n82 a_n21540_12270.n81 3.388
R10635 a_n21540_12270.n9 a_n21540_12270.n8 3.388
R10636 a_n21540_12270.n6 a_n21540_12270.n13 3.388
R10637 a_n21540_12270.n18 a_n21540_12270.n17 3.388
R10638 a_n21540_12270.n30 a_n21540_12270.n29 3.388
R10639 a_n21540_12270.n22 a_n21540_12270.n21 3.36
R10640 a_n21540_12270.n56 a_n21540_12270.n54 3.011
R10641 a_n21540_12270.n47 a_n21540_12270.n44 3.011
R10642 a_n21540_12270.n82 a_n21540_12270.n80 3.011
R10643 a_n21540_12270.n10 a_n21540_12270.n9 3.011
R10644 a_n21540_12270.n13 a_n21540_12270.n12 3.011
R10645 a_n21540_12270.n16 a_n21540_12270.n15 3.011
R10646 a_n21540_12270.n21 a_n21540_12270.n20 3.011
R10647 a_n21540_12270.n19 a_n21540_12270.n18 3.011
R10648 a_n21540_12270.n31 a_n21540_12270.n30 3.011
R10649 a_n21540_12270.n60 a_n21540_12270.n59 2.635
R10650 a_n21540_12270.n69 a_n21540_12270.n68 2.635
R10651 a_n21540_12270.n78 a_n21540_12270.n77 2.635
R10652 a_n21540_12270.n93 a_n21540_12270.n92 2.635
R10653 a_n21540_12270.n95 a_n21540_12270.n94 2.635
R10654 a_n21540_12270.n37 a_n21540_12270.n36 2.635
R10655 a_n21540_12270.n34 a_n21540_12270.n33 2.635
R10656 a_n21540_12270.n83 a_n21540_12270.n40 2.35
R10657 a_n21540_12270.n99 a_n21540_12270.n98 2.258
R10658 a_n21540_12270.n25 a_n21540_12270.n24 2.258
R10659 a_n21540_12270.n5 a_n21540_12270.n89 1.619
R10660 a_n21540_12270.n86 a_n21540_12270.n87 1.588
R10661 a_n21540_12270.n5 a_n21540_12270.n104 1.88
R10662 a_n21540_12270.n3 a_n21540_12270.n0 2.375
R10663 a_n21540_12270.n7 a_n21540_12270.n37 2.257
R10664 a_n21540_12270.n6 a_n21540_12270.n16 2.257
R10665 a_n21540_12270.n36 a_n21540_12270.n35 1.505
R10666 a_n21540_12270.n42 a_n21540_12270.n1 1.5
R10667 a_n21540_12270.n15 a_n21540_12270.n14 1.129
R10668 a_n21540_12270.n50 a_n21540_12270.n49 0.752
R10669 a_n21540_12270.n73 a_n21540_12270.n72 0.752
R10670 a_n21540_12270.n42 a_n21540_12270.n41 0.24
R10671 a_n21540_12270.n102 a_n21540_12270.n101 0.155
R10672 a_n21540_12270.n28 a_n21540_12270.n27 0.155
R10673 a_n21540_12270.n11 a_n21540_12270.n10 0.144
R10674 a_n21540_12270.n32 a_n21540_12270.n31 0.144
R10675 a_n21540_12270.n100 a_n21540_12270.n99 0.133
R10676 a_n21540_12270.n26 a_n21540_12270.n25 0.132
R10677 a_n21540_12270.n67 a_n21540_12270.n66 0.082
R10678 a_n21540_12270.n43 a_n21540_12270.n48 0.071
R10679 a_n21540_12270.n70 a_n21540_12270.n67 0.042
R10680 a_n21540_12270.n87 a_n21540_12270.n88 0.024
R10681 a_n21540_12270.n22 a_n21540_12270.n19 0.024
R10682 a_n21540_12270.n96 a_n21540_12270.n93 0.024
R10683 a_n21540_12270.n85 a_n21540_12270.n86 0.147
R10684 a_n21540_12270.n86 a_n21540_12270.n5 0.124
R10685 a_n21540_12270.n85 a_n21540_12270.n84 2.702
R10686 a_n21540_12270.n3 a_n21540_12270.n42 0.955
R10687 a_n21540_12270.n0 a_n21540_12270.n70 0.127
R10688 a_n21540_12270.n1 a_n21540_12270.n4 0.11
R10689 a_n21540_12270.n4 a_n21540_12270.n43 0.058
R10690 a_n21540_12270.n66 a_n21540_12270.n2 0.042
R10691 a_n14372_11547.n97 a_n14372_11547.t4 730.681
R10692 a_n14372_11547.n97 a_n14372_11547.t3 395.834
R10693 a_n14372_11547.n50 a_n14372_11547.n49 13.176
R10694 a_n14372_11547.n98 a_n14372_11547.t1 11.724
R10695 a_n14372_11547.n98 a_n14372_11547.t0 10.994
R10696 a_n14372_11547.n137 a_n14372_11547.n39 9.3
R10697 a_n14372_11547.n137 a_n14372_11547.n133 9.3
R10698 a_n14372_11547.n137 a_n14372_11547.n127 9.3
R10699 a_n14372_11547.n137 a_n14372_11547.n58 9.3
R10700 a_n14372_11547.n137 a_n14372_11547.n66 9.3
R10701 a_n14372_11547.n137 a_n14372_11547.n122 9.3
R10702 a_n14372_11547.n137 a_n14372_11547.n117 8.47
R10703 a_n14372_11547.n137 a_n14372_11547.n136 8.469
R10704 a_n14372_11547.n137 a_n14372_11547.n114 8.124
R10705 a_n14372_11547.n137 a_n14372_11547.n29 8.124
R10706 a_n14372_11547.n137 a_n14372_11547.n34 8.097
R10707 a_n14372_11547.n137 a_n14372_11547.n109 8.097
R10708 a_n14372_11547.n137 a_n14372_11547.n61 8.016
R10709 a_n14372_11547.n137 a_n14372_11547.n44 8.016
R10710 a_n14372_11547.n137 a_n14372_11547.n53 7.964
R10711 a_n14372_11547.n137 a_n14372_11547.n48 7.964
R10712 a_n14372_11547.n60 a_n14372_11547.n59 6.4
R10713 a_n14372_11547.n108 a_n14372_11547.n67 6.4
R10714 a_n14372_11547.n32 a_n14372_11547.n31 6.023
R10715 a_n14372_11547.n42 a_n14372_11547.n41 6.023
R10716 a_n14372_11547.n127 a_n14372_11547.n126 6.023
R10717 a_n14372_11547.n47 a_n14372_11547.n46 6.023
R10718 a_n14372_11547.n52 a_n14372_11547.n51 6.023
R10719 a_n14372_11547.n135 a_n14372_11547.n134 5.647
R10720 a_n14372_11547.n58 a_n14372_11547.n55 5.647
R10721 a_n14372_11547.n112 a_n14372_11547.n111 5.647
R10722 a_n14372_11547.n116 a_n14372_11547.n115 5.647
R10723 a_n14372_11547.n124 a_n14372_11547.n123 5.457
R10724 a_n14372_11547.n27 a_n14372_11547.n26 5.27
R10725 a_n14372_11547.n57 a_n14372_11547.n56 5.08
R10726 a_n14372_11547.n39 a_n14372_11547.n38 4.517
R10727 a_n14372_11547.n122 a_n14372_11547.n119 4.517
R10728 a_n14372_11547.n75 a_n14372_11547.n74 4.5
R10729 a_n14372_11547.n2 a_n14372_11547.n1 4.5
R10730 a_n14372_11547.n36 a_n14372_11547.n35 4.314
R10731 a_n14372_11547.n132 a_n14372_11547.n131 4.141
R10732 a_n14372_11547.n63 a_n14372_11547.n62 4.141
R10733 a_n14372_11547.n129 a_n14372_11547.n128 3.944
R10734 a_n14372_11547.n121 a_n14372_11547.n120 3.937
R10735 a_n14372_11547.n65 a_n14372_11547.n64 3.567
R10736 a_n14372_11547.n108 a_n14372_11547.n107 3.033
R10737 a_n14372_11547.t2 a_n14372_11547.n137 2.9
R10738 a_n14372_11547.n133 a_n14372_11547.n132 2.258
R10739 a_n14372_11547.n66 a_n14372_11547.n63 2.258
R10740 a_n14372_11547.n100 a_n14372_11547.n99 1.903
R10741 a_n14372_11547.n38 a_n14372_11547.n37 1.882
R10742 a_n14372_11547.n119 a_n14372_11547.n118 1.882
R10743 a_n14372_11547.n66 a_n14372_11547.n65 1.505
R10744 a_n14372_11547.n94 a_n14372_11547.n101 1.5
R10745 a_n14372_11547.n76 a_n14372_11547.n78 1.5
R10746 a_n14372_11547.n75 a_n14372_11547.n73 1.5
R10747 a_n14372_11547.n21 a_n14372_11547.n24 1.5
R10748 a_n14372_11547.n12 a_n14372_11547.n11 1.5
R10749 a_n14372_11547.n107 a_n14372_11547.n92 1.5
R10750 a_n14372_11547.n99 a_n14372_11547.n98 1.223
R10751 a_n14372_11547.n28 a_n14372_11547.n27 1.129
R10752 a_n14372_11547.n26 a_n14372_11547.n25 1.129
R10753 a_n14372_11547.n133 a_n14372_11547.n129 1.129
R10754 a_n14372_11547.n131 a_n14372_11547.n130 1.129
R10755 a_n14372_11547.n136 a_n14372_11547.n135 0.752
R10756 a_n14372_11547.n55 a_n14372_11547.n54 0.752
R10757 a_n14372_11547.n58 a_n14372_11547.n57 0.752
R10758 a_n14372_11547.n122 a_n14372_11547.n121 0.752
R10759 a_n14372_11547.n111 a_n14372_11547.n110 0.752
R10760 a_n14372_11547.n113 a_n14372_11547.n112 0.752
R10761 a_n14372_11547.n117 a_n14372_11547.n116 0.752
R10762 a_n14372_11547.n99 a_n14372_11547.n97 0.637
R10763 a_n14372_11547.n53 a_n14372_11547.n52 0.536
R10764 a_n14372_11547.n48 a_n14372_11547.n47 0.536
R10765 a_n14372_11547.n61 a_n14372_11547.n60 0.475
R10766 a_n14372_11547.n44 a_n14372_11547.n43 0.475
R10767 a_n14372_11547.n34 a_n14372_11547.n33 0.382
R10768 a_n14372_11547.n109 a_n14372_11547.n108 0.382
R10769 a_n14372_11547.n33 a_n14372_11547.n32 0.376
R10770 a_n14372_11547.n31 a_n14372_11547.n30 0.376
R10771 a_n14372_11547.n39 a_n14372_11547.n36 0.376
R10772 a_n14372_11547.n43 a_n14372_11547.n42 0.376
R10773 a_n14372_11547.n41 a_n14372_11547.n40 0.376
R10774 a_n14372_11547.n127 a_n14372_11547.n124 0.376
R10775 a_n14372_11547.n126 a_n14372_11547.n125 0.376
R10776 a_n14372_11547.n46 a_n14372_11547.n45 0.376
R10777 a_n14372_11547.n51 a_n14372_11547.n50 0.376
R10778 a_n14372_11547.n29 a_n14372_11547.n28 0.349
R10779 a_n14372_11547.n114 a_n14372_11547.n113 0.349
R10780 a_n14372_11547.n94 a_n14372_11547.n93 0.15
R10781 a_n14372_11547.n100 a_n14372_11547.n95 0.148
R10782 a_n14372_11547.n2 a_n14372_11547.n0 0.066
R10783 a_n14372_11547.n84 a_n14372_11547.n83 0.043
R10784 a_n14372_11547.n80 a_n14372_11547.n79 0.043
R10785 a_n14372_11547.n76 a_n14372_11547.n75 0.041
R10786 a_n14372_11547.n91 a_n14372_11547.n90 0.035
R10787 a_n14372_11547.n106 a_n14372_11547.n105 0.035
R10788 a_n14372_11547.n19 a_n14372_11547.n18 0.034
R10789 a_n14372_11547.n23 a_n14372_11547.n22 0.034
R10790 a_n14372_11547.n8 a_n14372_11547.n7 0.034
R10791 a_n14372_11547.n89 a_n14372_11547.n88 0.034
R10792 a_n14372_11547.n104 a_n14372_11547.n103 0.034
R10793 a_n14372_11547.n12 a_n14372_11547.n6 0.032
R10794 a_n14372_11547.n107 a_n14372_11547.n82 0.032
R10795 a_n14372_11547.n9 a_n14372_11547.n8 0.03
R10796 a_n14372_11547.n87 a_n14372_11547.n86 0.03
R10797 a_n14372_11547.n11 a_n14372_11547.n10 0.028
R10798 a_n14372_11547.n72 a_n14372_11547.n70 0.028
R10799 a_n14372_11547.n85 a_n14372_11547.n84 0.028
R10800 a_n14372_11547.n13 a_n14372_11547.n12 0.028
R10801 a_n14372_11547.n69 a_n14372_11547.n68 0.028
R10802 a_n14372_11547.n81 a_n14372_11547.n80 0.028
R10803 a_n14372_11547.n102 a_n14372_11547.n94 0.028
R10804 a_n14372_11547.n17 a_n14372_11547.n15 0.026
R10805 a_n14372_11547.n78 a_n14372_11547.n77 0.026
R10806 a_n14372_11547.n4 a_n14372_11547.n3 0.026
R10807 a_n14372_11547.n18 a_n14372_11547.n17 0.024
R10808 a_n14372_11547.n6 a_n14372_11547.n5 0.024
R10809 a_n14372_11547.n15 a_n14372_11547.n16 0.022
R10810 a_n14372_11547.n5 a_n14372_11547.n4 0.022
R10811 a_n14372_11547.n3 a_n14372_11547.n2 0.022
R10812 a_n14372_11547.n20 a_n14372_11547.n19 0.02
R10813 a_n14372_11547.n10 a_n14372_11547.n9 0.02
R10814 a_n14372_11547.n14 a_n14372_11547.n13 0.02
R10815 a_n14372_11547.n101 a_n14372_11547.n100 0.018
R10816 a_n14372_11547.n82 a_n14372_11547.n81 0.018
R10817 a_n14372_11547.n24 a_n14372_11547.n23 0.017
R10818 a_n14372_11547.n86 a_n14372_11547.n85 0.017
R10819 a_n14372_11547.n70 a_n14372_11547.n71 0.015
R10820 a_n14372_11547.n73 a_n14372_11547.n72 0.015
R10821 a_n14372_11547.n68 a_n14372_11547.n0 0.015
R10822 a_n14372_11547.n75 a_n14372_11547.n69 0.015
R10823 a_n14372_11547.n92 a_n14372_11547.n91 0.013
R10824 a_n14372_11547.n90 a_n14372_11547.n89 0.013
R10825 a_n14372_11547.n107 a_n14372_11547.n106 0.013
R10826 a_n14372_11547.n105 a_n14372_11547.n104 0.013
R10827 a_n14372_11547.n95 a_n14372_11547.n96 0.007
R10828 a_n14372_11547.n21 a_n14372_11547.n20 1.424
R10829 a_n14372_11547.n79 a_n14372_11547.n76 0.005
R10830 a_n14372_11547.n92 a_n14372_11547.n87 0.003
R10831 a_n14372_11547.n103 a_n14372_11547.n102 0.003
R10832 a_n14372_11547.n14 a_n14372_11547.n21 0.47
R10833 a_n15755_12275.n40 a_n15755_12275.t3 732.457
R10834 a_n15755_12275.n40 a_n15755_12275.t2 397.579
R10835 a_n15755_12275.n46 a_n15755_12275.n45 92.5
R10836 a_n15755_12275.n64 a_n15755_12275.n63 92.5
R10837 a_n15755_12275.n45 a_n15755_12275.t1 70.344
R10838 a_n15755_12275.n53 a_n15755_12275.n52 31.034
R10839 a_n15755_12275.n76 a_n15755_12275.n75 31.034
R10840 a_n15755_12275.n1 a_n15755_12275.n57 9.3
R10841 a_n15755_12275.n0 a_n15755_12275.n79 9.3
R10842 a_n15755_12275.n77 a_n15755_12275.n76 9.3
R10843 a_n15755_12275.n54 a_n15755_12275.n53 9.3
R10844 a_n15755_12275.n103 a_n15755_12275.n90 9.154
R10845 a_n15755_12275.n103 a_n15755_12275.n7 9.143
R10846 a_n15755_12275.n103 a_n15755_12275.n6 9.143
R10847 a_n15755_12275.n103 a_n15755_12275.n22 9.132
R10848 a_n15755_12275.n103 a_n15755_12275.n96 9.132
R10849 a_n15755_12275.n103 a_n15755_12275.n100 8.886
R10850 a_n15755_12275.n103 a_n15755_12275.n26 8.885
R10851 a_n15755_12275.n103 a_n15755_12275.n11 8.875
R10852 a_n15755_12275.n103 a_n15755_12275.n32 8.875
R10853 a_n15755_12275.n103 a_n15755_12275.n102 8.864
R10854 a_n15755_12275.n103 a_n15755_12275.n28 8.864
R10855 a_n15755_12275.n47 a_n15755_12275.n46 8.282
R10856 a_n15755_12275.n65 a_n15755_12275.n64 8.282
R10857 a_n15755_12275.t0 a_n15755_12275.n103 7.141
R10858 a_n15755_12275.n54 a_n15755_12275.n50 5.647
R10859 a_n15755_12275.n77 a_n15755_12275.n73 5.647
R10860 a_n15755_12275.n84 a_n15755_12275.n83 4.722
R10861 a_n15755_12275.n2 a_n15755_12275.n62 4.65
R10862 a_n15755_12275.n90 a_n15755_12275.n85 4.65
R10863 a_n15755_12275.n83 a_n15755_12275.n3 4.565
R10864 a_n15755_12275.n90 a_n15755_12275.n39 4.517
R10865 a_n15755_12275.n66 a_n15755_12275.n65 4.5
R10866 a_n15755_12275.n67 a_n15755_12275.n69 4.5
R10867 a_n15755_12275.n43 a_n15755_12275.n47 4.5
R10868 a_n15755_12275.n70 a_n15755_12275.n78 4.5
R10869 a_n15755_12275.n2 a_n15755_12275.n61 4.5
R10870 a_n15755_12275.n4 a_n15755_12275.n56 4.5
R10871 a_n15755_12275.n0 a_n15755_12275.n82 4.5
R10872 a_n15755_12275.n1 a_n15755_12275.n60 4.5
R10873 a_n15755_12275.n98 a_n15755_12275.n97 4.141
R10874 a_n15755_12275.n90 a_n15755_12275.n38 4.141
R10875 a_n15755_12275.n24 a_n15755_12275.n23 4.141
R10876 a_n15755_12275.n52 a_n15755_12275.n51 4.137
R10877 a_n15755_12275.n75 a_n15755_12275.n74 4.137
R10878 a_n15755_12275.n60 a_n15755_12275.n58 3.764
R10879 a_n15755_12275.n78 a_n15755_12275.n71 3.764
R10880 a_n15755_12275.n92 a_n15755_12275.n91 3.764
R10881 a_n15755_12275.n7 a_n15755_12275.n34 3.764
R10882 a_n15755_12275.n96 a_n15755_12275.n95 3.736
R10883 a_n15755_12275.n56 a_n15755_12275.n55 3.388
R10884 a_n15755_12275.n82 a_n15755_12275.n81 3.388
R10885 a_n15755_12275.n9 a_n15755_12275.n8 3.388
R10886 a_n15755_12275.n6 a_n15755_12275.n13 3.388
R10887 a_n15755_12275.n18 a_n15755_12275.n17 3.388
R10888 a_n15755_12275.n30 a_n15755_12275.n29 3.388
R10889 a_n15755_12275.n22 a_n15755_12275.n21 3.36
R10890 a_n15755_12275.n56 a_n15755_12275.n54 3.011
R10891 a_n15755_12275.n47 a_n15755_12275.n44 3.011
R10892 a_n15755_12275.n82 a_n15755_12275.n80 3.011
R10893 a_n15755_12275.n10 a_n15755_12275.n9 3.011
R10894 a_n15755_12275.n13 a_n15755_12275.n12 3.011
R10895 a_n15755_12275.n16 a_n15755_12275.n15 3.011
R10896 a_n15755_12275.n21 a_n15755_12275.n20 3.011
R10897 a_n15755_12275.n19 a_n15755_12275.n18 3.011
R10898 a_n15755_12275.n31 a_n15755_12275.n30 3.011
R10899 a_n15755_12275.n60 a_n15755_12275.n59 2.635
R10900 a_n15755_12275.n69 a_n15755_12275.n68 2.635
R10901 a_n15755_12275.n78 a_n15755_12275.n77 2.635
R10902 a_n15755_12275.n93 a_n15755_12275.n92 2.635
R10903 a_n15755_12275.n95 a_n15755_12275.n94 2.635
R10904 a_n15755_12275.n37 a_n15755_12275.n36 2.635
R10905 a_n15755_12275.n34 a_n15755_12275.n33 2.635
R10906 a_n15755_12275.n83 a_n15755_12275.n40 2.349
R10907 a_n15755_12275.n99 a_n15755_12275.n98 2.258
R10908 a_n15755_12275.n25 a_n15755_12275.n24 2.258
R10909 a_n15755_12275.n5 a_n15755_12275.n89 1.619
R10910 a_n15755_12275.n86 a_n15755_12275.n87 1.588
R10911 a_n15755_12275.n5 a_n15755_12275.n104 1.88
R10912 a_n15755_12275.n3 a_n15755_12275.n0 2.375
R10913 a_n15755_12275.n7 a_n15755_12275.n37 2.257
R10914 a_n15755_12275.n6 a_n15755_12275.n16 2.257
R10915 a_n15755_12275.n36 a_n15755_12275.n35 1.505
R10916 a_n15755_12275.n42 a_n15755_12275.n1 1.5
R10917 a_n15755_12275.n15 a_n15755_12275.n14 1.129
R10918 a_n15755_12275.n50 a_n15755_12275.n49 0.752
R10919 a_n15755_12275.n73 a_n15755_12275.n72 0.752
R10920 a_n15755_12275.n42 a_n15755_12275.n41 0.24
R10921 a_n15755_12275.n102 a_n15755_12275.n101 0.155
R10922 a_n15755_12275.n28 a_n15755_12275.n27 0.155
R10923 a_n15755_12275.n11 a_n15755_12275.n10 0.144
R10924 a_n15755_12275.n32 a_n15755_12275.n31 0.144
R10925 a_n15755_12275.n100 a_n15755_12275.n99 0.133
R10926 a_n15755_12275.n26 a_n15755_12275.n25 0.132
R10927 a_n15755_12275.n67 a_n15755_12275.n66 0.082
R10928 a_n15755_12275.n43 a_n15755_12275.n48 0.071
R10929 a_n15755_12275.n70 a_n15755_12275.n67 0.042
R10930 a_n15755_12275.n87 a_n15755_12275.n88 0.024
R10931 a_n15755_12275.n22 a_n15755_12275.n19 0.024
R10932 a_n15755_12275.n96 a_n15755_12275.n93 0.024
R10933 a_n15755_12275.n85 a_n15755_12275.n86 0.147
R10934 a_n15755_12275.n86 a_n15755_12275.n5 0.124
R10935 a_n15755_12275.n85 a_n15755_12275.n84 2.702
R10936 a_n15755_12275.n3 a_n15755_12275.n42 0.955
R10937 a_n15755_12275.n0 a_n15755_12275.n70 0.127
R10938 a_n15755_12275.n1 a_n15755_12275.n4 0.11
R10939 a_n15755_12275.n4 a_n15755_12275.n43 0.058
R10940 a_n15755_12275.n66 a_n15755_12275.n2 0.042
R10941 a_n17562_12353.n60 a_n17562_12353.t3 735.929
R10942 a_n17562_12353.n54 a_n17562_12353.t5 396.755
R10943 a_n17562_12353.n66 a_n17562_12353.t2 396.755
R10944 a_n17562_12353.n80 a_n17562_12353.n79 92.5
R10945 a_n17562_12353.n98 a_n17562_12353.n97 92.5
R10946 a_n17562_12353.n79 a_n17562_12353.t1 70.344
R10947 a_n17562_12353.n87 a_n17562_12353.n86 31.034
R10948 a_n17562_12353.n110 a_n17562_12353.n109 31.034
R10949 a_n17562_12353.n1 a_n17562_12353.n91 9.3
R10950 a_n17562_12353.n0 a_n17562_12353.n113 9.3
R10951 a_n17562_12353.n111 a_n17562_12353.n110 9.3
R10952 a_n17562_12353.n88 a_n17562_12353.n87 9.3
R10953 a_n17562_12353.n137 a_n17562_12353.n124 9.154
R10954 a_n17562_12353.n137 a_n17562_12353.n7 9.143
R10955 a_n17562_12353.n137 a_n17562_12353.n6 9.143
R10956 a_n17562_12353.n137 a_n17562_12353.n30 9.132
R10957 a_n17562_12353.n137 a_n17562_12353.n130 9.132
R10958 a_n17562_12353.n137 a_n17562_12353.n134 8.886
R10959 a_n17562_12353.n137 a_n17562_12353.n34 8.885
R10960 a_n17562_12353.n137 a_n17562_12353.n19 8.875
R10961 a_n17562_12353.n137 a_n17562_12353.n40 8.875
R10962 a_n17562_12353.n137 a_n17562_12353.n136 8.864
R10963 a_n17562_12353.n137 a_n17562_12353.n36 8.864
R10964 a_n17562_12353.n81 a_n17562_12353.n80 8.282
R10965 a_n17562_12353.n99 a_n17562_12353.n98 8.282
R10966 a_n17562_12353.t0 a_n17562_12353.n137 7.141
R10967 a_n17562_12353.n118 a_n17562_12353.n117 6.622
R10968 a_n17562_12353.n88 a_n17562_12353.n84 5.647
R10969 a_n17562_12353.n111 a_n17562_12353.n107 5.647
R10970 a_n17562_12353.n2 a_n17562_12353.n96 4.65
R10971 a_n17562_12353.n124 a_n17562_12353.n119 4.65
R10972 a_n17562_12353.n124 a_n17562_12353.n47 4.517
R10973 a_n17562_12353.n100 a_n17562_12353.n99 4.5
R10974 a_n17562_12353.n101 a_n17562_12353.n103 4.5
R10975 a_n17562_12353.n77 a_n17562_12353.n81 4.5
R10976 a_n17562_12353.n104 a_n17562_12353.n112 4.5
R10977 a_n17562_12353.n2 a_n17562_12353.n95 4.5
R10978 a_n17562_12353.n4 a_n17562_12353.n90 4.5
R10979 a_n17562_12353.n0 a_n17562_12353.n116 4.5
R10980 a_n17562_12353.n1 a_n17562_12353.n94 4.5
R10981 a_n17562_12353.n132 a_n17562_12353.n131 4.141
R10982 a_n17562_12353.n124 a_n17562_12353.n46 4.141
R10983 a_n17562_12353.n32 a_n17562_12353.n31 4.141
R10984 a_n17562_12353.n86 a_n17562_12353.n85 4.137
R10985 a_n17562_12353.n109 a_n17562_12353.n108 4.137
R10986 a_n17562_12353.n94 a_n17562_12353.n92 3.764
R10987 a_n17562_12353.n112 a_n17562_12353.n105 3.764
R10988 a_n17562_12353.n126 a_n17562_12353.n125 3.764
R10989 a_n17562_12353.n7 a_n17562_12353.n42 3.764
R10990 a_n17562_12353.n13 a_n17562_12353.n55 3.758
R10991 a_n17562_12353.n130 a_n17562_12353.n129 3.736
R10992 a_n17562_12353.n12 a_n17562_12353.n66 3.633
R10993 a_n17562_12353.n90 a_n17562_12353.n89 3.388
R10994 a_n17562_12353.n116 a_n17562_12353.n115 3.388
R10995 a_n17562_12353.n17 a_n17562_12353.n16 3.388
R10996 a_n17562_12353.n6 a_n17562_12353.n21 3.388
R10997 a_n17562_12353.n26 a_n17562_12353.n25 3.388
R10998 a_n17562_12353.n38 a_n17562_12353.n37 3.388
R10999 a_n17562_12353.n30 a_n17562_12353.n29 3.36
R11000 a_n17562_12353.n90 a_n17562_12353.n88 3.011
R11001 a_n17562_12353.n81 a_n17562_12353.n78 3.011
R11002 a_n17562_12353.n116 a_n17562_12353.n114 3.011
R11003 a_n17562_12353.n18 a_n17562_12353.n17 3.011
R11004 a_n17562_12353.n21 a_n17562_12353.n20 3.011
R11005 a_n17562_12353.n24 a_n17562_12353.n23 3.011
R11006 a_n17562_12353.n29 a_n17562_12353.n28 3.011
R11007 a_n17562_12353.n27 a_n17562_12353.n26 3.011
R11008 a_n17562_12353.n39 a_n17562_12353.n38 3.011
R11009 a_n17562_12353.n94 a_n17562_12353.n93 2.635
R11010 a_n17562_12353.n103 a_n17562_12353.n102 2.635
R11011 a_n17562_12353.n112 a_n17562_12353.n111 2.635
R11012 a_n17562_12353.n127 a_n17562_12353.n126 2.635
R11013 a_n17562_12353.n129 a_n17562_12353.n128 2.635
R11014 a_n17562_12353.n45 a_n17562_12353.n44 2.635
R11015 a_n17562_12353.n42 a_n17562_12353.n41 2.635
R11016 a_n17562_12353.n117 a_n17562_12353.n3 2.631
R11017 a_n17562_12353.n74 a_n17562_12353.n71 2.621
R11018 a_n17562_12353.n15 a_n17562_12353.n54 3.627
R11019 a_n17562_12353.n133 a_n17562_12353.n132 2.258
R11020 a_n17562_12353.n33 a_n17562_12353.n32 2.258
R11021 a_n17562_12353.n5 a_n17562_12353.n123 1.619
R11022 a_n17562_12353.n120 a_n17562_12353.n121 1.588
R11023 a_n17562_12353.n5 a_n17562_12353.n138 1.88
R11024 a_n17562_12353.n3 a_n17562_12353.n0 2.375
R11025 a_n17562_12353.n44 a_n17562_12353.n43 1.505
R11026 a_n17562_12353.n76 a_n17562_12353.n1 1.5
R11027 a_n17562_12353.n7 a_n17562_12353.n45 2.257
R11028 a_n17562_12353.n6 a_n17562_12353.n24 2.257
R11029 a_n17562_12353.n9 a_n17562_12353.n8 1.149
R11030 a_n17562_12353.n59 a_n17562_12353.n57 1.149
R11031 a_n17562_12353.n11 a_n17562_12353.n10 1.149
R11032 a_n17562_12353.n12 a_n17562_12353.n63 1.148
R11033 a_n17562_12353.n15 a_n17562_12353.n9 1.138
R11034 a_n17562_12353.n14 a_n17562_12353.t4 737.068
R11035 a_n17562_12353.n63 a_n17562_12353.n61 1.137
R11036 a_n17562_12353.n11 a_n17562_12353.n67 1.137
R11037 a_n17562_12353.n14 a_n17562_12353.n74 1.136
R11038 a_n17562_12353.n13 a_n17562_12353.n59 1.136
R11039 a_n17562_12353.n23 a_n17562_12353.n22 1.129
R11040 a_n17562_12353.n84 a_n17562_12353.n83 0.752
R11041 a_n17562_12353.n107 a_n17562_12353.n106 0.752
R11042 a_n17562_12353.n9 a_n17562_12353.n48 1.149
R11043 a_n17562_12353.n14 a_n17562_12353.n11 1.148
R11044 a_n17562_12353.n76 a_n17562_12353.n75 0.24
R11045 a_n17562_12353.n136 a_n17562_12353.n135 0.155
R11046 a_n17562_12353.n36 a_n17562_12353.n35 0.155
R11047 a_n17562_12353.n19 a_n17562_12353.n18 0.144
R11048 a_n17562_12353.n40 a_n17562_12353.n39 0.144
R11049 a_n17562_12353.n134 a_n17562_12353.n133 0.133
R11050 a_n17562_12353.n34 a_n17562_12353.n33 0.132
R11051 a_n17562_12353.n54 a_n17562_12353.n52 0.126
R11052 a_n17562_12353.n66 a_n17562_12353.n64 0.126
R11053 a_n17562_12353.n13 a_n17562_12353.n15 0.114
R11054 a_n17562_12353.n14 a_n17562_12353.n12 0.11
R11055 a_n17562_12353.n12 a_n17562_12353.n13 0.107
R11056 a_n17562_12353.n101 a_n17562_12353.n100 0.082
R11057 a_n17562_12353.n77 a_n17562_12353.n82 0.071
R11058 a_n17562_12353.n104 a_n17562_12353.n101 0.042
R11059 a_n17562_12353.n59 a_n17562_12353.n60 0.059
R11060 a_n17562_12353.n8 a_n17562_12353.n50 0.032
R11061 a_n17562_12353.n10 a_n17562_12353.n69 0.032
R11062 a_n17562_12353.n52 a_n17562_12353.n53 0.028
R11063 a_n17562_12353.n48 a_n17562_12353.n49 0.028
R11064 a_n17562_12353.n8 a_n17562_12353.n51 0.028
R11065 a_n17562_12353.n55 a_n17562_12353.n56 0.028
R11066 a_n17562_12353.n57 a_n17562_12353.n58 0.028
R11067 a_n17562_12353.n64 a_n17562_12353.n65 0.028
R11068 a_n17562_12353.n61 a_n17562_12353.n62 0.028
R11069 a_n17562_12353.n71 a_n17562_12353.n72 0.028
R11070 a_n17562_12353.n67 a_n17562_12353.n68 0.028
R11071 a_n17562_12353.n10 a_n17562_12353.n70 0.028
R11072 a_n17562_12353.n74 a_n17562_12353.n73 0.027
R11073 a_n17562_12353.n121 a_n17562_12353.n122 0.024
R11074 a_n17562_12353.n30 a_n17562_12353.n27 0.024
R11075 a_n17562_12353.n130 a_n17562_12353.n127 0.024
R11076 a_n17562_12353.n119 a_n17562_12353.n120 0.147
R11077 a_n17562_12353.n120 a_n17562_12353.n5 0.124
R11078 a_n17562_12353.n117 a_n17562_12353.n14 0.072
R11079 a_n17562_12353.n119 a_n17562_12353.n118 2.702
R11080 a_n17562_12353.n3 a_n17562_12353.n76 0.955
R11081 a_n17562_12353.n0 a_n17562_12353.n104 0.127
R11082 a_n17562_12353.n1 a_n17562_12353.n4 0.11
R11083 a_n17562_12353.n4 a_n17562_12353.n77 0.058
R11084 a_n17562_12353.n100 a_n17562_12353.n2 0.042
R11085 a_n8507_11550.n97 a_n8507_11550.t3 730.676
R11086 a_n8507_11550.n97 a_n8507_11550.t4 395.824
R11087 a_n8507_11550.n50 a_n8507_11550.n49 13.176
R11088 a_n8507_11550.n98 a_n8507_11550.t0 11.725
R11089 a_n8507_11550.n98 a_n8507_11550.t2 10.988
R11090 a_n8507_11550.n137 a_n8507_11550.n39 9.3
R11091 a_n8507_11550.n137 a_n8507_11550.n133 9.3
R11092 a_n8507_11550.n137 a_n8507_11550.n127 9.3
R11093 a_n8507_11550.n137 a_n8507_11550.n58 9.3
R11094 a_n8507_11550.n137 a_n8507_11550.n66 9.3
R11095 a_n8507_11550.n137 a_n8507_11550.n122 9.3
R11096 a_n8507_11550.n137 a_n8507_11550.n117 8.47
R11097 a_n8507_11550.n137 a_n8507_11550.n136 8.469
R11098 a_n8507_11550.n137 a_n8507_11550.n114 8.124
R11099 a_n8507_11550.n137 a_n8507_11550.n29 8.124
R11100 a_n8507_11550.n137 a_n8507_11550.n34 8.097
R11101 a_n8507_11550.n137 a_n8507_11550.n109 8.097
R11102 a_n8507_11550.n137 a_n8507_11550.n61 8.016
R11103 a_n8507_11550.n137 a_n8507_11550.n44 8.016
R11104 a_n8507_11550.n137 a_n8507_11550.n53 7.964
R11105 a_n8507_11550.n137 a_n8507_11550.n48 7.964
R11106 a_n8507_11550.n60 a_n8507_11550.n59 6.4
R11107 a_n8507_11550.n108 a_n8507_11550.n67 6.4
R11108 a_n8507_11550.n32 a_n8507_11550.n31 6.023
R11109 a_n8507_11550.n42 a_n8507_11550.n41 6.023
R11110 a_n8507_11550.n127 a_n8507_11550.n126 6.023
R11111 a_n8507_11550.n47 a_n8507_11550.n46 6.023
R11112 a_n8507_11550.n52 a_n8507_11550.n51 6.023
R11113 a_n8507_11550.n135 a_n8507_11550.n134 5.647
R11114 a_n8507_11550.n58 a_n8507_11550.n55 5.647
R11115 a_n8507_11550.n112 a_n8507_11550.n111 5.647
R11116 a_n8507_11550.n116 a_n8507_11550.n115 5.647
R11117 a_n8507_11550.n124 a_n8507_11550.n123 5.457
R11118 a_n8507_11550.n27 a_n8507_11550.n26 5.27
R11119 a_n8507_11550.n57 a_n8507_11550.n56 5.08
R11120 a_n8507_11550.n39 a_n8507_11550.n38 4.517
R11121 a_n8507_11550.n122 a_n8507_11550.n119 4.517
R11122 a_n8507_11550.n75 a_n8507_11550.n74 4.5
R11123 a_n8507_11550.n2 a_n8507_11550.n1 4.5
R11124 a_n8507_11550.n36 a_n8507_11550.n35 4.314
R11125 a_n8507_11550.n132 a_n8507_11550.n131 4.141
R11126 a_n8507_11550.n63 a_n8507_11550.n62 4.141
R11127 a_n8507_11550.n129 a_n8507_11550.n128 3.944
R11128 a_n8507_11550.n121 a_n8507_11550.n120 3.937
R11129 a_n8507_11550.n65 a_n8507_11550.n64 3.567
R11130 a_n8507_11550.n108 a_n8507_11550.n107 3.033
R11131 a_n8507_11550.t1 a_n8507_11550.n137 2.9
R11132 a_n8507_11550.n133 a_n8507_11550.n132 2.258
R11133 a_n8507_11550.n66 a_n8507_11550.n63 2.258
R11134 a_n8507_11550.n100 a_n8507_11550.n99 1.903
R11135 a_n8507_11550.n38 a_n8507_11550.n37 1.882
R11136 a_n8507_11550.n119 a_n8507_11550.n118 1.882
R11137 a_n8507_11550.n66 a_n8507_11550.n65 1.505
R11138 a_n8507_11550.n94 a_n8507_11550.n101 1.5
R11139 a_n8507_11550.n76 a_n8507_11550.n78 1.5
R11140 a_n8507_11550.n75 a_n8507_11550.n73 1.5
R11141 a_n8507_11550.n21 a_n8507_11550.n24 1.5
R11142 a_n8507_11550.n12 a_n8507_11550.n11 1.5
R11143 a_n8507_11550.n107 a_n8507_11550.n92 1.5
R11144 a_n8507_11550.n99 a_n8507_11550.n98 1.345
R11145 a_n8507_11550.n28 a_n8507_11550.n27 1.129
R11146 a_n8507_11550.n26 a_n8507_11550.n25 1.129
R11147 a_n8507_11550.n133 a_n8507_11550.n129 1.129
R11148 a_n8507_11550.n131 a_n8507_11550.n130 1.129
R11149 a_n8507_11550.n136 a_n8507_11550.n135 0.752
R11150 a_n8507_11550.n55 a_n8507_11550.n54 0.752
R11151 a_n8507_11550.n58 a_n8507_11550.n57 0.752
R11152 a_n8507_11550.n122 a_n8507_11550.n121 0.752
R11153 a_n8507_11550.n111 a_n8507_11550.n110 0.752
R11154 a_n8507_11550.n113 a_n8507_11550.n112 0.752
R11155 a_n8507_11550.n117 a_n8507_11550.n116 0.752
R11156 a_n8507_11550.n99 a_n8507_11550.n97 0.637
R11157 a_n8507_11550.n53 a_n8507_11550.n52 0.536
R11158 a_n8507_11550.n48 a_n8507_11550.n47 0.536
R11159 a_n8507_11550.n61 a_n8507_11550.n60 0.475
R11160 a_n8507_11550.n44 a_n8507_11550.n43 0.475
R11161 a_n8507_11550.n34 a_n8507_11550.n33 0.382
R11162 a_n8507_11550.n109 a_n8507_11550.n108 0.382
R11163 a_n8507_11550.n33 a_n8507_11550.n32 0.376
R11164 a_n8507_11550.n31 a_n8507_11550.n30 0.376
R11165 a_n8507_11550.n39 a_n8507_11550.n36 0.376
R11166 a_n8507_11550.n43 a_n8507_11550.n42 0.376
R11167 a_n8507_11550.n41 a_n8507_11550.n40 0.376
R11168 a_n8507_11550.n127 a_n8507_11550.n124 0.376
R11169 a_n8507_11550.n126 a_n8507_11550.n125 0.376
R11170 a_n8507_11550.n46 a_n8507_11550.n45 0.376
R11171 a_n8507_11550.n51 a_n8507_11550.n50 0.376
R11172 a_n8507_11550.n29 a_n8507_11550.n28 0.349
R11173 a_n8507_11550.n114 a_n8507_11550.n113 0.349
R11174 a_n8507_11550.n94 a_n8507_11550.n93 0.15
R11175 a_n8507_11550.n100 a_n8507_11550.n95 0.148
R11176 a_n8507_11550.n2 a_n8507_11550.n0 0.066
R11177 a_n8507_11550.n84 a_n8507_11550.n83 0.043
R11178 a_n8507_11550.n80 a_n8507_11550.n79 0.043
R11179 a_n8507_11550.n76 a_n8507_11550.n75 0.041
R11180 a_n8507_11550.n91 a_n8507_11550.n90 0.035
R11181 a_n8507_11550.n106 a_n8507_11550.n105 0.035
R11182 a_n8507_11550.n19 a_n8507_11550.n18 0.034
R11183 a_n8507_11550.n23 a_n8507_11550.n22 0.034
R11184 a_n8507_11550.n8 a_n8507_11550.n7 0.034
R11185 a_n8507_11550.n89 a_n8507_11550.n88 0.034
R11186 a_n8507_11550.n104 a_n8507_11550.n103 0.034
R11187 a_n8507_11550.n12 a_n8507_11550.n6 0.032
R11188 a_n8507_11550.n107 a_n8507_11550.n82 0.032
R11189 a_n8507_11550.n9 a_n8507_11550.n8 0.03
R11190 a_n8507_11550.n87 a_n8507_11550.n86 0.03
R11191 a_n8507_11550.n11 a_n8507_11550.n10 0.028
R11192 a_n8507_11550.n72 a_n8507_11550.n70 0.028
R11193 a_n8507_11550.n85 a_n8507_11550.n84 0.028
R11194 a_n8507_11550.n13 a_n8507_11550.n12 0.028
R11195 a_n8507_11550.n69 a_n8507_11550.n68 0.028
R11196 a_n8507_11550.n81 a_n8507_11550.n80 0.028
R11197 a_n8507_11550.n102 a_n8507_11550.n94 0.028
R11198 a_n8507_11550.n17 a_n8507_11550.n15 0.026
R11199 a_n8507_11550.n78 a_n8507_11550.n77 0.026
R11200 a_n8507_11550.n4 a_n8507_11550.n3 0.026
R11201 a_n8507_11550.n18 a_n8507_11550.n17 0.024
R11202 a_n8507_11550.n6 a_n8507_11550.n5 0.024
R11203 a_n8507_11550.n15 a_n8507_11550.n16 0.022
R11204 a_n8507_11550.n5 a_n8507_11550.n4 0.022
R11205 a_n8507_11550.n3 a_n8507_11550.n2 0.022
R11206 a_n8507_11550.n20 a_n8507_11550.n19 0.02
R11207 a_n8507_11550.n10 a_n8507_11550.n9 0.02
R11208 a_n8507_11550.n14 a_n8507_11550.n13 0.02
R11209 a_n8507_11550.n101 a_n8507_11550.n100 0.018
R11210 a_n8507_11550.n82 a_n8507_11550.n81 0.018
R11211 a_n8507_11550.n24 a_n8507_11550.n23 0.017
R11212 a_n8507_11550.n86 a_n8507_11550.n85 0.017
R11213 a_n8507_11550.n70 a_n8507_11550.n71 0.015
R11214 a_n8507_11550.n73 a_n8507_11550.n72 0.015
R11215 a_n8507_11550.n68 a_n8507_11550.n0 0.015
R11216 a_n8507_11550.n75 a_n8507_11550.n69 0.015
R11217 a_n8507_11550.n92 a_n8507_11550.n91 0.013
R11218 a_n8507_11550.n90 a_n8507_11550.n89 0.013
R11219 a_n8507_11550.n107 a_n8507_11550.n106 0.013
R11220 a_n8507_11550.n105 a_n8507_11550.n104 0.013
R11221 a_n8507_11550.n95 a_n8507_11550.n96 0.007
R11222 a_n8507_11550.n21 a_n8507_11550.n20 1.424
R11223 a_n8507_11550.n79 a_n8507_11550.n76 0.005
R11224 a_n8507_11550.n92 a_n8507_11550.n87 0.003
R11225 a_n8507_11550.n103 a_n8507_11550.n102 0.003
R11226 a_n8507_11550.n14 a_n8507_11550.n21 0.47
R11227 a_n9889_12279.n40 a_n9889_12279.t3 732.452
R11228 a_n9889_12279.n40 a_n9889_12279.t2 397.573
R11229 a_n9889_12279.n46 a_n9889_12279.n45 92.5
R11230 a_n9889_12279.n64 a_n9889_12279.n63 92.5
R11231 a_n9889_12279.n45 a_n9889_12279.t1 70.344
R11232 a_n9889_12279.n53 a_n9889_12279.n52 31.034
R11233 a_n9889_12279.n76 a_n9889_12279.n75 31.034
R11234 a_n9889_12279.n1 a_n9889_12279.n57 9.3
R11235 a_n9889_12279.n0 a_n9889_12279.n79 9.3
R11236 a_n9889_12279.n77 a_n9889_12279.n76 9.3
R11237 a_n9889_12279.n54 a_n9889_12279.n53 9.3
R11238 a_n9889_12279.n103 a_n9889_12279.n90 9.154
R11239 a_n9889_12279.n103 a_n9889_12279.n7 9.143
R11240 a_n9889_12279.n103 a_n9889_12279.n6 9.143
R11241 a_n9889_12279.n103 a_n9889_12279.n22 9.132
R11242 a_n9889_12279.n103 a_n9889_12279.n96 9.132
R11243 a_n9889_12279.n103 a_n9889_12279.n100 8.886
R11244 a_n9889_12279.n103 a_n9889_12279.n26 8.885
R11245 a_n9889_12279.n103 a_n9889_12279.n11 8.875
R11246 a_n9889_12279.n103 a_n9889_12279.n32 8.875
R11247 a_n9889_12279.n103 a_n9889_12279.n102 8.864
R11248 a_n9889_12279.n103 a_n9889_12279.n28 8.864
R11249 a_n9889_12279.n47 a_n9889_12279.n46 8.282
R11250 a_n9889_12279.n65 a_n9889_12279.n64 8.282
R11251 a_n9889_12279.t0 a_n9889_12279.n103 7.141
R11252 a_n9889_12279.n54 a_n9889_12279.n50 5.647
R11253 a_n9889_12279.n77 a_n9889_12279.n73 5.647
R11254 a_n9889_12279.n84 a_n9889_12279.n83 4.723
R11255 a_n9889_12279.n2 a_n9889_12279.n62 4.65
R11256 a_n9889_12279.n90 a_n9889_12279.n85 4.65
R11257 a_n9889_12279.n83 a_n9889_12279.n3 4.566
R11258 a_n9889_12279.n90 a_n9889_12279.n39 4.517
R11259 a_n9889_12279.n66 a_n9889_12279.n65 4.5
R11260 a_n9889_12279.n67 a_n9889_12279.n69 4.5
R11261 a_n9889_12279.n43 a_n9889_12279.n47 4.5
R11262 a_n9889_12279.n70 a_n9889_12279.n78 4.5
R11263 a_n9889_12279.n2 a_n9889_12279.n61 4.5
R11264 a_n9889_12279.n4 a_n9889_12279.n56 4.5
R11265 a_n9889_12279.n0 a_n9889_12279.n82 4.5
R11266 a_n9889_12279.n1 a_n9889_12279.n60 4.5
R11267 a_n9889_12279.n98 a_n9889_12279.n97 4.141
R11268 a_n9889_12279.n90 a_n9889_12279.n38 4.141
R11269 a_n9889_12279.n24 a_n9889_12279.n23 4.141
R11270 a_n9889_12279.n52 a_n9889_12279.n51 4.137
R11271 a_n9889_12279.n75 a_n9889_12279.n74 4.137
R11272 a_n9889_12279.n60 a_n9889_12279.n58 3.764
R11273 a_n9889_12279.n78 a_n9889_12279.n71 3.764
R11274 a_n9889_12279.n92 a_n9889_12279.n91 3.764
R11275 a_n9889_12279.n7 a_n9889_12279.n34 3.764
R11276 a_n9889_12279.n96 a_n9889_12279.n95 3.736
R11277 a_n9889_12279.n56 a_n9889_12279.n55 3.388
R11278 a_n9889_12279.n82 a_n9889_12279.n81 3.388
R11279 a_n9889_12279.n9 a_n9889_12279.n8 3.388
R11280 a_n9889_12279.n6 a_n9889_12279.n13 3.388
R11281 a_n9889_12279.n18 a_n9889_12279.n17 3.388
R11282 a_n9889_12279.n30 a_n9889_12279.n29 3.388
R11283 a_n9889_12279.n22 a_n9889_12279.n21 3.36
R11284 a_n9889_12279.n56 a_n9889_12279.n54 3.011
R11285 a_n9889_12279.n47 a_n9889_12279.n44 3.011
R11286 a_n9889_12279.n82 a_n9889_12279.n80 3.011
R11287 a_n9889_12279.n10 a_n9889_12279.n9 3.011
R11288 a_n9889_12279.n13 a_n9889_12279.n12 3.011
R11289 a_n9889_12279.n16 a_n9889_12279.n15 3.011
R11290 a_n9889_12279.n21 a_n9889_12279.n20 3.011
R11291 a_n9889_12279.n19 a_n9889_12279.n18 3.011
R11292 a_n9889_12279.n31 a_n9889_12279.n30 3.011
R11293 a_n9889_12279.n60 a_n9889_12279.n59 2.635
R11294 a_n9889_12279.n69 a_n9889_12279.n68 2.635
R11295 a_n9889_12279.n78 a_n9889_12279.n77 2.635
R11296 a_n9889_12279.n93 a_n9889_12279.n92 2.635
R11297 a_n9889_12279.n95 a_n9889_12279.n94 2.635
R11298 a_n9889_12279.n37 a_n9889_12279.n36 2.635
R11299 a_n9889_12279.n34 a_n9889_12279.n33 2.635
R11300 a_n9889_12279.n83 a_n9889_12279.n40 2.35
R11301 a_n9889_12279.n99 a_n9889_12279.n98 2.258
R11302 a_n9889_12279.n25 a_n9889_12279.n24 2.258
R11303 a_n9889_12279.n5 a_n9889_12279.n89 1.619
R11304 a_n9889_12279.n86 a_n9889_12279.n87 1.588
R11305 a_n9889_12279.n5 a_n9889_12279.n104 1.88
R11306 a_n9889_12279.n3 a_n9889_12279.n0 2.375
R11307 a_n9889_12279.n7 a_n9889_12279.n37 2.257
R11308 a_n9889_12279.n6 a_n9889_12279.n16 2.257
R11309 a_n9889_12279.n36 a_n9889_12279.n35 1.505
R11310 a_n9889_12279.n42 a_n9889_12279.n1 1.5
R11311 a_n9889_12279.n15 a_n9889_12279.n14 1.129
R11312 a_n9889_12279.n50 a_n9889_12279.n49 0.752
R11313 a_n9889_12279.n73 a_n9889_12279.n72 0.752
R11314 a_n9889_12279.n42 a_n9889_12279.n41 0.24
R11315 a_n9889_12279.n102 a_n9889_12279.n101 0.155
R11316 a_n9889_12279.n28 a_n9889_12279.n27 0.155
R11317 a_n9889_12279.n11 a_n9889_12279.n10 0.144
R11318 a_n9889_12279.n32 a_n9889_12279.n31 0.144
R11319 a_n9889_12279.n100 a_n9889_12279.n99 0.133
R11320 a_n9889_12279.n26 a_n9889_12279.n25 0.132
R11321 a_n9889_12279.n67 a_n9889_12279.n66 0.082
R11322 a_n9889_12279.n43 a_n9889_12279.n48 0.071
R11323 a_n9889_12279.n70 a_n9889_12279.n67 0.042
R11324 a_n9889_12279.n87 a_n9889_12279.n88 0.024
R11325 a_n9889_12279.n22 a_n9889_12279.n19 0.024
R11326 a_n9889_12279.n96 a_n9889_12279.n93 0.024
R11327 a_n9889_12279.n85 a_n9889_12279.n86 0.147
R11328 a_n9889_12279.n86 a_n9889_12279.n5 0.124
R11329 a_n9889_12279.n85 a_n9889_12279.n84 2.702
R11330 a_n9889_12279.n3 a_n9889_12279.n42 0.955
R11331 a_n9889_12279.n0 a_n9889_12279.n70 0.127
R11332 a_n9889_12279.n1 a_n9889_12279.n4 0.11
R11333 a_n9889_12279.n4 a_n9889_12279.n43 0.058
R11334 a_n9889_12279.n66 a_n9889_12279.n2 0.042
R11335 a_n18722_2907.n95 a_n18722_2907.t3 730.679
R11336 a_n18722_2907.n95 a_n18722_2907.t4 395.833
R11337 a_n18722_2907.n41 a_n18722_2907.n40 13.176
R11338 a_n18722_2907.n96 a_n18722_2907.t1 11.724
R11339 a_n18722_2907.n96 a_n18722_2907.t0 10.997
R11340 a_n18722_2907.n150 a_n18722_2907.n34 9.3
R11341 a_n18722_2907.n150 a_n18722_2907.n141 9.3
R11342 a_n18722_2907.n150 a_n18722_2907.n135 9.3
R11343 a_n18722_2907.n150 a_n18722_2907.n49 9.3
R11344 a_n18722_2907.n150 a_n18722_2907.n54 9.3
R11345 a_n18722_2907.n150 a_n18722_2907.n123 9.3
R11346 a_n18722_2907.n150 a_n18722_2907.n149 8.469
R11347 a_n18722_2907.n150 a_n18722_2907.n113 8.469
R11348 a_n18722_2907.n150 a_n18722_2907.n118 8.125
R11349 a_n18722_2907.n150 a_n18722_2907.n29 8.124
R11350 a_n18722_2907.n150 a_n18722_2907.n110 8.097
R11351 a_n18722_2907.n150 a_n18722_2907.n146 8.096
R11352 a_n18722_2907.n150 a_n18722_2907.n126 8.016
R11353 a_n18722_2907.n150 a_n18722_2907.n39 8.016
R11354 a_n18722_2907.n150 a_n18722_2907.n130 7.964
R11355 a_n18722_2907.n150 a_n18722_2907.n44 7.964
R11356 a_n18722_2907.n125 a_n18722_2907.n124 6.4
R11357 a_n18722_2907.n109 a_n18722_2907.n55 6.4
R11358 a_n18722_2907.n144 a_n18722_2907.n143 6.023
R11359 a_n18722_2907.n37 a_n18722_2907.n36 6.023
R11360 a_n18722_2907.n135 a_n18722_2907.n134 6.023
R11361 a_n18722_2907.n43 a_n18722_2907.n42 6.023
R11362 a_n18722_2907.n129 a_n18722_2907.n128 6.023
R11363 a_n18722_2907.n148 a_n18722_2907.n147 5.647
R11364 a_n18722_2907.n49 a_n18722_2907.n46 5.647
R11365 a_n18722_2907.n116 a_n18722_2907.n115 5.647
R11366 a_n18722_2907.n112 a_n18722_2907.n111 5.647
R11367 a_n18722_2907.n132 a_n18722_2907.n131 5.457
R11368 a_n18722_2907.n27 a_n18722_2907.n26 5.27
R11369 a_n18722_2907.n48 a_n18722_2907.n47 5.08
R11370 a_n18722_2907.n34 a_n18722_2907.n33 4.517
R11371 a_n18722_2907.n123 a_n18722_2907.n120 4.517
R11372 a_n18722_2907.n63 a_n18722_2907.n62 4.5
R11373 a_n18722_2907.n2 a_n18722_2907.n1 4.5
R11374 a_n18722_2907.n31 a_n18722_2907.n30 4.314
R11375 a_n18722_2907.n140 a_n18722_2907.n139 4.141
R11376 a_n18722_2907.n51 a_n18722_2907.n50 4.141
R11377 a_n18722_2907.n137 a_n18722_2907.n136 3.944
R11378 a_n18722_2907.n122 a_n18722_2907.n121 3.937
R11379 a_n18722_2907.n53 a_n18722_2907.n52 3.567
R11380 a_n18722_2907.n109 a_n18722_2907.n108 3.033
R11381 a_n18722_2907.t2 a_n18722_2907.n150 2.9
R11382 a_n18722_2907.n141 a_n18722_2907.n140 2.258
R11383 a_n18722_2907.n54 a_n18722_2907.n51 2.258
R11384 a_n18722_2907.n33 a_n18722_2907.n32 1.882
R11385 a_n18722_2907.n120 a_n18722_2907.n119 1.882
R11386 a_n18722_2907.n98 a_n18722_2907.n97 1.657
R11387 a_n18722_2907.n54 a_n18722_2907.n53 1.505
R11388 a_n18722_2907.n82 a_n18722_2907.n102 1.5
R11389 a_n18722_2907.n64 a_n18722_2907.n66 1.5
R11390 a_n18722_2907.n63 a_n18722_2907.n61 1.5
R11391 a_n18722_2907.n21 a_n18722_2907.n24 1.5
R11392 a_n18722_2907.n12 a_n18722_2907.n11 1.5
R11393 a_n18722_2907.n108 a_n18722_2907.n80 1.5
R11394 a_n18722_2907.n97 a_n18722_2907.n96 1.221
R11395 a_n18722_2907.n28 a_n18722_2907.n27 1.129
R11396 a_n18722_2907.n26 a_n18722_2907.n25 1.129
R11397 a_n18722_2907.n141 a_n18722_2907.n137 1.129
R11398 a_n18722_2907.n139 a_n18722_2907.n138 1.129
R11399 a_n18722_2907.n101 a_n18722_2907.n100 0.853
R11400 a_n18722_2907.n149 a_n18722_2907.n148 0.752
R11401 a_n18722_2907.n46 a_n18722_2907.n45 0.752
R11402 a_n18722_2907.n49 a_n18722_2907.n48 0.752
R11403 a_n18722_2907.n123 a_n18722_2907.n122 0.752
R11404 a_n18722_2907.n115 a_n18722_2907.n114 0.752
R11405 a_n18722_2907.n117 a_n18722_2907.n116 0.752
R11406 a_n18722_2907.n113 a_n18722_2907.n112 0.752
R11407 a_n18722_2907.n89 a_n18722_2907.n88 0.716
R11408 a_n18722_2907.n97 a_n18722_2907.n95 0.637
R11409 a_n18722_2907.n130 a_n18722_2907.n129 0.536
R11410 a_n18722_2907.n44 a_n18722_2907.n43 0.536
R11411 a_n18722_2907.n126 a_n18722_2907.n125 0.476
R11412 a_n18722_2907.n39 a_n18722_2907.n38 0.475
R11413 a_n18722_2907.n110 a_n18722_2907.n109 0.382
R11414 a_n18722_2907.n146 a_n18722_2907.n145 0.382
R11415 a_n18722_2907.n145 a_n18722_2907.n144 0.376
R11416 a_n18722_2907.n143 a_n18722_2907.n142 0.376
R11417 a_n18722_2907.n34 a_n18722_2907.n31 0.376
R11418 a_n18722_2907.n38 a_n18722_2907.n37 0.376
R11419 a_n18722_2907.n36 a_n18722_2907.n35 0.376
R11420 a_n18722_2907.n135 a_n18722_2907.n132 0.376
R11421 a_n18722_2907.n134 a_n18722_2907.n133 0.376
R11422 a_n18722_2907.n42 a_n18722_2907.n41 0.376
R11423 a_n18722_2907.n128 a_n18722_2907.n127 0.376
R11424 a_n18722_2907.n118 a_n18722_2907.n117 0.35
R11425 a_n18722_2907.n29 a_n18722_2907.n28 0.349
R11426 a_n18722_2907.n2 a_n18722_2907.n0 0.066
R11427 a_n18722_2907.n87 a_n18722_2907.n86 0.047
R11428 a_n18722_2907.n72 a_n18722_2907.n71 0.043
R11429 a_n18722_2907.n68 a_n18722_2907.n67 0.043
R11430 a_n18722_2907.n64 a_n18722_2907.n63 0.041
R11431 a_n18722_2907.n79 a_n18722_2907.n78 0.035
R11432 a_n18722_2907.n107 a_n18722_2907.n106 0.035
R11433 a_n18722_2907.n19 a_n18722_2907.n18 0.034
R11434 a_n18722_2907.n23 a_n18722_2907.n22 0.034
R11435 a_n18722_2907.n8 a_n18722_2907.n7 0.034
R11436 a_n18722_2907.n77 a_n18722_2907.n76 0.034
R11437 a_n18722_2907.n105 a_n18722_2907.n104 0.034
R11438 a_n18722_2907.n12 a_n18722_2907.n6 0.032
R11439 a_n18722_2907.n108 a_n18722_2907.n70 0.032
R11440 a_n18722_2907.n99 a_n18722_2907.n98 0.031
R11441 a_n18722_2907.n9 a_n18722_2907.n8 0.03
R11442 a_n18722_2907.n75 a_n18722_2907.n74 0.03
R11443 a_n18722_2907.n101 a_n18722_2907.n94 0.03
R11444 a_n18722_2907.n81 a_n18722_2907.n87 0.03
R11445 a_n18722_2907.n11 a_n18722_2907.n10 0.028
R11446 a_n18722_2907.n60 a_n18722_2907.n58 0.028
R11447 a_n18722_2907.n73 a_n18722_2907.n72 0.028
R11448 a_n18722_2907.n91 a_n18722_2907.n90 0.028
R11449 a_n18722_2907.n13 a_n18722_2907.n12 0.028
R11450 a_n18722_2907.n57 a_n18722_2907.n56 0.028
R11451 a_n18722_2907.n69 a_n18722_2907.n68 0.028
R11452 a_n18722_2907.n103 a_n18722_2907.n82 0.028
R11453 a_n18722_2907.n85 a_n18722_2907.n83 0.028
R11454 a_n18722_2907.n17 a_n18722_2907.n15 0.026
R11455 a_n18722_2907.n66 a_n18722_2907.n65 0.026
R11456 a_n18722_2907.n93 a_n18722_2907.n92 0.026
R11457 a_n18722_2907.n4 a_n18722_2907.n3 0.026
R11458 a_n18722_2907.n90 a_n18722_2907.n89 0.024
R11459 a_n18722_2907.n18 a_n18722_2907.n17 0.024
R11460 a_n18722_2907.n6 a_n18722_2907.n5 0.024
R11461 a_n18722_2907.n15 a_n18722_2907.n16 0.022
R11462 a_n18722_2907.n5 a_n18722_2907.n4 0.022
R11463 a_n18722_2907.n3 a_n18722_2907.n2 0.022
R11464 a_n18722_2907.n20 a_n18722_2907.n19 0.02
R11465 a_n18722_2907.n10 a_n18722_2907.n9 0.02
R11466 a_n18722_2907.n94 a_n18722_2907.n93 0.02
R11467 a_n18722_2907.n14 a_n18722_2907.n13 0.02
R11468 a_n18722_2907.n100 a_n18722_2907.n99 0.019
R11469 a_n18722_2907.n82 a_n18722_2907.n81 0.018
R11470 a_n18722_2907.n102 a_n18722_2907.n101 0.018
R11471 a_n18722_2907.n70 a_n18722_2907.n69 0.018
R11472 a_n18722_2907.n24 a_n18722_2907.n23 0.017
R11473 a_n18722_2907.n74 a_n18722_2907.n73 0.017
R11474 a_n18722_2907.n58 a_n18722_2907.n59 0.015
R11475 a_n18722_2907.n61 a_n18722_2907.n60 0.015
R11476 a_n18722_2907.n56 a_n18722_2907.n0 0.015
R11477 a_n18722_2907.n63 a_n18722_2907.n57 0.015
R11478 a_n18722_2907.n80 a_n18722_2907.n79 0.013
R11479 a_n18722_2907.n78 a_n18722_2907.n77 0.013
R11480 a_n18722_2907.n108 a_n18722_2907.n107 0.013
R11481 a_n18722_2907.n106 a_n18722_2907.n105 0.013
R11482 a_n18722_2907.n92 a_n18722_2907.n91 0.007
R11483 a_n18722_2907.n86 a_n18722_2907.n85 0.007
R11484 a_n18722_2907.n21 a_n18722_2907.n20 1.424
R11485 a_n18722_2907.n67 a_n18722_2907.n64 0.005
R11486 a_n18722_2907.n80 a_n18722_2907.n75 0.003
R11487 a_n18722_2907.n104 a_n18722_2907.n103 0.003
R11488 a_n18722_2907.n83 a_n18722_2907.n84 0.003
R11489 a_n18722_2907.n14 a_n18722_2907.n21 0.47
R11490 a_n18744_6000.n13 a_n18744_6000.t2 732.456
R11491 a_n18744_6000.n13 a_n18744_6000.t3 397.58
R11492 a_n18744_6000.n51 a_n18744_6000.n50 92.5
R11493 a_n18744_6000.n9 a_n18744_6000.n8 92.5
R11494 a_n18744_6000.n50 a_n18744_6000.t1 70.344
R11495 a_n18744_6000.n45 a_n18744_6000.n44 31.034
R11496 a_n18744_6000.n24 a_n18744_6000.n23 31.034
R11497 a_n18744_6000.n27 a_n18744_6000.n28 9.3
R11498 a_n18744_6000.n38 a_n18744_6000.n39 9.3
R11499 a_n18744_6000.n46 a_n18744_6000.n45 9.3
R11500 a_n18744_6000.n25 a_n18744_6000.n24 9.3
R11501 a_n18744_6000.n105 a_n18744_6000.n98 9.154
R11502 a_n18744_6000.n105 a_n18744_6000.n4 9.143
R11503 a_n18744_6000.n105 a_n18744_6000.n3 9.143
R11504 a_n18744_6000.n105 a_n18744_6000.n78 9.132
R11505 a_n18744_6000.n105 a_n18744_6000.n62 9.132
R11506 a_n18744_6000.n105 a_n18744_6000.n102 8.885
R11507 a_n18744_6000.n105 a_n18744_6000.n82 8.885
R11508 a_n18744_6000.n105 a_n18744_6000.n86 8.875
R11509 a_n18744_6000.n105 a_n18744_6000.n56 8.875
R11510 a_n18744_6000.n105 a_n18744_6000.n104 8.864
R11511 a_n18744_6000.n105 a_n18744_6000.n88 8.864
R11512 a_n18744_6000.n52 a_n18744_6000.n51 8.282
R11513 a_n18744_6000.n10 a_n18744_6000.n9 8.282
R11514 a_n18744_6000.t0 a_n18744_6000.n105 7.141
R11515 a_n18744_6000.n46 a_n18744_6000.n42 5.647
R11516 a_n18744_6000.n25 a_n18744_6000.n21 5.647
R11517 a_n18744_6000.n1 a_n18744_6000.n11 4.65
R11518 a_n18744_6000.n16 a_n18744_6000.n15 4.566
R11519 a_n18744_6000.n98 a_n18744_6000.n90 4.517
R11520 a_n18744_6000.n0 a_n18744_6000.n10 4.5
R11521 a_n18744_6000.n1 a_n18744_6000.n7 4.5
R11522 a_n18744_6000.n6 a_n18744_6000.n52 4.5
R11523 a_n18744_6000.n40 a_n18744_6000.n48 4.5
R11524 a_n18744_6000.n12 a_n18744_6000.n37 4.5
R11525 a_n18744_6000.n17 a_n18744_6000.n32 4.5
R11526 a_n18744_6000.n15 a_n18744_6000.n14 4.482
R11527 a_n18744_6000.n100 a_n18744_6000.n99 4.141
R11528 a_n18744_6000.n98 a_n18744_6000.n89 4.141
R11529 a_n18744_6000.n80 a_n18744_6000.n79 4.141
R11530 a_n18744_6000.n44 a_n18744_6000.n43 4.137
R11531 a_n18744_6000.n23 a_n18744_6000.n22 4.137
R11532 a_n18744_6000.n37 a_n18744_6000.n35 3.764
R11533 a_n18744_6000.n26 a_n18744_6000.n19 3.764
R11534 a_n18744_6000.n58 a_n18744_6000.n57 3.764
R11535 a_n18744_6000.n3 a_n18744_6000.n69 3.764
R11536 a_n18744_6000.n62 a_n18744_6000.n61 3.736
R11537 a_n18744_6000.n48 a_n18744_6000.n47 3.388
R11538 a_n18744_6000.n32 a_n18744_6000.n31 3.388
R11539 a_n18744_6000.n54 a_n18744_6000.n53 3.388
R11540 a_n18744_6000.n4 a_n18744_6000.n67 3.388
R11541 a_n18744_6000.n76 a_n18744_6000.n75 3.388
R11542 a_n18744_6000.n84 a_n18744_6000.n83 3.388
R11543 a_n18744_6000.n78 a_n18744_6000.n74 3.36
R11544 a_n18744_6000.n48 a_n18744_6000.n46 3.011
R11545 a_n18744_6000.n52 a_n18744_6000.n49 3.011
R11546 a_n18744_6000.n32 a_n18744_6000.n30 3.011
R11547 a_n18744_6000.n55 a_n18744_6000.n54 3.011
R11548 a_n18744_6000.n67 a_n18744_6000.n66 3.011
R11549 a_n18744_6000.n65 a_n18744_6000.n64 3.011
R11550 a_n18744_6000.n74 a_n18744_6000.n73 3.011
R11551 a_n18744_6000.n77 a_n18744_6000.n76 3.011
R11552 a_n18744_6000.n85 a_n18744_6000.n84 3.011
R11553 a_n18744_6000.n91 a_n18744_6000.n14 2.921
R11554 a_n18744_6000.n37 a_n18744_6000.n36 2.635
R11555 a_n18744_6000.n26 a_n18744_6000.n25 2.635
R11556 a_n18744_6000.n59 a_n18744_6000.n58 2.635
R11557 a_n18744_6000.n61 a_n18744_6000.n60 2.635
R11558 a_n18744_6000.n72 a_n18744_6000.n71 2.635
R11559 a_n18744_6000.n69 a_n18744_6000.n68 2.635
R11560 a_n18744_6000.n15 a_n18744_6000.n13 2.349
R11561 a_n18744_6000.n101 a_n18744_6000.n100 2.258
R11562 a_n18744_6000.n81 a_n18744_6000.n80 2.258
R11563 a_n18744_6000.n5 a_n18744_6000.n96 1.633
R11564 a_n18744_6000.n2 a_n18744_6000.n95 1.619
R11565 a_n18744_6000.n92 a_n18744_6000.n93 1.588
R11566 a_n18744_6000.n5 a_n18744_6000.n106 1.587
R11567 a_n18744_6000.n71 a_n18744_6000.n70 1.505
R11568 a_n18744_6000.n12 a_n18744_6000.n34 1.5
R11569 a_n18744_6000.n64 a_n18744_6000.n63 1.129
R11570 a_n18744_6000.n42 a_n18744_6000.n41 0.752
R11571 a_n18744_6000.n21 a_n18744_6000.n20 0.752
R11572 a_n18744_6000.n104 a_n18744_6000.n103 0.155
R11573 a_n18744_6000.n88 a_n18744_6000.n87 0.155
R11574 a_n18744_6000.n56 a_n18744_6000.n55 0.144
R11575 a_n18744_6000.n86 a_n18744_6000.n85 0.144
R11576 a_n18744_6000.n102 a_n18744_6000.n101 0.132
R11577 a_n18744_6000.n82 a_n18744_6000.n81 0.132
R11578 a_n18744_6000.n91 a_n18744_6000.n92 0.125
R11579 a_n18744_6000.n106 a_n18744_6000.n107 0.037
R11580 a_n18744_6000.n96 a_n18744_6000.n97 0.034
R11581 a_n18744_6000.n40 a_n18744_6000.n38 0.094
R11582 a_n18744_6000.n34 a_n18744_6000.n33 0.293
R11583 a_n18744_6000.n34 a_n18744_6000.n18 0.877
R11584 a_n18744_6000.n93 a_n18744_6000.n94 0.024
R11585 a_n18744_6000.n62 a_n18744_6000.n59 0.024
R11586 a_n18744_6000.n78 a_n18744_6000.n77 0.024
R11587 a_n18744_6000.n98 a_n18744_6000.n91 4.672
R11588 a_n18744_6000.n18 a_n18744_6000.n16 0.019
R11589 a_n18744_6000.n18 a_n18744_6000.n17 2.433
R11590 a_n18744_6000.n6 a_n18744_6000.n40 0.044
R11591 a_n18744_6000.n17 a_n18744_6000.n27 0.032
R11592 a_n18744_6000.n38 a_n18744_6000.n12 0.031
R11593 a_n18744_6000.n17 a_n18744_6000.n29 0.017
R11594 a_n18744_6000.n27 a_n18744_6000.n26 4.595
R11595 a_n18744_6000.n4 a_n18744_6000.n65 2.257
R11596 a_n18744_6000.n3 a_n18744_6000.n72 2.257
R11597 a_n18744_6000.n2 a_n18744_6000.n5 0.256
R11598 a_n18744_6000.n92 a_n18744_6000.n2 0.124
R11599 a_n18744_6000.n6 a_n18744_6000.n1 0.07
R11600 a_n18744_6000.n1 a_n18744_6000.n0 0.053
R11601 modi1.n266 modi1.t4 1037.94
R11602 modi1.n257 modi1.t3 1037.29
R11603 modi1.n257 modi1.t5 797.574
R11604 modi1.n266 modi1.t2 796.922
R11605 modi1.n30 modi1.n29 92.5
R11606 modi1.n46 modi1.n45 92.5
R11607 modi1.n45 modi1.t1 70.344
R11608 modi1.n8 modi1.n7 31.034
R11609 modi1.n65 modi1.n64 31.034
R11610 modi1.n113 modi1.n112 9.3
R11611 modi1.n190 modi1.n189 9.3
R11612 modi1.n15 modi1.n14 9.3
R11613 modi1.n66 modi1.n65 9.3
R11614 modi1.n9 modi1.n8 9.3
R11615 modi1.n77 modi1.n76 9.3
R11616 modi1.n229 modi1.n228 9.154
R11617 modi1.n31 modi1.n30 8.282
R11618 modi1.n47 modi1.n46 8.282
R11619 modi1.n228 modi1.t0 7.141
R11620 modi1.n149 modi1.n148 7.033
R11621 modi1.n92 modi1.n91 7.033
R11622 modi1.n258 modi1.n256 6.465
R11623 modi1.n9 modi1.n5 5.647
R11624 modi1.n66 modi1.n62 5.647
R11625 modi1.n230 modi1.n229 4.65
R11626 modi1.n44 modi1.n43 4.65
R11627 modi1.n176 modi1.n175 4.5
R11628 modi1.n196 modi1.n195 4.5
R11629 modi1.n209 modi1.n208 4.5
R11630 modi1.n216 modi1.n213 4.5
R11631 modi1.n225 modi1.n224 4.5
R11632 modi1.n231 modi1.n227 4.5
R11633 modi1.n100 modi1.n97 4.5
R11634 modi1.n107 modi1.n106 4.5
R11635 modi1.n119 modi1.n118 4.5
R11636 modi1.n129 modi1.n128 4.5
R11637 modi1.n139 modi1.n138 4.5
R11638 modi1.n163 modi1.n162 4.5
R11639 modi1.n83 modi1.n81 4.5
R11640 modi1.n70 modi1.n67 4.5
R11641 modi1.n57 modi1.n55 4.5
R11642 modi1.n32 modi1.n31 4.5
R11643 modi1.n39 modi1.n38 4.5
R11644 modi1.n48 modi1.n47 4.5
R11645 modi1.n12 modi1.n11 4.5
R11646 modi1.n20 modi1.n19 4.5
R11647 modi1.n128 modi1.n125 4.141
R11648 modi1.n162 modi1.n161 4.141
R11649 modi1.n7 modi1.n6 4.137
R11650 modi1.n64 modi1.n63 4.137
R11651 modi1.n118 modi1.n115 3.764
R11652 modi1.n208 modi1.n206 3.764
R11653 modi1.n19 modi1.n17 3.764
R11654 modi1.n67 modi1.n60 3.764
R11655 modi1.n271 modi1.n266 3.463
R11656 modi1.n138 modi1.n135 3.388
R11657 modi1.n106 modi1.n105 3.388
R11658 modi1.n195 modi1.n194 3.388
R11659 modi1.n175 modi1.n174 3.388
R11660 modi1.n11 modi1.n10 3.388
R11661 modi1.n81 modi1.n80 3.388
R11662 modi1 modi1.n258 3.022
R11663 modi1.n138 modi1.n137 3.011
R11664 modi1.n106 modi1.n103 3.011
R11665 modi1.n97 modi1.n95 3.011
R11666 modi1.n189 modi1.n188 3.011
R11667 modi1.n195 modi1.n193 3.011
R11668 modi1.n175 modi1.n173 3.011
R11669 modi1.n11 modi1.n9 3.011
R11670 modi1.n31 modi1.n28 3.011
R11671 modi1.n81 modi1.n79 3.011
R11672 modi1.n118 modi1.n117 2.635
R11673 modi1.n112 modi1.n111 2.635
R11674 modi1.n213 modi1.n212 2.635
R11675 modi1.n208 modi1.n207 2.635
R11676 modi1.n19 modi1.n18 2.635
R11677 modi1.n55 modi1.n54 2.635
R11678 modi1.n67 modi1.n66 2.635
R11679 modi1.n128 modi1.n127 2.258
R11680 modi1.n162 modi1.n160 2.258
R11681 modi1.n258 modi1.n257 2.25
R11682 modi1.n25 modi1.n0 1.754
R11683 modi1.n179 modi1.n150 1.754
R11684 modi1.n25 modi1.n24 1.705
R11685 modi1.n42 modi1.n41 1.705
R11686 modi1.n72 modi1.n71 1.705
R11687 modi1.n86 modi1.n85 1.705
R11688 modi1.n255 modi1.n144 1.705
R11689 modi1.n199 modi1.n198 1.705
R11690 modi1.n219 modi1.n218 1.705
R11691 modi1.n248 modi1.n247 1.705
R11692 modi1.n254 modi1.n253 1.705
R11693 modi1.n242 modi1.n241 1.705
R11694 modi1.n236 modi1.n235 1.705
R11695 modi1.n185 modi1.n184 1.705
R11696 modi1.n179 modi1.n178 1.705
R11697 modi1.n213 modi1.n211 1.505
R11698 modi1.n197 modi1.n196 1.5
R11699 modi1.n210 modi1.n209 1.5
R11700 modi1.n217 modi1.n216 1.5
R11701 modi1.n226 modi1.n225 1.5
R11702 modi1.n232 modi1.n231 1.5
R11703 modi1.n84 modi1.n83 1.5
R11704 modi1.n71 modi1.n70 1.5
R11705 modi1.n33 modi1.n32 1.5
R11706 modi1.n58 modi1.n57 1.5
R11707 modi1.n40 modi1.n39 1.5
R11708 modi1.n49 modi1.n48 1.5
R11709 modi1.n24 modi1.n12 1.5
R11710 modi1.n21 modi1.n20 1.5
R11711 modi1.n287 modi1.n286 1.402
R11712 modi1.n272 modi1.n271 1.355
R11713 modi1.n256 modi1.n255 1.268
R11714 modi1.n288 modi1.n287 1.141
R11715 modi1.n289 modi1.n288 1.137
R11716 modi1.n279 modi1.n278 1.137
R11717 modi1.n294 modi1.n293 1.137
R11718 modi1.n273 modi1.n272 1.137
R11719 modi1.n263 modi1.n262 1.137
R11720 modi1.n298 modi1.n297 1.137
R11721 modi1.n300 modi1.n299 1.136
R11722 modi1.n275 modi1.n274 1.136
R11723 modi1.n97 modi1.n96 1.129
R11724 modi1.n150 modi1.n149 1.127
R11725 modi1.n144 modi1.n92 1.127
R11726 modi1.n140 modi1.n139 1.125
R11727 modi1.n177 modi1.n176 1.125
R11728 modi1.n5 modi1.n4 0.752
R11729 modi1.n62 modi1.n61 0.752
R11730 modi1.n256 modi1.n86 0.709
R11731 modi1.n91 modi1.n90 0.155
R11732 modi1.n148 modi1.n147 0.155
R11733 modi1.n137 modi1.n136 0.144
R11734 modi1.n173 modi1.n172 0.144
R11735 modi1.n127 modi1.n126 0.133
R11736 modi1.n160 modi1.n159 0.132
R11737 modi1.n133 modi1.n132 0.053
R11738 modi1.n123 modi1.n122 0.053
R11739 modi1.n113 modi1.n110 0.053
R11740 modi1.n157 modi1.n156 0.053
R11741 modi1.n167 modi1.n166 0.053
R11742 modi1.n170 modi1.n169 0.053
R11743 modi1.n77 modi1.n75 0.053
R11744 modi1.n42 modi1.n25 0.049
R11745 modi1.n72 modi1.n42 0.049
R11746 modi1.n86 modi1.n72 0.049
R11747 modi1.n255 modi1.n254 0.049
R11748 modi1.n254 modi1.n248 0.049
R11749 modi1.n248 modi1.n242 0.049
R11750 modi1.n242 modi1.n236 0.049
R11751 modi1.n236 modi1.n219 0.049
R11752 modi1.n219 modi1.n199 0.049
R11753 modi1.n199 modi1.n185 0.049
R11754 modi1.n185 modi1.n179 0.049
R11755 modi1.n271 modi1.n270 0.048
R11756 modi1.n39 modi1.n37 0.045
R11757 modi1.n57 modi1.n53 0.045
R11758 modi1.n100 modi1.n99 0.043
R11759 modi1.n225 modi1.n223 0.043
R11760 modi1.n88 modi1.n87 0.034
R11761 modi1.n166 modi1.n165 0.032
R11762 modi1.n134 modi1.n133 0.03
R11763 modi1.n132 modi1.n131 0.03
R11764 modi1.n156 modi1.n155 0.03
R11765 modi1.n22 modi1.n21 0.03
R11766 modi1.n84 modi1.n74 0.03
R11767 modi1.n122 modi1.n121 0.028
R11768 modi1.n168 modi1.n167 0.028
R11769 modi1.n171 modi1.n170 0.028
R11770 modi1.n94 modi1.n93 0.025
R11771 modi1.n124 modi1.n123 0.025
R11772 modi1.n48 modi1.n44 0.025
R11773 modi1.n117 modi1.n116 0.024
R11774 modi1.n193 modi1.n192 0.024
R11775 modi1.n231 modi1.n230 0.023
R11776 modi1.n158 modi1.n157 0.023
R11777 modi1.n120 modi1.n119 0.021
R11778 modi1.n114 modi1.n113 0.021
R11779 modi1.n203 modi1.n202 0.021
R11780 modi1.n20 modi1.n13 0.021
R11781 modi1.n16 modi1.n15 0.021
R11782 modi1.n70 modi1.n59 0.021
R11783 modi1.n293 modi1.n292 0.021
R11784 modi1.n139 modi1.n94 0.019
R11785 modi1.n110 modi1.n109 0.019
R11786 modi1.n109 modi1.n108 0.019
R11787 modi1.n107 modi1.n102 0.019
R11788 modi1.n204 modi1.n203 0.019
R11789 modi1.n191 modi1.n190 0.019
R11790 modi1.n176 modi1.n171 0.019
R11791 modi1.n2 modi1.n1 0.019
R11792 modi1.n3 modi1.n2 0.019
R11793 modi1.n69 modi1.n68 0.019
R11794 modi1.n78 modi1.n77 0.019
R11795 modi1.n83 modi1.n82 0.019
R11796 modi1.n92 modi1.n89 0.019
R11797 modi1.n149 modi1.n146 0.019
R11798 modi1.n198 modi1.n197 0.018
R11799 modi1.n278 modi1.n277 0.018
R11800 modi1.n293 modi1.n291 0.018
R11801 modi1.n297 modi1.n296 0.018
R11802 modi1.n262 modi1.n260 0.018
R11803 modi1.n139 modi1.n134 0.017
R11804 modi1.n130 modi1.n129 0.017
R11805 modi1.n108 modi1.n107 0.017
R11806 modi1.n101 modi1.n100 0.017
R11807 modi1.n196 modi1.n191 0.017
R11808 modi1.n164 modi1.n163 0.017
R11809 modi1.n176 modi1.n168 0.017
R11810 modi1.n12 modi1.n3 0.017
R11811 modi1.n32 modi1.n27 0.017
R11812 modi1.n83 modi1.n78 0.017
R11813 modi1.n142 modi1.n141 0.016
R11814 modi1.n252 modi1.n251 0.016
R11815 modi1.n246 modi1.n245 0.016
R11816 modi1.n181 modi1.n180 0.016
R11817 modi1.n153 modi1.n152 0.016
R11818 modi1.n71 modi1.n58 0.016
R11819 modi1.n286 modi1.n285 0.016
R11820 modi1.n284 modi1.n283 0.016
R11821 modi1.n268 modi1.n267 0.016
R11822 modi1.n270 modi1.n269 0.016
R11823 modi1.n119 modi1.n114 0.015
R11824 modi1.n216 modi1.n215 0.015
R11825 modi1.n209 modi1.n204 0.015
R11826 modi1.n238 modi1.n237 0.015
R11827 modi1.n232 modi1.n226 0.015
R11828 modi1.n217 modi1.n210 0.015
R11829 modi1.n20 modi1.n16 0.015
R11830 modi1.n57 modi1.n56 0.015
R11831 modi1.n70 modi1.n69 0.015
R11832 modi1.n40 modi1.n35 0.015
R11833 modi1.n58 modi1.n51 0.015
R11834 modi1.n177 modi1.n153 0.014
R11835 modi1.n34 modi1.n33 0.014
R11836 modi1.n50 modi1.n49 0.014
R11837 modi1.n141 modi1.n140 0.013
R11838 modi1.n233 modi1.n232 0.013
R11839 modi1.n226 modi1.n221 0.013
R11840 modi1.n105 modi1.n104 0.012
R11841 modi1.n206 modi1.n205 0.012
R11842 modi1.n129 modi1.n124 0.012
R11843 modi1.n102 modi1.n101 0.012
R11844 modi1.n215 modi1.n214 0.012
R11845 modi1.n163 modi1.n158 0.012
R11846 modi1.n27 modi1.n26 0.012
R11847 modi1.n143 modi1.n142 0.011
R11848 modi1.n251 modi1.n250 0.011
R11849 modi1.n239 modi1.n238 0.011
R11850 modi1.n218 modi1.n217 0.011
R11851 modi1.n182 modi1.n181 0.011
R11852 modi1.n152 modi1.n151 0.011
R11853 modi1.n24 modi1.n23 0.011
R11854 modi1.n287 modi1.n282 0.011
R11855 modi1.n278 modi1.n276 0.011
R11856 modi1.n262 modi1.n261 0.011
R11857 modi1.n272 modi1.n265 0.011
R11858 modi1.n294 modi1.n290 0.011
R11859 modi1.n298 modi1.n295 0.011
R11860 modi1.n210 modi1.n201 0.01
R11861 modi1.n184 modi1.n183 0.01
R11862 modi1.n253 modi1.n252 0.009
R11863 modi1.n241 modi1.n240 0.009
R11864 modi1.n187 modi1.n186 0.009
R11865 modi1.n99 modi1.n98 0.008
R11866 modi1.n223 modi1.n222 0.008
R11867 modi1.n245 modi1.n244 0.008
R11868 modi1.n244 modi1.n243 0.008
R11869 modi1.n37 modi1.n36 0.008
R11870 modi1.n53 modi1.n52 0.008
R11871 modi1.n85 modi1.n84 0.008
R11872 modi1.n285 modi1.n284 0.008
R11873 modi1.n269 modi1.n268 0.008
R11874 modi1.n197 modi1.n187 0.007
R11875 modi1.n41 modi1.n40 0.007
R11876 modi1.n74 modi1.n73 0.007
R11877 modi1.n281 modi1.n280 0.007
R11878 modi1.n299 modi1.n294 0.007
R11879 modi1.n299 modi1.n298 0.007
R11880 modi1.n274 modi1.n264 0.007
R11881 modi1.n131 modi1.n130 0.006
R11882 modi1.n121 modi1.n120 0.006
R11883 modi1.n155 modi1.n154 0.006
R11884 modi1.n165 modi1.n164 0.006
R11885 modi1.n201 modi1.n200 0.006
R11886 modi1.n23 modi1.n22 0.006
R11887 modi1.n144 modi1.n143 0.005
R11888 modi1.n250 modi1.n249 0.005
R11889 modi1.n240 modi1.n239 0.005
R11890 modi1.n183 modi1.n182 0.005
R11891 modi1.n178 modi1.n177 0.005
R11892 modi1 modi1.n301 0.005
R11893 modi1.n89 modi1.n88 0.004
R11894 modi1.n146 modi1.n145 0.004
R11895 modi1.n280 modi1.n279 0.004
R11896 modi1.n264 modi1.n263 0.004
R11897 modi1.n274 modi1.n273 0.004
R11898 modi1.n301 modi1.n300 0.004
R11899 modi1.n275 modi1.n259 0.003
R11900 modi1.n300 modi1.n289 0.002
R11901 modi1.n288 modi1.n281 0.002
R11902 modi1.n235 modi1.n234 0.002
R11903 modi1.n234 modi1.n233 0.002
R11904 modi1.n221 modi1.n220 0.002
R11905 modi1.n35 modi1.n34 0.002
R11906 modi1.n51 modi1.n50 0.002
R11907 modi1.n289 modi1.n275 0.002
R11908 modi1.n247 modi1.n246 0.001
R11909 fout0.n109 fout0.t11 1038.92
R11910 fout0.n519 fout0.t6 1037.29
R11911 fout0.n520 fout0.t12 798.832
R11912 fout0.n125 fout0.t5 795.548
R11913 fout0.n479 fout0.t8 732.329
R11914 fout0.n37 fout0.t3 731.671
R11915 fout0.n12 fout0.t9 731.671
R11916 fout0.n0 fout0.t7 730.671
R11917 fout0.n57 fout0.t4 400.617
R11918 fout0.n86 fout0.t13 400.598
R11919 fout0.n494 fout0.t14 397.317
R11920 fout0.n0 fout0.t10 395.839
R11921 fout0.n319 fout0.n318 13.176
R11922 fout0.n131 fout0.t2 11.723
R11923 fout0.n131 fout0.t1 10.996
R11924 fout0.n139 fout0.n137 9.3
R11925 fout0.n441 fout0.n440 9.3
R11926 fout0.n187 fout0.n186 9.3
R11927 fout0.n189 fout0.n188 9.3
R11928 fout0.n246 fout0.n245 9.3
R11929 fout0.n243 fout0.n242 9.3
R11930 fout0.n201 fout0.n200 9.3
R11931 fout0.n199 fout0.n198 9.3
R11932 fout0.n325 fout0.n324 9.3
R11933 fout0.n224 fout0.n223 9.3
R11934 fout0.n232 fout0.n231 9.3
R11935 fout0.n235 fout0.n234 9.3
R11936 fout0.n355 fout0.n354 9.3
R11937 fout0.n352 fout0.n351 9.3
R11938 fout0.n436 fout0.n435 9.3
R11939 fout0.n434 fout0.n433 9.3
R11940 fout0.n427 fout0.n426 8.097
R11941 fout0.n234 fout0.n233 5.457
R11942 fout0.n354 fout0.n353 5.08
R11943 fout0.n425 fout0.n424 4.65
R11944 fout0.n364 fout0.n363 4.65
R11945 fout0.n446 fout0.n439 4.5
R11946 fout0.n420 fout0.n419 4.5
R11947 fout0.n413 fout0.n412 4.5
R11948 fout0.n344 fout0.n343 4.5
R11949 fout0.n334 fout0.n333 4.5
R11950 fout0.n321 fout0.n320 4.5
R11951 fout0.n297 fout0.n296 4.5
R11952 fout0.n229 fout0.n221 4.5
R11953 fout0.n252 fout0.n251 4.5
R11954 fout0.n197 fout0.n196 4.5
R11955 fout0.n209 fout0.n208 4.5
R11956 fout0.n216 fout0.n215 4.5
R11957 fout0.n260 fout0.n259 4.5
R11958 fout0.n240 fout0.n239 4.5
R11959 fout0.n406 fout0.n405 4.5
R11960 fout0.n185 fout0.n184 4.5
R11961 fout0.n455 fout0.n452 4.5
R11962 fout0.n142 fout0.n141 4.5
R11963 fout0.n208 fout0.n206 4.314
R11964 fout0.n259 fout0.n256 3.944
R11965 fout0.n419 fout0.n418 3.937
R11966 fout0.n405 fout0.n404 3.567
R11967 fout0.n365 fout0.n358 3.033
R11968 fout0.n429 fout0.n428 3.033
R11969 fout0.n426 fout0.t0 2.9
R11970 fout0.n258 fout0.n257 2.258
R11971 fout0.n403 fout0.n402 2.258
R11972 fout0.n214 fout0.n213 1.882
R11973 fout0.n215 fout0.n214 1.882
R11974 fout0.n411 fout0.n410 1.882
R11975 fout0.n467 fout0.n131 1.516
R11976 fout0.n405 fout0.n403 1.505
R11977 fout0.n412 fout0.n411 1.505
R11978 fout0.n447 fout0.n446 1.5
R11979 fout0.n298 fout0.n297 1.5
R11980 fout0.n335 fout0.n334 1.5
R11981 fout0.n366 fout0.n365 1.5
R11982 fout0.n345 fout0.n344 1.5
R11983 fout0.n456 fout0.n455 1.5
R11984 fout0.n143 fout0.n142 1.5
R11985 fout0.n46 fout0.n45 1.435
R11986 fout0.n75 fout0.n74 1.435
R11987 fout0.n533 fout0.n519 1.388
R11988 fout0.n111 fout0.n109 1.355
R11989 fout0.n126 fout0.n125 1.355
R11990 fout0.n521 fout0.n520 1.354
R11991 fout0.n496 fout0.n494 1.354
R11992 fout0.n480 fout0.n479 1.354
R11993 fout0.n38 fout0.n37 1.354
R11994 fout0.n13 fout0.n12 1.354
R11995 fout0.n497 fout0.n496 1.142
R11996 fout0.n112 fout0.n111 1.142
R11997 fout0.n39 fout0.n38 1.142
R11998 fout0.n14 fout0.n13 1.142
R11999 fout0.n498 fout0.n497 1.138
R12000 fout0.n40 fout0.n39 1.138
R12001 fout0.n69 fout0.n14 1.138
R12002 fout0.n113 fout0.n112 1.138
R12003 fout0.n481 fout0.n480 1.137
R12004 fout0.n507 fout0.n506 1.137
R12005 fout0.n472 fout0.n471 1.137
R12006 fout0.n502 fout0.n501 1.137
R12007 fout0.n487 fout0.n486 1.137
R12008 fout0.n23 fout0.n22 1.137
R12009 fout0.n52 fout0.n51 1.137
R12010 fout0.n19 fout0.n18 1.137
R12011 fout0.n29 fout0.n28 1.137
R12012 fout0.n47 fout0.n46 1.137
R12013 fout0.n66 fout0.n65 1.137
R12014 fout0.n81 fout0.n80 1.137
R12015 fout0.n62 fout0.n61 1.137
R12016 fout0.n4 fout0.n3 1.137
R12017 fout0.n76 fout0.n75 1.137
R12018 fout0.n127 fout0.n126 1.137
R12019 fout0.n95 fout0.n94 1.137
R12020 fout0.n118 fout0.n117 1.137
R12021 fout0.n92 fout0.n91 1.137
R12022 fout0.n102 fout0.n101 1.137
R12023 fout0.n509 fout0.n508 1.136
R12024 fout0.n97 fout0.n96 1.136
R12025 fout0.n483 fout0.n482 1.136
R12026 fout0.n129 fout0.n128 1.136
R12027 fout0.n84 fout0.n83 1.136
R12028 fout0.n68 fout0.n67 1.136
R12029 fout0.n55 fout0.n54 1.136
R12030 fout0.n25 fout0.n24 1.136
R12031 fout0.n184 fout0.n183 1.129
R12032 fout0.n259 fout0.n258 1.129
R12033 fout0.n251 fout0.n250 1.129
R12034 fout0.n261 fout0.n260 1.042
R12035 fout0.n278 fout0.n277 0.853
R12036 fout0.n368 fout0.n367 0.853
R12037 fout0.n462 fout0.n461 0.853
R12038 fout0.n155 fout0.n154 0.853
R12039 fout0.n541 fout0.n540 0.827
R12040 fout0.n141 fout0.n140 0.752
R12041 fout0.n333 fout0.n332 0.752
R12042 fout0.n343 fout0.n342 0.752
R12043 fout0.n419 fout0.n417 0.752
R12044 fout0.n439 fout0.n438 0.752
R12045 fout0.n452 fout0.n451 0.752
R12046 fout0.n145 fout0.n144 0.717
R12047 fout0.n467 fout0.n466 0.69
R12048 fout0.n468 fout0.n467 0.68
R12049 fout0.n324 fout0.n323 0.536
R12050 fout0.n223 fout0.n222 0.536
R12051 fout0.n245 fout0.n244 0.475
R12052 fout0.n363 fout0.n362 0.475
R12053 fout0.n541 fout0.n510 0.471
R12054 fout0.n534 fout0.n533 0.44
R12055 fout0.n428 fout0.n427 0.382
R12056 fout0.n195 fout0.n194 0.382
R12057 fout0.n196 fout0.n195 0.376
R12058 fout0.n208 fout0.n207 0.376
R12059 fout0.n239 fout0.n238 0.376
R12060 fout0.n221 fout0.n220 0.376
R12061 fout0.n296 fout0.n295 0.376
R12062 fout0.n320 fout0.n319 0.376
R12063 fout0.n183 fout0.n182 0.349
R12064 fout0.n438 fout0.n437 0.349
R12065 fout0 fout0.n541 0.229
R12066 fout0.n88 fout0.n87 0.152
R12067 fout0.n57 fout0.n56 0.123
R12068 fout0.n86 fout0.n85 0.123
R12069 fout0.n58 fout0.n57 0.091
R12070 fout0.n494 fout0.n493 0.083
R12071 fout0.n479 fout0.n478 0.083
R12072 fout0.n37 fout0.n36 0.083
R12073 fout0.n12 fout0.n11 0.083
R12074 fout0.n519 fout0.n518 0.076
R12075 fout0 fout0.n130 0.076
R12076 fout0.n109 fout0.n108 0.075
R12077 fout0.n125 fout0.n124 0.075
R12078 fout0.n87 fout0.n86 0.07
R12079 fout0.n515 fout0.n514 0.059
R12080 fout0.n236 fout0.n235 0.047
R12081 fout0.n226 fout0.n225 0.047
R12082 fout0.n315 fout0.n314 0.047
R12083 fout0.n328 fout0.n327 0.047
R12084 fout0.n356 fout0.n355 0.047
R12085 fout0.n443 fout0.n442 0.047
R12086 fout0.n422 fout0.n421 0.043
R12087 fout0.n391 fout0.n390 0.043
R12088 fout0.n205 fout0.n204 0.041
R12089 fout0.n172 fout0.n171 0.041
R12090 fout0.n431 fout0.n430 0.035
R12091 fout0.n299 fout0.n298 0.035
R12092 fout0.n304 fout0.n303 0.035
R12093 fout0.n397 fout0.n396 0.035
R12094 fout0.n192 fout0.n191 0.034
R12095 fout0.n313 fout0.n312 0.034
R12096 fout0.n317 fout0.n316 0.034
R12097 fout0.n434 fout0.n432 0.034
R12098 fout0.n152 fout0.n151 0.034
R12099 fout0.n150 fout0.n149 0.034
R12100 fout0.n268 fout0.n267 0.034
R12101 fout0.n275 fout0.n274 0.034
R12102 fout0.n335 fout0.n311 0.034
R12103 fout0.n337 fout0.n336 0.034
R12104 fout0.n350 fout0.n349 0.034
R12105 fout0.n399 fout0.n398 0.034
R12106 fout0.n529 fout0.n528 0.032
R12107 fout0.n528 fout0.n527 0.032
R12108 fout0.n506 fout0.n504 0.032
R12109 fout0.n190 fout0.n189 0.032
R12110 fout0.n365 fout0.n364 0.032
R12111 fout0.n429 fout0.n425 0.032
R12112 fout0.n273 fout0.n272 0.032
R12113 fout0.n447 fout0.n399 0.032
R12114 fout0.n18 fout0.n17 0.032
R12115 fout0.n61 fout0.n60 0.032
R12116 fout0.n91 fout0.n90 0.032
R12117 fout0.n533 fout0.n532 0.032
R12118 fout0.n157 fout0.n156 0.031
R12119 fout0.n168 fout0.n167 0.031
R12120 fout0.n280 fout0.n279 0.031
R12121 fout0.n291 fout0.n290 0.031
R12122 fout0.n370 fout0.n369 0.031
R12123 fout0.n381 fout0.n380 0.031
R12124 fout0.n464 fout0.n463 0.031
R12125 fout0.n523 fout0.n522 0.03
R12126 fout0.n199 fout0.n197 0.03
R12127 fout0.n243 fout0.n241 0.03
R12128 fout0.n228 fout0.n227 0.03
R12129 fout0.n330 fout0.n329 0.03
R12130 fout0.n444 fout0.n443 0.03
R12131 fout0.n153 fout0.n152 0.03
R12132 fout0.n147 fout0.n146 0.03
R12133 fout0.n271 fout0.n270 0.03
R12134 fout0.n309 fout0.n308 0.03
R12135 fout0.n338 fout0.n337 0.03
R12136 fout0.n394 fout0.n393 0.03
R12137 fout0.n461 fout0.n460 0.03
R12138 fout0.n532 fout0.n531 0.028
R12139 fout0.n530 fout0.n529 0.028
R12140 fout0.n527 fout0.n526 0.028
R12141 fout0.n525 fout0.n524 0.028
R12142 fout0.n493 fout0.n492 0.028
R12143 fout0.n491 fout0.n490 0.028
R12144 fout0.n476 fout0.n475 0.028
R12145 fout0.n478 fout0.n477 0.028
R12146 fout0.n486 fout0.n485 0.028
R12147 fout0.n501 fout0.n500 0.028
R12148 fout0.n506 fout0.n505 0.028
R12149 fout0.n471 fout0.n469 0.028
R12150 fout0.n142 fout0.n139 0.028
R12151 fout0.n180 fout0.n179 0.028
R12152 fout0.n203 fout0.n202 0.028
R12153 fout0.n218 fout0.n217 0.028
R12154 fout0.n260 fout0.n219 0.028
R12155 fout0.n249 fout0.n248 0.028
R12156 fout0.n365 fout0.n357 0.028
R12157 fout0.n409 fout0.n408 0.028
R12158 fout0.n423 fout0.n422 0.028
R12159 fout0.n446 fout0.n436 0.028
R12160 fout0.n143 fout0.n135 0.028
R12161 fout0.n170 fout0.n169 0.028
R12162 fout0.n177 fout0.n176 0.028
R12163 fout0.n261 fout0.n178 0.028
R12164 fout0.n266 fout0.n265 0.028
R12165 fout0.n276 fout0.n275 0.028
R12166 fout0.n293 fout0.n292 0.028
R12167 fout0.n306 fout0.n305 0.028
R12168 fout0.n367 fout0.n366 0.028
R12169 fout0.n386 fout0.n385 0.028
R12170 fout0.n392 fout0.n391 0.028
R12171 fout0.n457 fout0.n456 0.028
R12172 fout0.n45 fout0.n44 0.028
R12173 fout0.n43 fout0.n42 0.028
R12174 fout0.n34 fout0.n33 0.028
R12175 fout0.n36 fout0.n35 0.028
R12176 fout0.n51 fout0.n50 0.028
R12177 fout0.n18 fout0.n16 0.028
R12178 fout0.n22 fout0.n21 0.028
R12179 fout0.n28 fout0.n26 0.028
R12180 fout0.n74 fout0.n73 0.028
R12181 fout0.n72 fout0.n71 0.028
R12182 fout0.n9 fout0.n8 0.028
R12183 fout0.n11 fout0.n10 0.028
R12184 fout0.n80 fout0.n79 0.028
R12185 fout0.n61 fout0.n59 0.028
R12186 fout0.n65 fout0.n64 0.028
R12187 fout0.n3 fout0.n1 0.028
R12188 fout0.n101 fout0.n100 0.028
R12189 fout0.n91 fout0.n89 0.028
R12190 fout0.n94 fout0.n93 0.028
R12191 fout0.n117 fout0.n115 0.028
R12192 fout0.n161 fout0.n160 0.027
R12193 fout0.n164 fout0.n163 0.027
R12194 fout0.n284 fout0.n283 0.027
R12195 fout0.n287 fout0.n286 0.027
R12196 fout0.n374 fout0.n373 0.027
R12197 fout0.n377 fout0.n376 0.027
R12198 fout0.n518 fout0.n517 0.026
R12199 fout0.n516 fout0.n515 0.026
R12200 fout0.n514 fout0.n513 0.026
R12201 fout0.n512 fout0.n511 0.026
R12202 fout0.n187 fout0.n185 0.026
R12203 fout0.n240 fout0.n237 0.026
R12204 fout0.n360 fout0.n359 0.026
R12205 fout0.n407 fout0.n406 0.026
R12206 fout0.n263 fout0.n262 0.026
R12207 fout0.n277 fout0.n269 0.026
R12208 fout0.n348 fout0.n347 0.026
R12209 fout0.n384 fout0.n383 0.026
R12210 fout0.n389 fout0.n388 0.026
R12211 fout0.n459 fout0.n458 0.026
R12212 fout0.n108 fout0.n107 0.025
R12213 fout0.n106 fout0.n105 0.025
R12214 fout0.n122 fout0.n121 0.025
R12215 fout0.n124 fout0.n123 0.025
R12216 fout0.n144 fout0.n143 0.024
R12217 fout0.n247 fout0.n246 0.024
R12218 fout0.n364 fout0.n361 0.024
R12219 fout0.n134 fout0.n133 0.024
R12220 fout0.n174 fout0.n173 0.024
R12221 fout0.n269 fout0.n268 0.024
R12222 fout0.n302 fout0.n301 0.024
R12223 fout0.n345 fout0.n339 0.024
R12224 fout0.n537 fout0.n536 0.023
R12225 fout0.n211 fout0.n210 0.022
R12226 fout0.n237 fout0.n236 0.022
R12227 fout0.n325 fout0.n322 0.022
R12228 fout0.n361 fout0.n360 0.022
R12229 fout0.n416 fout0.n415 0.022
R12230 fout0.n133 fout0.n132 0.022
R12231 fout0.n277 fout0.n276 0.022
R12232 fout0.n301 fout0.n300 0.022
R12233 fout0.n366 fout0.n350 0.022
R12234 fout0.n349 fout0.n348 0.022
R12235 fout0.n254 fout0.n253 0.02
R12236 fout0.n252 fout0.n249 0.02
R12237 fout0.n248 fout0.n247 0.02
R12238 fout0.n357 fout0.n356 0.02
R12239 fout0.n341 fout0.n340 0.02
R12240 fout0.n154 fout0.n153 0.02
R12241 fout0.n267 fout0.n266 0.02
R12242 fout0.n367 fout0.n338 0.02
R12243 fout0.n460 fout0.n459 0.02
R12244 fout0.n456 fout0.n450 0.02
R12245 fout0.n155 fout0.n145 0.019
R12246 fout0.n156 fout0.n155 0.019
R12247 fout0.n278 fout0.n168 0.019
R12248 fout0.n279 fout0.n278 0.019
R12249 fout0.n368 fout0.n291 0.019
R12250 fout0.n369 fout0.n368 0.019
R12251 fout0.n462 fout0.n381 0.019
R12252 fout0.n463 fout0.n462 0.019
R12253 fout0.n425 fout0.n423 0.018
R12254 fout0.n175 fout0.n174 0.018
R12255 fout0.n461 fout0.n447 0.018
R12256 fout0.n524 fout0.n523 0.017
R12257 fout0.n522 fout0.n521 0.017
R12258 fout0.n496 fout0.n495 0.017
R12259 fout0.n486 fout0.n484 0.017
R12260 fout0.n471 fout0.n470 0.017
R12261 fout0.n480 fout0.n474 0.017
R12262 fout0.n202 fout0.n201 0.017
R12263 fout0.n230 fout0.n229 0.017
R12264 fout0.n227 fout0.n226 0.017
R12265 fout0.n454 fout0.n453 0.017
R12266 fout0.n262 fout0.n261 0.017
R12267 fout0.n265 fout0.n264 0.017
R12268 fout0.n274 fout0.n273 0.017
R12269 fout0.n272 fout0.n271 0.017
R12270 fout0.n347 fout0.n346 0.017
R12271 fout0.n388 fout0.n387 0.017
R12272 fout0.n393 fout0.n392 0.017
R12273 fout0.n450 fout0.n449 0.017
R12274 fout0.n46 fout0.n41 0.017
R12275 fout0.n51 fout0.n49 0.017
R12276 fout0.n28 fout0.n27 0.017
R12277 fout0.n38 fout0.n32 0.017
R12278 fout0.n75 fout0.n70 0.017
R12279 fout0.n80 fout0.n78 0.017
R12280 fout0.n3 fout0.n2 0.017
R12281 fout0.n13 fout0.n7 0.017
R12282 fout0.n111 fout0.n110 0.017
R12283 fout0.n101 fout0.n99 0.017
R12284 fout0.n117 fout0.n116 0.017
R12285 fout0.n126 fout0.n120 0.017
R12286 fout0.n502 fout0.n499 0.016
R12287 fout0.n507 fout0.n503 0.016
R12288 fout0.n23 fout0.n20 0.016
R12289 fout0.n66 fout0.n63 0.016
R12290 fout0.n531 fout0.n530 0.015
R12291 fout0.n526 fout0.n525 0.015
R12292 fout0.n492 fout0.n491 0.015
R12293 fout0.n477 fout0.n476 0.015
R12294 fout0.n181 fout0.n180 0.015
R12295 fout0.n191 fout0.n190 0.015
R12296 fout0.n219 fout0.n218 0.015
R12297 fout0.n329 fout0.n328 0.015
R12298 fout0.n334 fout0.n331 0.015
R12299 fout0.n408 fout0.n407 0.015
R12300 fout0.n413 fout0.n409 0.015
R12301 fout0.n445 fout0.n444 0.015
R12302 fout0.n151 fout0.n150 0.015
R12303 fout0.n149 fout0.n148 0.015
R12304 fout0.n178 fout0.n177 0.015
R12305 fout0.n308 fout0.n307 0.015
R12306 fout0.n311 fout0.n310 0.015
R12307 fout0.n336 fout0.n335 0.015
R12308 fout0.n385 fout0.n384 0.015
R12309 fout0.n387 fout0.n386 0.015
R12310 fout0.n44 fout0.n43 0.015
R12311 fout0.n35 fout0.n34 0.015
R12312 fout0.n73 fout0.n72 0.015
R12313 fout0.n10 fout0.n9 0.015
R12314 fout0.n517 fout0.n516 0.013
R12315 fout0.n513 fout0.n512 0.013
R12316 fout0.n193 fout0.n192 0.013
R12317 fout0.n217 fout0.n216 0.013
R12318 fout0.n232 fout0.n230 0.013
R12319 fout0.n430 fout0.n429 0.013
R12320 fout0.n432 fout0.n431 0.013
R12321 fout0.n176 fout0.n175 0.013
R12322 fout0.n396 fout0.n395 0.013
R12323 fout0.n398 fout0.n397 0.013
R12324 fout0.n466 fout0.n465 0.013
R12325 fout0.n107 fout0.n106 0.013
R12326 fout0.n123 fout0.n122 0.013
R12327 fout0.n508 fout0.n502 0.012
R12328 fout0.n508 fout0.n507 0.012
R12329 fout0.n162 fout0.n161 0.012
R12330 fout0.n163 fout0.n162 0.012
R12331 fout0.n285 fout0.n284 0.012
R12332 fout0.n286 fout0.n285 0.012
R12333 fout0.n375 fout0.n374 0.012
R12334 fout0.n376 fout0.n375 0.012
R12335 fout0.n24 fout0.n19 0.012
R12336 fout0.n24 fout0.n23 0.012
R12337 fout0.n67 fout0.n62 0.012
R12338 fout0.n67 fout0.n66 0.012
R12339 fout0.n96 fout0.n92 0.012
R12340 fout0.n96 fout0.n95 0.012
R12341 fout0.n489 fout0.n488 0.011
R12342 fout0.n482 fout0.n473 0.011
R12343 fout0.n255 fout0.n254 0.011
R12344 fout0.n159 fout0.n158 0.011
R12345 fout0.n166 fout0.n165 0.011
R12346 fout0.n282 fout0.n281 0.011
R12347 fout0.n289 fout0.n288 0.011
R12348 fout0.n372 fout0.n371 0.011
R12349 fout0.n379 fout0.n378 0.011
R12350 fout0.n54 fout0.n53 0.011
R12351 fout0.n31 fout0.n30 0.011
R12352 fout0.n83 fout0.n82 0.011
R12353 fout0.n6 fout0.n5 0.011
R12354 fout0.n104 fout0.n103 0.011
R12355 fout0.n128 fout0.n119 0.011
R12356 fout0.n52 fout0.n48 0.01
R12357 fout0.n81 fout0.n77 0.01
R12358 fout0.n102 fout0.n98 0.01
R12359 fout0.n118 fout0.n114 0.01
R12360 fout0.n535 fout0.n534 0.01
R12361 fout0.n536 fout0.n535 0.01
R12362 fout0.n539 fout0.n538 0.009
R12363 fout0.n139 fout0.n138 0.009
R12364 fout0.n212 fout0.n211 0.009
R12365 fout0.n216 fout0.n212 0.009
R12366 fout0.n314 fout0.n313 0.009
R12367 fout0.n415 fout0.n414 0.009
R12368 fout0.n135 fout0.n134 0.009
R12369 fout0.n300 fout0.n299 0.009
R12370 fout0.n209 fout0.n205 0.007
R12371 fout0.n297 fout0.n294 0.007
R12372 fout0.n316 fout0.n315 0.007
R12373 fout0.n322 fout0.n321 0.007
R12374 fout0.n414 fout0.n413 0.007
R12375 fout0.n442 fout0.n441 0.007
R12376 fout0.n173 fout0.n172 0.007
R12377 fout0.n298 fout0.n293 0.007
R12378 fout0.n303 fout0.n302 0.007
R12379 fout0.n305 fout0.n304 0.007
R12380 fout0.n458 fout0.n457 0.007
R12381 fout0.n449 fout0.n448 0.007
R12382 fout0.n488 fout0.n487 0.006
R12383 fout0.n473 fout0.n472 0.006
R12384 fout0.n482 fout0.n481 0.006
R12385 fout0.n158 fout0.n157 0.006
R12386 fout0.n160 fout0.n159 0.006
R12387 fout0.n165 fout0.n164 0.006
R12388 fout0.n167 fout0.n166 0.006
R12389 fout0.n281 fout0.n280 0.006
R12390 fout0.n283 fout0.n282 0.006
R12391 fout0.n288 fout0.n287 0.006
R12392 fout0.n290 fout0.n289 0.006
R12393 fout0.n371 fout0.n370 0.006
R12394 fout0.n373 fout0.n372 0.006
R12395 fout0.n378 fout0.n377 0.006
R12396 fout0.n380 fout0.n379 0.006
R12397 fout0.n465 fout0.n464 0.006
R12398 fout0.n54 fout0.n47 0.006
R12399 fout0.n53 fout0.n52 0.006
R12400 fout0.n30 fout0.n29 0.006
R12401 fout0.n83 fout0.n76 0.006
R12402 fout0.n82 fout0.n81 0.006
R12403 fout0.n5 fout0.n4 0.006
R12404 fout0.n103 fout0.n102 0.006
R12405 fout0.n119 fout0.n118 0.006
R12406 fout0.n128 fout0.n127 0.006
R12407 fout0.n538 fout0.n537 0.005
R12408 fout0.n540 fout0.n539 0.005
R12409 fout0.n185 fout0.n181 0.005
R12410 fout0.n189 fout0.n187 0.005
R12411 fout0.n260 fout0.n255 0.005
R12412 fout0.n253 fout0.n252 0.005
R12413 fout0.n225 fout0.n224 0.005
R12414 fout0.n326 fout0.n325 0.005
R12415 fout0.n401 fout0.n400 0.005
R12416 fout0.n421 fout0.n420 0.005
R12417 fout0.n346 fout0.n345 0.005
R12418 fout0.n390 fout0.n389 0.005
R12419 fout0.n510 fout0.n509 0.004
R12420 fout0.n97 fout0.n88 0.004
R12421 fout0.n483 fout0.n468 0.003
R12422 fout0.n25 fout0.n15 0.003
R12423 fout0.n56 fout0.n55 0.003
R12424 fout0.n68 fout0.n58 0.003
R12425 fout0.n85 fout0.n84 0.003
R12426 fout0.n130 fout0.n129 0.003
R12427 fout0.n142 fout0.n136 0.003
R12428 fout0.n334 fout0.n330 0.003
R12429 fout0.n355 fout0.n352 0.003
R12430 fout0.n344 fout0.n341 0.003
R12431 fout0.n420 fout0.n416 0.003
R12432 fout0.n436 fout0.n434 0.003
R12433 fout0.n446 fout0.n445 0.003
R12434 fout0.n455 fout0.n454 0.003
R12435 fout0.n264 fout0.n263 0.003
R12436 fout0.n395 fout0.n394 0.003
R12437 fout0.n497 fout0.n489 0.003
R12438 fout0.n112 fout0.n104 0.003
R12439 fout0.n14 fout0.n6 0.003
R12440 fout0.n39 fout0.n31 0.003
R12441 fout0.n509 fout0.n498 0.002
R12442 fout0.n113 fout0.n97 0.002
R12443 fout0.n498 fout0.n483 0.002
R12444 fout0.n129 fout0.n113 0.002
R12445 fout0.n84 fout0.n69 0.002
R12446 fout0.n55 fout0.n40 0.002
R12447 fout0.n69 fout0.n68 0.002
R12448 fout0.n40 fout0.n25 0.002
R12449 fout0.n197 fout0.n193 0.001
R12450 fout0.n201 fout0.n199 0.001
R12451 fout0.n204 fout0.n203 0.001
R12452 fout0.n210 fout0.n209 0.001
R12453 fout0.n246 fout0.n243 0.001
R12454 fout0.n241 fout0.n240 0.001
R12455 fout0.n235 fout0.n232 0.001
R12456 fout0.n229 fout0.n228 0.001
R12457 fout0.n321 fout0.n317 0.001
R12458 fout0.n327 fout0.n326 0.001
R12459 fout0.n406 fout0.n401 0.001
R12460 fout0.n148 fout0.n147 0.001
R12461 fout0.n171 fout0.n170 0.001
R12462 fout0.n307 fout0.n306 0.001
R12463 fout0.n310 fout0.n309 0.001
R12464 fout0.n383 fout0.n382 0.001
R12465 fout0.n87 fout0.n0 0.001
R12466 modi0.n267 modi0.t5 1037.92
R12467 modi0.n258 modi0.t3 1037.28
R12468 modi0.n267 modi0.t2 798.492
R12469 modi0.n258 modi0.t4 797.528
R12470 modi0.n31 modi0.n30 92.5
R12471 modi0.n59 modi0.n58 92.5
R12472 modi0.n58 modi0.t0 70.344
R12473 modi0.n19 modi0.n18 31.034
R12474 modi0.n50 modi0.n49 31.034
R12475 modi0.n114 modi0.n113 9.3
R12476 modi0.n191 modi0.n190 9.3
R12477 modi0.n3 modi0.n2 9.3
R12478 modi0.n51 modi0.n50 9.3
R12479 modi0.n20 modi0.n19 9.3
R12480 modi0.n78 modi0.n77 9.3
R12481 modi0.n230 modi0.n229 9.154
R12482 modi0.n32 modi0.n31 8.282
R12483 modi0.n60 modi0.n59 8.282
R12484 modi0.n229 modi0.t1 7.141
R12485 modi0.n150 modi0.n149 7.033
R12486 modi0.n93 modi0.n92 7.033
R12487 modi0.n259 modi0.n257 6.416
R12488 modi0.n20 modi0.n16 5.647
R12489 modi0.n51 modi0.n47 5.647
R12490 modi0.n231 modi0.n230 4.65
R12491 modi0.n57 modi0.n56 4.65
R12492 modi0.n177 modi0.n176 4.5
R12493 modi0.n197 modi0.n196 4.5
R12494 modi0.n210 modi0.n209 4.5
R12495 modi0.n217 modi0.n214 4.5
R12496 modi0.n226 modi0.n225 4.5
R12497 modi0.n232 modi0.n228 4.5
R12498 modi0.n101 modi0.n98 4.5
R12499 modi0.n108 modi0.n107 4.5
R12500 modi0.n120 modi0.n119 4.5
R12501 modi0.n130 modi0.n129 4.5
R12502 modi0.n140 modi0.n139 4.5
R12503 modi0.n164 modi0.n163 4.5
R12504 modi0.n84 modi0.n82 4.5
R12505 modi0.n55 modi0.n52 4.5
R12506 modi0.n70 modi0.n68 4.5
R12507 modi0.n33 modi0.n32 4.5
R12508 modi0.n40 modi0.n39 4.5
R12509 modi0.n61 modi0.n60 4.5
R12510 modi0.n23 modi0.n22 4.5
R12511 modi0.n8 modi0.n7 4.5
R12512 modi0.n129 modi0.n126 4.141
R12513 modi0.n163 modi0.n162 4.141
R12514 modi0.n18 modi0.n17 4.137
R12515 modi0.n49 modi0.n48 4.137
R12516 modi0 modi0.n259 3.871
R12517 modi0.n119 modi0.n116 3.764
R12518 modi0.n209 modi0.n207 3.764
R12519 modi0.n7 modi0.n5 3.764
R12520 modi0.n52 modi0.n45 3.764
R12521 modi0.n272 modi0.n267 3.461
R12522 modi0.n139 modi0.n136 3.388
R12523 modi0.n107 modi0.n106 3.388
R12524 modi0.n196 modi0.n195 3.388
R12525 modi0.n176 modi0.n175 3.388
R12526 modi0.n22 modi0.n21 3.388
R12527 modi0.n82 modi0.n81 3.388
R12528 modi0.n139 modi0.n138 3.011
R12529 modi0.n107 modi0.n104 3.011
R12530 modi0.n98 modi0.n96 3.011
R12531 modi0.n190 modi0.n189 3.011
R12532 modi0.n196 modi0.n194 3.011
R12533 modi0.n176 modi0.n174 3.011
R12534 modi0.n22 modi0.n20 3.011
R12535 modi0.n32 modi0.n29 3.011
R12536 modi0.n82 modi0.n80 3.011
R12537 modi0.n119 modi0.n118 2.635
R12538 modi0.n113 modi0.n112 2.635
R12539 modi0.n214 modi0.n213 2.635
R12540 modi0.n209 modi0.n208 2.635
R12541 modi0.n7 modi0.n6 2.635
R12542 modi0.n68 modi0.n67 2.635
R12543 modi0.n52 modi0.n51 2.635
R12544 modi0.n129 modi0.n128 2.258
R12545 modi0.n163 modi0.n161 2.258
R12546 modi0.n259 modi0.n258 2.25
R12547 modi0.n26 modi0.n0 1.754
R12548 modi0.n180 modi0.n151 1.754
R12549 modi0.n26 modi0.n25 1.705
R12550 modi0.n43 modi0.n42 1.705
R12551 modi0.n73 modi0.n72 1.705
R12552 modi0.n87 modi0.n86 1.705
R12553 modi0.n256 modi0.n145 1.705
R12554 modi0.n200 modi0.n199 1.705
R12555 modi0.n220 modi0.n219 1.705
R12556 modi0.n249 modi0.n248 1.705
R12557 modi0.n255 modi0.n254 1.705
R12558 modi0.n243 modi0.n242 1.705
R12559 modi0.n237 modi0.n236 1.705
R12560 modi0.n186 modi0.n185 1.705
R12561 modi0.n180 modi0.n179 1.705
R12562 modi0.n214 modi0.n212 1.505
R12563 modi0.n198 modi0.n197 1.5
R12564 modi0.n211 modi0.n210 1.5
R12565 modi0.n218 modi0.n217 1.5
R12566 modi0.n227 modi0.n226 1.5
R12567 modi0.n233 modi0.n232 1.5
R12568 modi0.n85 modi0.n84 1.5
R12569 modi0.n72 modi0.n55 1.5
R12570 modi0.n34 modi0.n33 1.5
R12571 modi0.n71 modi0.n70 1.5
R12572 modi0.n41 modi0.n40 1.5
R12573 modi0.n62 modi0.n61 1.5
R12574 modi0.n24 modi0.n23 1.5
R12575 modi0.n9 modi0.n8 1.5
R12576 modi0.n288 modi0.n287 1.402
R12577 modi0.n273 modi0.n272 1.355
R12578 modi0.n257 modi0.n256 1.267
R12579 modi0.n289 modi0.n288 1.141
R12580 modi0.n290 modi0.n289 1.137
R12581 modi0.n280 modi0.n279 1.137
R12582 modi0.n295 modi0.n294 1.137
R12583 modi0.n274 modi0.n273 1.137
R12584 modi0.n264 modi0.n263 1.137
R12585 modi0.n299 modi0.n298 1.137
R12586 modi0.n301 modi0.n300 1.136
R12587 modi0.n276 modi0.n275 1.136
R12588 modi0.n98 modi0.n97 1.129
R12589 modi0.n151 modi0.n150 1.127
R12590 modi0.n145 modi0.n93 1.127
R12591 modi0.n141 modi0.n140 1.125
R12592 modi0.n178 modi0.n177 1.125
R12593 modi0.n16 modi0.n15 0.752
R12594 modi0.n47 modi0.n46 0.752
R12595 modi0.n257 modi0.n87 0.71
R12596 modi0.n92 modi0.n91 0.155
R12597 modi0.n149 modi0.n148 0.155
R12598 modi0.n138 modi0.n137 0.144
R12599 modi0.n174 modi0.n173 0.144
R12600 modi0.n128 modi0.n127 0.133
R12601 modi0.n161 modi0.n160 0.132
R12602 modi0.n134 modi0.n133 0.053
R12603 modi0.n124 modi0.n123 0.053
R12604 modi0.n114 modi0.n111 0.053
R12605 modi0.n158 modi0.n157 0.053
R12606 modi0.n168 modi0.n167 0.053
R12607 modi0.n171 modi0.n170 0.053
R12608 modi0.n78 modi0.n76 0.053
R12609 modi0.n43 modi0.n26 0.049
R12610 modi0.n73 modi0.n43 0.049
R12611 modi0.n87 modi0.n73 0.049
R12612 modi0.n256 modi0.n255 0.049
R12613 modi0.n255 modi0.n249 0.049
R12614 modi0.n249 modi0.n243 0.049
R12615 modi0.n243 modi0.n237 0.049
R12616 modi0.n237 modi0.n220 0.049
R12617 modi0.n220 modi0.n200 0.049
R12618 modi0.n200 modi0.n186 0.049
R12619 modi0.n186 modi0.n180 0.049
R12620 modi0.n272 modi0.n271 0.048
R12621 modi0.n40 modi0.n38 0.045
R12622 modi0.n70 modi0.n66 0.045
R12623 modi0.n101 modi0.n100 0.043
R12624 modi0.n226 modi0.n224 0.043
R12625 modi0.n89 modi0.n88 0.034
R12626 modi0.n167 modi0.n166 0.032
R12627 modi0.n135 modi0.n134 0.03
R12628 modi0.n133 modi0.n132 0.03
R12629 modi0.n157 modi0.n156 0.03
R12630 modi0.n10 modi0.n9 0.03
R12631 modi0.n85 modi0.n75 0.03
R12632 modi0.n123 modi0.n122 0.028
R12633 modi0.n169 modi0.n168 0.028
R12634 modi0.n172 modi0.n171 0.028
R12635 modi0.n95 modi0.n94 0.025
R12636 modi0.n125 modi0.n124 0.025
R12637 modi0.n61 modi0.n57 0.025
R12638 modi0.n118 modi0.n117 0.024
R12639 modi0.n194 modi0.n193 0.024
R12640 modi0.n232 modi0.n231 0.023
R12641 modi0.n159 modi0.n158 0.023
R12642 modi0.n121 modi0.n120 0.021
R12643 modi0.n115 modi0.n114 0.021
R12644 modi0.n204 modi0.n203 0.021
R12645 modi0.n8 modi0.n1 0.021
R12646 modi0.n4 modi0.n3 0.021
R12647 modi0.n55 modi0.n44 0.021
R12648 modi0.n294 modi0.n293 0.021
R12649 modi0.n140 modi0.n95 0.019
R12650 modi0.n111 modi0.n110 0.019
R12651 modi0.n110 modi0.n109 0.019
R12652 modi0.n108 modi0.n103 0.019
R12653 modi0.n205 modi0.n204 0.019
R12654 modi0.n192 modi0.n191 0.019
R12655 modi0.n177 modi0.n172 0.019
R12656 modi0.n199 modi0.n198 0.019
R12657 modi0.n13 modi0.n12 0.019
R12658 modi0.n14 modi0.n13 0.019
R12659 modi0.n54 modi0.n53 0.019
R12660 modi0.n79 modi0.n78 0.019
R12661 modi0.n84 modi0.n83 0.019
R12662 modi0.n93 modi0.n90 0.019
R12663 modi0.n150 modi0.n147 0.019
R12664 modi0.n279 modi0.n278 0.018
R12665 modi0.n294 modi0.n292 0.018
R12666 modi0.n298 modi0.n297 0.018
R12667 modi0.n263 modi0.n261 0.018
R12668 modi0.n140 modi0.n135 0.017
R12669 modi0.n131 modi0.n130 0.017
R12670 modi0.n109 modi0.n108 0.017
R12671 modi0.n102 modi0.n101 0.017
R12672 modi0.n197 modi0.n192 0.017
R12673 modi0.n165 modi0.n164 0.017
R12674 modi0.n177 modi0.n169 0.017
R12675 modi0.n23 modi0.n14 0.017
R12676 modi0.n33 modi0.n28 0.017
R12677 modi0.n84 modi0.n79 0.017
R12678 modi0.n143 modi0.n142 0.016
R12679 modi0.n253 modi0.n252 0.016
R12680 modi0.n247 modi0.n246 0.016
R12681 modi0.n182 modi0.n181 0.016
R12682 modi0.n154 modi0.n153 0.016
R12683 modi0.n287 modi0.n286 0.016
R12684 modi0.n285 modi0.n284 0.016
R12685 modi0.n269 modi0.n268 0.016
R12686 modi0.n271 modi0.n270 0.016
R12687 modi0.n120 modi0.n115 0.015
R12688 modi0.n217 modi0.n216 0.015
R12689 modi0.n210 modi0.n205 0.015
R12690 modi0.n239 modi0.n238 0.015
R12691 modi0.n233 modi0.n227 0.015
R12692 modi0.n218 modi0.n211 0.015
R12693 modi0.n8 modi0.n4 0.015
R12694 modi0.n70 modi0.n69 0.015
R12695 modi0.n55 modi0.n54 0.015
R12696 modi0.n41 modi0.n36 0.015
R12697 modi0.n71 modi0.n64 0.015
R12698 modi0.n72 modi0.n71 0.015
R12699 modi0.n178 modi0.n154 0.014
R12700 modi0.n35 modi0.n34 0.014
R12701 modi0.n63 modi0.n62 0.014
R12702 modi0.n142 modi0.n141 0.013
R12703 modi0.n234 modi0.n233 0.013
R12704 modi0.n227 modi0.n222 0.013
R12705 modi0.n106 modi0.n105 0.012
R12706 modi0.n207 modi0.n206 0.012
R12707 modi0.n130 modi0.n125 0.012
R12708 modi0.n103 modi0.n102 0.012
R12709 modi0.n216 modi0.n215 0.012
R12710 modi0.n164 modi0.n159 0.012
R12711 modi0.n28 modi0.n27 0.012
R12712 modi0.n144 modi0.n143 0.011
R12713 modi0.n252 modi0.n251 0.011
R12714 modi0.n240 modi0.n239 0.011
R12715 modi0.n219 modi0.n218 0.011
R12716 modi0.n185 modi0.n184 0.011
R12717 modi0.n183 modi0.n182 0.011
R12718 modi0.n153 modi0.n152 0.011
R12719 modi0.n288 modi0.n283 0.011
R12720 modi0.n279 modi0.n277 0.011
R12721 modi0.n263 modi0.n262 0.011
R12722 modi0.n273 modi0.n266 0.011
R12723 modi0.n295 modi0.n291 0.011
R12724 modi0.n299 modi0.n296 0.011
R12725 modi0.n242 modi0.n241 0.01
R12726 modi0.n211 modi0.n202 0.01
R12727 modi0.n25 modi0.n11 0.01
R12728 modi0.n254 modi0.n253 0.009
R12729 modi0.n188 modi0.n187 0.009
R12730 modi0.n100 modi0.n99 0.008
R12731 modi0.n224 modi0.n223 0.008
R12732 modi0.n246 modi0.n245 0.008
R12733 modi0.n245 modi0.n244 0.008
R12734 modi0.n38 modi0.n37 0.008
R12735 modi0.n66 modi0.n65 0.008
R12736 modi0.n286 modi0.n285 0.008
R12737 modi0.n270 modi0.n269 0.008
R12738 modi0.n198 modi0.n188 0.007
R12739 modi0.n42 modi0.n41 0.007
R12740 modi0.n75 modi0.n74 0.007
R12741 modi0.n86 modi0.n85 0.007
R12742 modi0.n282 modi0.n281 0.007
R12743 modi0.n300 modi0.n295 0.007
R12744 modi0.n300 modi0.n299 0.007
R12745 modi0.n275 modi0.n265 0.007
R12746 modi0.n132 modi0.n131 0.006
R12747 modi0.n122 modi0.n121 0.006
R12748 modi0.n156 modi0.n155 0.006
R12749 modi0.n166 modi0.n165 0.006
R12750 modi0.n202 modi0.n201 0.006
R12751 modi0.n11 modi0.n10 0.006
R12752 modi0.n145 modi0.n144 0.005
R12753 modi0.n251 modi0.n250 0.005
R12754 modi0.n241 modi0.n240 0.005
R12755 modi0.n184 modi0.n183 0.005
R12756 modi0.n179 modi0.n178 0.005
R12757 modi0 modi0.n302 0.005
R12758 modi0.n90 modi0.n89 0.004
R12759 modi0.n147 modi0.n146 0.004
R12760 modi0.n281 modi0.n280 0.004
R12761 modi0.n265 modi0.n264 0.004
R12762 modi0.n275 modi0.n274 0.004
R12763 modi0.n302 modi0.n301 0.004
R12764 modi0.n276 modi0.n260 0.003
R12765 modi0.n236 modi0.n235 0.003
R12766 modi0.n301 modi0.n290 0.002
R12767 modi0.n289 modi0.n282 0.002
R12768 modi0.n235 modi0.n234 0.002
R12769 modi0.n222 modi0.n221 0.002
R12770 modi0.n36 modi0.n35 0.002
R12771 modi0.n64 modi0.n63 0.002
R12772 modi0.n290 modi0.n276 0.002
R12773 modi0.n248 modi0.n247 0.001
R12774 modi0.n25 modi0.n24 0.001
R12775 modi4.n6 modi4.t2 1037.92
R12776 modi4.n43 modi4.t4 1037.28
R12777 modi4.n43 modi4.t3 797.53
R12778 modi4.n6 modi4.t5 796.885
R12779 modi4.n291 modi4.n290 92.5
R12780 modi4.n263 modi4.n262 92.5
R12781 modi4.n290 modi4.t0 70.344
R12782 modi4.n277 modi4.n276 31.034
R12783 modi4.n243 modi4.n242 31.034
R12784 modi4.n218 modi4.n217 9.3
R12785 modi4.n278 modi4.n277 9.3
R12786 modi4.n244 modi4.n243 9.3
R12787 modi4.n228 modi4.n227 9.3
R12788 modi4.n90 modi4.n89 9.3
R12789 modi4.n172 modi4.n171 9.3
R12790 modi4.n128 modi4.n127 9.154
R12791 modi4.n292 modi4.n291 8.282
R12792 modi4.n264 modi4.n263 8.282
R12793 modi4.n127 modi4.t1 7.141
R12794 modi4.n48 modi4.n47 7.033
R12795 modi4.n210 modi4.n209 7.032
R12796 modi4.n301 modi4.n300 6.465
R12797 modi4.n278 modi4.n274 5.647
R12798 modi4.n244 modi4.n240 5.647
R12799 modi4.n284 modi4.n283 4.65
R12800 modi4.n129 modi4.n128 4.65
R12801 modi4.n234 modi4.n232 4.5
R12802 modi4.n249 modi4.n245 4.5
R12803 modi4.n256 modi4.n253 4.5
R12804 modi4.n281 modi4.n280 4.5
R12805 modi4.n295 modi4.n292 4.5
R12806 modi4.n285 modi4.n282 4.5
R12807 modi4.n265 modi4.n264 4.5
R12808 modi4.n223 modi4.n222 4.5
R12809 modi4.n200 modi4.n199 4.5
R12810 modi4.n188 modi4.n187 4.5
R12811 modi4.n178 modi4.n177 4.5
R12812 modi4.n166 modi4.n165 4.5
R12813 modi4.n159 modi4.n158 4.5
R12814 modi4.n131 modi4.n130 4.5
R12815 modi4.n125 modi4.n124 4.5
R12816 modi4.n116 modi4.n115 4.5
R12817 modi4.n109 modi4.n108 4.5
R12818 modi4.n96 modi4.n95 4.5
R12819 modi4.n65 modi4.n64 4.5
R12820 modi4.n75 modi4.n74 4.5
R12821 modi4.n64 modi4.n61 4.141
R12822 modi4.n187 modi4.n186 4.141
R12823 modi4.n276 modi4.n275 4.137
R12824 modi4.n242 modi4.n241 4.137
R12825 modi4.n222 modi4.n220 3.764
R12826 modi4.n245 modi4.n238 3.764
R12827 modi4.n95 modi4.n92 3.764
R12828 modi4.n165 modi4.n163 3.764
R12829 modi4.n11 modi4.n6 3.464
R12830 modi4.n280 modi4.n279 3.388
R12831 modi4.n232 modi4.n231 3.388
R12832 modi4.n74 modi4.n71 3.388
R12833 modi4.n108 modi4.n107 3.388
R12834 modi4.n177 modi4.n176 3.388
R12835 modi4.n199 modi4.n198 3.388
R12836 modi4 modi4.n301 3.014
R12837 modi4.n280 modi4.n278 3.011
R12838 modi4.n292 modi4.n289 3.011
R12839 modi4.n232 modi4.n230 3.011
R12840 modi4.n74 modi4.n73 3.011
R12841 modi4.n108 modi4.n105 3.011
R12842 modi4.n115 modi4.n113 3.011
R12843 modi4.n171 modi4.n170 3.011
R12844 modi4.n177 modi4.n175 3.011
R12845 modi4.n199 modi4.n197 3.011
R12846 modi4.n222 modi4.n221 2.635
R12847 modi4.n253 modi4.n252 2.635
R12848 modi4.n245 modi4.n244 2.635
R12849 modi4.n95 modi4.n94 2.635
R12850 modi4.n89 modi4.n88 2.635
R12851 modi4.n158 modi4.n157 2.635
R12852 modi4.n165 modi4.n164 2.635
R12853 modi4.n64 modi4.n63 2.258
R12854 modi4.n187 modi4.n185 2.258
R12855 modi4.n301 modi4.n43 2.25
R12856 modi4.n78 modi4.n49 1.754
R12857 modi4.n251 modi4.n226 1.754
R12858 modi4.n78 modi4.n77 1.705
R12859 modi4.n153 modi4.n152 1.705
R12860 modi4.n147 modi4.n146 1.705
R12861 modi4.n142 modi4.n141 1.705
R12862 modi4.n136 modi4.n135 1.705
R12863 modi4.n119 modi4.n118 1.705
R12864 modi4.n99 modi4.n98 1.705
R12865 modi4.n84 modi4.n83 1.705
R12866 modi4.n299 modi4.n225 1.705
R12867 modi4.n298 modi4.n297 1.705
R12868 modi4.n268 modi4.n267 1.705
R12869 modi4.n251 modi4.n250 1.705
R12870 modi4.n212 modi4.n211 1.705
R12871 modi4.n158 modi4.n156 1.505
R12872 modi4.n235 modi4.n234 1.5
R12873 modi4.n250 modi4.n249 1.5
R12874 modi4.n297 modi4.n281 1.5
R12875 modi4.n296 modi4.n295 1.5
R12876 modi4.n257 modi4.n256 1.5
R12877 modi4.n286 modi4.n285 1.5
R12878 modi4.n266 modi4.n265 1.5
R12879 modi4.n224 modi4.n223 1.5
R12880 modi4.n132 modi4.n131 1.5
R12881 modi4.n126 modi4.n125 1.5
R12882 modi4.n117 modi4.n116 1.5
R12883 modi4.n110 modi4.n109 1.5
R12884 modi4.n97 modi4.n96 1.5
R12885 modi4.n38 modi4.n37 1.402
R12886 modi4.n13 modi4.n11 1.355
R12887 modi4.n300 modi4.n212 1.268
R12888 modi4.n14 modi4.n13 1.141
R12889 modi4.n26 modi4.n14 1.137
R12890 modi4.n3 modi4.n2 1.137
R12891 modi4.n20 modi4.n19 1.137
R12892 modi4.n39 modi4.n38 1.137
R12893 modi4.n31 modi4.n30 1.137
R12894 modi4.n23 modi4.n22 1.137
R12895 modi4.n25 modi4.n24 1.136
R12896 modi4.n41 modi4.n40 1.136
R12897 modi4.n211 modi4.n210 1.129
R12898 modi4.n115 modi4.n114 1.129
R12899 modi4.n49 modi4.n48 1.127
R12900 modi4.n201 modi4.n200 1.125
R12901 modi4.n76 modi4.n75 1.125
R12902 modi4.n274 modi4.n273 0.752
R12903 modi4.n240 modi4.n239 0.752
R12904 modi4.n300 modi4.n299 0.709
R12905 modi4.n47 modi4.n46 0.155
R12906 modi4.n209 modi4.n208 0.155
R12907 modi4.n73 modi4.n72 0.144
R12908 modi4.n197 modi4.n196 0.144
R12909 modi4.n63 modi4.n62 0.133
R12910 modi4.n185 modi4.n184 0.132
R12911 modi4.n218 modi4.n216 0.053
R12912 modi4.n54 modi4.n53 0.053
R12913 modi4.n69 modi4.n68 0.053
R12914 modi4.n59 modi4.n58 0.053
R12915 modi4.n172 modi4.n169 0.053
R12916 modi4.n182 modi4.n181 0.053
R12917 modi4.n192 modi4.n191 0.053
R12918 modi4.n84 modi4.n78 0.049
R12919 modi4.n99 modi4.n84 0.049
R12920 modi4.n119 modi4.n99 0.049
R12921 modi4.n136 modi4.n119 0.049
R12922 modi4.n142 modi4.n136 0.049
R12923 modi4.n147 modi4.n142 0.049
R12924 modi4.n153 modi4.n147 0.049
R12925 modi4.n212 modi4.n153 0.049
R12926 modi4.n299 modi4.n298 0.049
R12927 modi4.n298 modi4.n268 0.049
R12928 modi4.n268 modi4.n251 0.049
R12929 modi4.n11 modi4.n10 0.048
R12930 modi4.n125 modi4.n123 0.045
R12931 modi4.n159 modi4.n155 0.045
R12932 modi4.n295 modi4.n294 0.043
R12933 modi4.n265 modi4.n261 0.043
R12934 modi4.n191 modi4.n190 0.032
R12935 modi4.n206 modi4.n205 0.032
R12936 modi4.n224 modi4.n214 0.03
R12937 modi4.n236 modi4.n235 0.03
R12938 modi4.n70 modi4.n69 0.03
R12939 modi4.n68 modi4.n67 0.03
R12940 modi4.n181 modi4.n180 0.03
R12941 modi4.n58 modi4.n57 0.028
R12942 modi4.n193 modi4.n192 0.028
R12943 modi4.n195 modi4.n194 0.028
R12944 modi4.n55 modi4.n54 0.025
R12945 modi4.n60 modi4.n59 0.025
R12946 modi4.n131 modi4.n129 0.025
R12947 modi4.n94 modi4.n93 0.024
R12948 modi4.n175 modi4.n174 0.024
R12949 modi4.n285 modi4.n284 0.023
R12950 modi4.n183 modi4.n182 0.023
R12951 modi4.n223 modi4.n215 0.021
R12952 modi4.n219 modi4.n218 0.021
R12953 modi4.n247 modi4.n246 0.021
R12954 modi4.n91 modi4.n90 0.021
R12955 modi4.n166 modi4.n161 0.021
R12956 modi4.n169 modi4.n168 0.021
R12957 modi4.n19 modi4.n18 0.021
R12958 modi4.n270 modi4.n269 0.019
R12959 modi4.n281 modi4.n272 0.019
R12960 modi4.n248 modi4.n247 0.019
R12961 modi4.n229 modi4.n228 0.019
R12962 modi4.n234 modi4.n233 0.019
R12963 modi4.n75 modi4.n55 0.019
R12964 modi4.n103 modi4.n102 0.019
R12965 modi4.n104 modi4.n103 0.019
R12966 modi4.n168 modi4.n167 0.019
R12967 modi4.n173 modi4.n172 0.019
R12968 modi4.n179 modi4.n178 0.019
R12969 modi4.n200 modi4.n195 0.019
R12970 modi4.n210 modi4.n207 0.019
R12971 modi4.n48 modi4.n45 0.019
R12972 modi4.n2 modi4.n1 0.018
R12973 modi4.n19 modi4.n17 0.018
R12974 modi4.n22 modi4.n21 0.018
R12975 modi4.n30 modi4.n28 0.018
R12976 modi4.n281 modi4.n270 0.017
R12977 modi4.n234 modi4.n229 0.017
R12978 modi4.n75 modi4.n70 0.017
R12979 modi4.n66 modi4.n65 0.017
R12980 modi4.n109 modi4.n104 0.017
R12981 modi4.n116 modi4.n112 0.017
R12982 modi4.n178 modi4.n173 0.017
R12983 modi4.n189 modi4.n188 0.017
R12984 modi4.n200 modi4.n193 0.017
R12985 modi4.n98 modi4.n97 0.017
R12986 modi4.n297 modi4.n296 0.016
R12987 modi4.n52 modi4.n51 0.016
R12988 modi4.n80 modi4.n79 0.016
R12989 modi4.n86 modi4.n85 0.016
R12990 modi4.n146 modi4.n145 0.016
R12991 modi4.n151 modi4.n150 0.016
R12992 modi4.n203 modi4.n202 0.016
R12993 modi4.n10 modi4.n9 0.016
R12994 modi4.n8 modi4.n7 0.016
R12995 modi4.n35 modi4.n34 0.016
R12996 modi4.n37 modi4.n36 0.016
R12997 modi4 modi4.n42 0.016
R12998 modi4.n223 modi4.n219 0.015
R12999 modi4.n256 modi4.n255 0.015
R13000 modi4.n249 modi4.n248 0.015
R13001 modi4.n287 modi4.n286 0.015
R13002 modi4.n258 modi4.n257 0.015
R13003 modi4.n96 modi4.n91 0.015
R13004 modi4.n160 modi4.n159 0.015
R13005 modi4.n167 modi4.n166 0.015
R13006 modi4.n117 modi4.n110 0.015
R13007 modi4.n132 modi4.n126 0.015
R13008 modi4.n138 modi4.n137 0.015
R13009 modi4.n296 modi4.n288 0.014
R13010 modi4.n266 modi4.n259 0.014
R13011 modi4.n202 modi4.n201 0.014
R13012 modi4.n76 modi4.n52 0.013
R13013 modi4.n126 modi4.n121 0.013
R13014 modi4.n133 modi4.n132 0.013
R13015 modi4.n107 modi4.n106 0.012
R13016 modi4.n163 modi4.n162 0.012
R13017 modi4.n272 modi4.n271 0.012
R13018 modi4.n255 modi4.n254 0.012
R13019 modi4.n65 modi4.n60 0.012
R13020 modi4.n112 modi4.n111 0.012
R13021 modi4.n161 modi4.n160 0.012
R13022 modi4.n188 modi4.n183 0.012
R13023 modi4.n250 modi4.n237 0.011
R13024 modi4.n51 modi4.n50 0.011
R13025 modi4.n81 modi4.n80 0.011
R13026 modi4.n110 modi4.n101 0.011
R13027 modi4.n150 modi4.n149 0.011
R13028 modi4.n204 modi4.n203 0.011
R13029 modi4.n13 modi4.n12 0.011
R13030 modi4.n2 modi4.n0 0.011
R13031 modi4.n30 modi4.n29 0.011
R13032 modi4.n38 modi4.n33 0.011
R13033 modi4.n20 modi4.n16 0.011
R13034 modi4.n83 modi4.n82 0.01
R13035 modi4.n118 modi4.n117 0.01
R13036 modi4.n139 modi4.n138 0.01
R13037 modi4.n225 modi4.n224 0.009
R13038 modi4.n141 modi4.n140 0.009
R13039 modi4.n145 modi4.n144 0.009
R13040 modi4.n294 modi4.n293 0.008
R13041 modi4.n261 modi4.n260 0.008
R13042 modi4.n267 modi4.n266 0.008
R13043 modi4.n123 modi4.n122 0.008
R13044 modi4.n155 modi4.n154 0.008
R13045 modi4.n87 modi4.n86 0.008
R13046 modi4.n97 modi4.n87 0.008
R13047 modi4.n152 modi4.n151 0.008
R13048 modi4.n9 modi4.n8 0.008
R13049 modi4.n36 modi4.n35 0.008
R13050 modi4.n237 modi4.n236 0.007
R13051 modi4.n144 modi4.n143 0.007
R13052 modi4.n5 modi4.n4 0.007
R13053 modi4.n24 modi4.n20 0.007
R13054 modi4.n24 modi4.n23 0.007
R13055 modi4.n40 modi4.n32 0.007
R13056 modi4.n31 modi4.n27 0.007
R13057 modi4.n214 modi4.n213 0.006
R13058 modi4.n67 modi4.n66 0.006
R13059 modi4.n57 modi4.n56 0.006
R13060 modi4.n180 modi4.n179 0.006
R13061 modi4.n190 modi4.n189 0.006
R13062 modi4.n140 modi4.n139 0.006
R13063 modi4.n77 modi4.n76 0.005
R13064 modi4.n82 modi4.n81 0.005
R13065 modi4.n101 modi4.n100 0.005
R13066 modi4.n149 modi4.n148 0.005
R13067 modi4.n211 modi4.n204 0.005
R13068 modi4.n45 modi4.n44 0.004
R13069 modi4.n207 modi4.n206 0.004
R13070 modi4.n4 modi4.n3 0.004
R13071 modi4.n32 modi4.n31 0.004
R13072 modi4.n40 modi4.n39 0.004
R13073 modi4.n25 modi4.n15 0.004
R13074 modi4.n42 modi4.n41 0.003
R13075 modi4.n26 modi4.n25 0.002
R13076 modi4.n14 modi4.n5 0.002
R13077 modi4.n288 modi4.n287 0.002
R13078 modi4.n259 modi4.n258 0.002
R13079 modi4.n121 modi4.n120 0.002
R13080 modi4.n134 modi4.n133 0.002
R13081 modi4.n135 modi4.n134 0.002
R13082 modi4.n41 modi4.n26 0.002
R13083 a_n7001_2908.n95 a_n7001_2908.t4 730.681
R13084 a_n7001_2908.n95 a_n7001_2908.t3 395.834
R13085 a_n7001_2908.n41 a_n7001_2908.n40 13.176
R13086 a_n7001_2908.n96 a_n7001_2908.t2 11.72
R13087 a_n7001_2908.n96 a_n7001_2908.t0 10.994
R13088 a_n7001_2908.n150 a_n7001_2908.n34 9.3
R13089 a_n7001_2908.n150 a_n7001_2908.n141 9.3
R13090 a_n7001_2908.n150 a_n7001_2908.n135 9.3
R13091 a_n7001_2908.n150 a_n7001_2908.n49 9.3
R13092 a_n7001_2908.n150 a_n7001_2908.n54 9.3
R13093 a_n7001_2908.n150 a_n7001_2908.n123 9.3
R13094 a_n7001_2908.n150 a_n7001_2908.n149 8.469
R13095 a_n7001_2908.n150 a_n7001_2908.n113 8.469
R13096 a_n7001_2908.n150 a_n7001_2908.n118 8.125
R13097 a_n7001_2908.n150 a_n7001_2908.n29 8.124
R13098 a_n7001_2908.n150 a_n7001_2908.n110 8.097
R13099 a_n7001_2908.n150 a_n7001_2908.n146 8.096
R13100 a_n7001_2908.n150 a_n7001_2908.n126 8.016
R13101 a_n7001_2908.n150 a_n7001_2908.n39 8.016
R13102 a_n7001_2908.n150 a_n7001_2908.n130 7.964
R13103 a_n7001_2908.n150 a_n7001_2908.n44 7.964
R13104 a_n7001_2908.n125 a_n7001_2908.n124 6.4
R13105 a_n7001_2908.n109 a_n7001_2908.n55 6.4
R13106 a_n7001_2908.n144 a_n7001_2908.n143 6.023
R13107 a_n7001_2908.n37 a_n7001_2908.n36 6.023
R13108 a_n7001_2908.n135 a_n7001_2908.n134 6.023
R13109 a_n7001_2908.n43 a_n7001_2908.n42 6.023
R13110 a_n7001_2908.n129 a_n7001_2908.n128 6.023
R13111 a_n7001_2908.n148 a_n7001_2908.n147 5.647
R13112 a_n7001_2908.n49 a_n7001_2908.n46 5.647
R13113 a_n7001_2908.n116 a_n7001_2908.n115 5.647
R13114 a_n7001_2908.n112 a_n7001_2908.n111 5.647
R13115 a_n7001_2908.n132 a_n7001_2908.n131 5.457
R13116 a_n7001_2908.n27 a_n7001_2908.n26 5.27
R13117 a_n7001_2908.n48 a_n7001_2908.n47 5.08
R13118 a_n7001_2908.n34 a_n7001_2908.n33 4.517
R13119 a_n7001_2908.n123 a_n7001_2908.n120 4.517
R13120 a_n7001_2908.n63 a_n7001_2908.n62 4.5
R13121 a_n7001_2908.n2 a_n7001_2908.n1 4.5
R13122 a_n7001_2908.n31 a_n7001_2908.n30 4.314
R13123 a_n7001_2908.n140 a_n7001_2908.n139 4.141
R13124 a_n7001_2908.n51 a_n7001_2908.n50 4.141
R13125 a_n7001_2908.n137 a_n7001_2908.n136 3.944
R13126 a_n7001_2908.n122 a_n7001_2908.n121 3.937
R13127 a_n7001_2908.n53 a_n7001_2908.n52 3.567
R13128 a_n7001_2908.n109 a_n7001_2908.n108 3.033
R13129 a_n7001_2908.t1 a_n7001_2908.n150 2.9
R13130 a_n7001_2908.n141 a_n7001_2908.n140 2.258
R13131 a_n7001_2908.n54 a_n7001_2908.n51 2.258
R13132 a_n7001_2908.n33 a_n7001_2908.n32 1.882
R13133 a_n7001_2908.n120 a_n7001_2908.n119 1.882
R13134 a_n7001_2908.n98 a_n7001_2908.n97 1.672
R13135 a_n7001_2908.n54 a_n7001_2908.n53 1.505
R13136 a_n7001_2908.n82 a_n7001_2908.n102 1.5
R13137 a_n7001_2908.n64 a_n7001_2908.n66 1.5
R13138 a_n7001_2908.n63 a_n7001_2908.n61 1.5
R13139 a_n7001_2908.n21 a_n7001_2908.n24 1.5
R13140 a_n7001_2908.n12 a_n7001_2908.n11 1.5
R13141 a_n7001_2908.n108 a_n7001_2908.n80 1.5
R13142 a_n7001_2908.n97 a_n7001_2908.n96 1.222
R13143 a_n7001_2908.n28 a_n7001_2908.n27 1.129
R13144 a_n7001_2908.n26 a_n7001_2908.n25 1.129
R13145 a_n7001_2908.n141 a_n7001_2908.n137 1.129
R13146 a_n7001_2908.n139 a_n7001_2908.n138 1.129
R13147 a_n7001_2908.n101 a_n7001_2908.n100 0.853
R13148 a_n7001_2908.n149 a_n7001_2908.n148 0.752
R13149 a_n7001_2908.n46 a_n7001_2908.n45 0.752
R13150 a_n7001_2908.n49 a_n7001_2908.n48 0.752
R13151 a_n7001_2908.n123 a_n7001_2908.n122 0.752
R13152 a_n7001_2908.n115 a_n7001_2908.n114 0.752
R13153 a_n7001_2908.n117 a_n7001_2908.n116 0.752
R13154 a_n7001_2908.n113 a_n7001_2908.n112 0.752
R13155 a_n7001_2908.n89 a_n7001_2908.n88 0.716
R13156 a_n7001_2908.n97 a_n7001_2908.n95 0.637
R13157 a_n7001_2908.n130 a_n7001_2908.n129 0.536
R13158 a_n7001_2908.n44 a_n7001_2908.n43 0.536
R13159 a_n7001_2908.n126 a_n7001_2908.n125 0.476
R13160 a_n7001_2908.n39 a_n7001_2908.n38 0.475
R13161 a_n7001_2908.n110 a_n7001_2908.n109 0.382
R13162 a_n7001_2908.n146 a_n7001_2908.n145 0.382
R13163 a_n7001_2908.n145 a_n7001_2908.n144 0.376
R13164 a_n7001_2908.n143 a_n7001_2908.n142 0.376
R13165 a_n7001_2908.n34 a_n7001_2908.n31 0.376
R13166 a_n7001_2908.n38 a_n7001_2908.n37 0.376
R13167 a_n7001_2908.n36 a_n7001_2908.n35 0.376
R13168 a_n7001_2908.n135 a_n7001_2908.n132 0.376
R13169 a_n7001_2908.n134 a_n7001_2908.n133 0.376
R13170 a_n7001_2908.n42 a_n7001_2908.n41 0.376
R13171 a_n7001_2908.n128 a_n7001_2908.n127 0.376
R13172 a_n7001_2908.n118 a_n7001_2908.n117 0.35
R13173 a_n7001_2908.n29 a_n7001_2908.n28 0.349
R13174 a_n7001_2908.n2 a_n7001_2908.n0 0.066
R13175 a_n7001_2908.n87 a_n7001_2908.n86 0.047
R13176 a_n7001_2908.n72 a_n7001_2908.n71 0.043
R13177 a_n7001_2908.n68 a_n7001_2908.n67 0.043
R13178 a_n7001_2908.n64 a_n7001_2908.n63 0.041
R13179 a_n7001_2908.n79 a_n7001_2908.n78 0.035
R13180 a_n7001_2908.n107 a_n7001_2908.n106 0.035
R13181 a_n7001_2908.n19 a_n7001_2908.n18 0.034
R13182 a_n7001_2908.n23 a_n7001_2908.n22 0.034
R13183 a_n7001_2908.n8 a_n7001_2908.n7 0.034
R13184 a_n7001_2908.n77 a_n7001_2908.n76 0.034
R13185 a_n7001_2908.n105 a_n7001_2908.n104 0.034
R13186 a_n7001_2908.n12 a_n7001_2908.n6 0.032
R13187 a_n7001_2908.n108 a_n7001_2908.n70 0.032
R13188 a_n7001_2908.n99 a_n7001_2908.n98 0.031
R13189 a_n7001_2908.n9 a_n7001_2908.n8 0.03
R13190 a_n7001_2908.n75 a_n7001_2908.n74 0.03
R13191 a_n7001_2908.n101 a_n7001_2908.n94 0.03
R13192 a_n7001_2908.n81 a_n7001_2908.n87 0.03
R13193 a_n7001_2908.n11 a_n7001_2908.n10 0.028
R13194 a_n7001_2908.n60 a_n7001_2908.n58 0.028
R13195 a_n7001_2908.n73 a_n7001_2908.n72 0.028
R13196 a_n7001_2908.n91 a_n7001_2908.n90 0.028
R13197 a_n7001_2908.n13 a_n7001_2908.n12 0.028
R13198 a_n7001_2908.n57 a_n7001_2908.n56 0.028
R13199 a_n7001_2908.n69 a_n7001_2908.n68 0.028
R13200 a_n7001_2908.n103 a_n7001_2908.n82 0.028
R13201 a_n7001_2908.n85 a_n7001_2908.n83 0.028
R13202 a_n7001_2908.n17 a_n7001_2908.n15 0.026
R13203 a_n7001_2908.n66 a_n7001_2908.n65 0.026
R13204 a_n7001_2908.n93 a_n7001_2908.n92 0.026
R13205 a_n7001_2908.n4 a_n7001_2908.n3 0.026
R13206 a_n7001_2908.n90 a_n7001_2908.n89 0.024
R13207 a_n7001_2908.n18 a_n7001_2908.n17 0.024
R13208 a_n7001_2908.n6 a_n7001_2908.n5 0.024
R13209 a_n7001_2908.n15 a_n7001_2908.n16 0.022
R13210 a_n7001_2908.n5 a_n7001_2908.n4 0.022
R13211 a_n7001_2908.n3 a_n7001_2908.n2 0.022
R13212 a_n7001_2908.n20 a_n7001_2908.n19 0.02
R13213 a_n7001_2908.n10 a_n7001_2908.n9 0.02
R13214 a_n7001_2908.n94 a_n7001_2908.n93 0.02
R13215 a_n7001_2908.n14 a_n7001_2908.n13 0.02
R13216 a_n7001_2908.n100 a_n7001_2908.n99 0.019
R13217 a_n7001_2908.n82 a_n7001_2908.n81 0.018
R13218 a_n7001_2908.n102 a_n7001_2908.n101 0.018
R13219 a_n7001_2908.n70 a_n7001_2908.n69 0.018
R13220 a_n7001_2908.n24 a_n7001_2908.n23 0.017
R13221 a_n7001_2908.n74 a_n7001_2908.n73 0.017
R13222 a_n7001_2908.n58 a_n7001_2908.n59 0.015
R13223 a_n7001_2908.n61 a_n7001_2908.n60 0.015
R13224 a_n7001_2908.n56 a_n7001_2908.n0 0.015
R13225 a_n7001_2908.n63 a_n7001_2908.n57 0.015
R13226 a_n7001_2908.n80 a_n7001_2908.n79 0.013
R13227 a_n7001_2908.n78 a_n7001_2908.n77 0.013
R13228 a_n7001_2908.n108 a_n7001_2908.n107 0.013
R13229 a_n7001_2908.n106 a_n7001_2908.n105 0.013
R13230 a_n7001_2908.n92 a_n7001_2908.n91 0.007
R13231 a_n7001_2908.n86 a_n7001_2908.n85 0.007
R13232 a_n7001_2908.n21 a_n7001_2908.n20 1.424
R13233 a_n7001_2908.n67 a_n7001_2908.n64 0.005
R13234 a_n7001_2908.n80 a_n7001_2908.n75 0.003
R13235 a_n7001_2908.n104 a_n7001_2908.n103 0.003
R13236 a_n7001_2908.n83 a_n7001_2908.n84 0.003
R13237 a_n7001_2908.n14 a_n7001_2908.n21 0.47
R13238 a_n2702_11550.n97 a_n2702_11550.t4 730.68
R13239 a_n2702_11550.n97 a_n2702_11550.t3 395.833
R13240 a_n2702_11550.n46 a_n2702_11550.n45 13.176
R13241 a_n2702_11550.n98 a_n2702_11550.t0 11.724
R13242 a_n2702_11550.n98 a_n2702_11550.t2 10.994
R13243 a_n2702_11550.n137 a_n2702_11550.n39 9.3
R13244 a_n2702_11550.n137 a_n2702_11550.n133 9.3
R13245 a_n2702_11550.n137 a_n2702_11550.n127 9.3
R13246 a_n2702_11550.n137 a_n2702_11550.n58 9.3
R13247 a_n2702_11550.n137 a_n2702_11550.n66 9.3
R13248 a_n2702_11550.n137 a_n2702_11550.n122 9.3
R13249 a_n2702_11550.n137 a_n2702_11550.n117 8.47
R13250 a_n2702_11550.n137 a_n2702_11550.n136 8.469
R13251 a_n2702_11550.n137 a_n2702_11550.n114 8.124
R13252 a_n2702_11550.n137 a_n2702_11550.n29 8.124
R13253 a_n2702_11550.n137 a_n2702_11550.n34 8.097
R13254 a_n2702_11550.n137 a_n2702_11550.n109 8.097
R13255 a_n2702_11550.n137 a_n2702_11550.n61 8.016
R13256 a_n2702_11550.n137 a_n2702_11550.n44 8.016
R13257 a_n2702_11550.n137 a_n2702_11550.n53 7.964
R13258 a_n2702_11550.n137 a_n2702_11550.n49 7.964
R13259 a_n2702_11550.n60 a_n2702_11550.n59 6.4
R13260 a_n2702_11550.n108 a_n2702_11550.n67 6.4
R13261 a_n2702_11550.n32 a_n2702_11550.n31 6.023
R13262 a_n2702_11550.n42 a_n2702_11550.n41 6.023
R13263 a_n2702_11550.n127 a_n2702_11550.n126 6.023
R13264 a_n2702_11550.n48 a_n2702_11550.n47 6.023
R13265 a_n2702_11550.n52 a_n2702_11550.n51 6.023
R13266 a_n2702_11550.n135 a_n2702_11550.n134 5.647
R13267 a_n2702_11550.n58 a_n2702_11550.n55 5.647
R13268 a_n2702_11550.n112 a_n2702_11550.n111 5.647
R13269 a_n2702_11550.n116 a_n2702_11550.n115 5.647
R13270 a_n2702_11550.n124 a_n2702_11550.n123 5.457
R13271 a_n2702_11550.n27 a_n2702_11550.n26 5.27
R13272 a_n2702_11550.n57 a_n2702_11550.n56 5.08
R13273 a_n2702_11550.n39 a_n2702_11550.n38 4.517
R13274 a_n2702_11550.n122 a_n2702_11550.n119 4.517
R13275 a_n2702_11550.n75 a_n2702_11550.n74 4.5
R13276 a_n2702_11550.n2 a_n2702_11550.n1 4.5
R13277 a_n2702_11550.n36 a_n2702_11550.n35 4.314
R13278 a_n2702_11550.n132 a_n2702_11550.n131 4.141
R13279 a_n2702_11550.n63 a_n2702_11550.n62 4.141
R13280 a_n2702_11550.n129 a_n2702_11550.n128 3.944
R13281 a_n2702_11550.n121 a_n2702_11550.n120 3.937
R13282 a_n2702_11550.n65 a_n2702_11550.n64 3.567
R13283 a_n2702_11550.n108 a_n2702_11550.n107 3.033
R13284 a_n2702_11550.t1 a_n2702_11550.n137 2.9
R13285 a_n2702_11550.n133 a_n2702_11550.n132 2.258
R13286 a_n2702_11550.n66 a_n2702_11550.n63 2.258
R13287 a_n2702_11550.n100 a_n2702_11550.n99 1.903
R13288 a_n2702_11550.n38 a_n2702_11550.n37 1.882
R13289 a_n2702_11550.n119 a_n2702_11550.n118 1.882
R13290 a_n2702_11550.n66 a_n2702_11550.n65 1.505
R13291 a_n2702_11550.n94 a_n2702_11550.n101 1.5
R13292 a_n2702_11550.n76 a_n2702_11550.n78 1.5
R13293 a_n2702_11550.n75 a_n2702_11550.n73 1.5
R13294 a_n2702_11550.n21 a_n2702_11550.n24 1.5
R13295 a_n2702_11550.n12 a_n2702_11550.n11 1.5
R13296 a_n2702_11550.n107 a_n2702_11550.n92 1.5
R13297 a_n2702_11550.n99 a_n2702_11550.n98 1.223
R13298 a_n2702_11550.n28 a_n2702_11550.n27 1.129
R13299 a_n2702_11550.n26 a_n2702_11550.n25 1.129
R13300 a_n2702_11550.n133 a_n2702_11550.n129 1.129
R13301 a_n2702_11550.n131 a_n2702_11550.n130 1.129
R13302 a_n2702_11550.n136 a_n2702_11550.n135 0.752
R13303 a_n2702_11550.n55 a_n2702_11550.n54 0.752
R13304 a_n2702_11550.n58 a_n2702_11550.n57 0.752
R13305 a_n2702_11550.n122 a_n2702_11550.n121 0.752
R13306 a_n2702_11550.n111 a_n2702_11550.n110 0.752
R13307 a_n2702_11550.n113 a_n2702_11550.n112 0.752
R13308 a_n2702_11550.n117 a_n2702_11550.n116 0.752
R13309 a_n2702_11550.n99 a_n2702_11550.n97 0.637
R13310 a_n2702_11550.n53 a_n2702_11550.n52 0.536
R13311 a_n2702_11550.n49 a_n2702_11550.n48 0.536
R13312 a_n2702_11550.n61 a_n2702_11550.n60 0.475
R13313 a_n2702_11550.n44 a_n2702_11550.n43 0.475
R13314 a_n2702_11550.n34 a_n2702_11550.n33 0.382
R13315 a_n2702_11550.n109 a_n2702_11550.n108 0.382
R13316 a_n2702_11550.n33 a_n2702_11550.n32 0.376
R13317 a_n2702_11550.n31 a_n2702_11550.n30 0.376
R13318 a_n2702_11550.n39 a_n2702_11550.n36 0.376
R13319 a_n2702_11550.n43 a_n2702_11550.n42 0.376
R13320 a_n2702_11550.n41 a_n2702_11550.n40 0.376
R13321 a_n2702_11550.n127 a_n2702_11550.n124 0.376
R13322 a_n2702_11550.n126 a_n2702_11550.n125 0.376
R13323 a_n2702_11550.n47 a_n2702_11550.n46 0.376
R13324 a_n2702_11550.n51 a_n2702_11550.n50 0.376
R13325 a_n2702_11550.n29 a_n2702_11550.n28 0.349
R13326 a_n2702_11550.n114 a_n2702_11550.n113 0.349
R13327 a_n2702_11550.n94 a_n2702_11550.n93 0.15
R13328 a_n2702_11550.n100 a_n2702_11550.n95 0.148
R13329 a_n2702_11550.n2 a_n2702_11550.n0 0.066
R13330 a_n2702_11550.n84 a_n2702_11550.n83 0.043
R13331 a_n2702_11550.n80 a_n2702_11550.n79 0.043
R13332 a_n2702_11550.n76 a_n2702_11550.n75 0.041
R13333 a_n2702_11550.n91 a_n2702_11550.n90 0.035
R13334 a_n2702_11550.n106 a_n2702_11550.n105 0.035
R13335 a_n2702_11550.n19 a_n2702_11550.n18 0.034
R13336 a_n2702_11550.n23 a_n2702_11550.n22 0.034
R13337 a_n2702_11550.n8 a_n2702_11550.n7 0.034
R13338 a_n2702_11550.n89 a_n2702_11550.n88 0.034
R13339 a_n2702_11550.n104 a_n2702_11550.n103 0.034
R13340 a_n2702_11550.n12 a_n2702_11550.n6 0.032
R13341 a_n2702_11550.n107 a_n2702_11550.n82 0.032
R13342 a_n2702_11550.n9 a_n2702_11550.n8 0.03
R13343 a_n2702_11550.n87 a_n2702_11550.n86 0.03
R13344 a_n2702_11550.n11 a_n2702_11550.n10 0.028
R13345 a_n2702_11550.n72 a_n2702_11550.n70 0.028
R13346 a_n2702_11550.n85 a_n2702_11550.n84 0.028
R13347 a_n2702_11550.n13 a_n2702_11550.n12 0.028
R13348 a_n2702_11550.n69 a_n2702_11550.n68 0.028
R13349 a_n2702_11550.n81 a_n2702_11550.n80 0.028
R13350 a_n2702_11550.n102 a_n2702_11550.n94 0.028
R13351 a_n2702_11550.n17 a_n2702_11550.n15 0.026
R13352 a_n2702_11550.n78 a_n2702_11550.n77 0.026
R13353 a_n2702_11550.n4 a_n2702_11550.n3 0.026
R13354 a_n2702_11550.n18 a_n2702_11550.n17 0.024
R13355 a_n2702_11550.n6 a_n2702_11550.n5 0.024
R13356 a_n2702_11550.n15 a_n2702_11550.n16 0.022
R13357 a_n2702_11550.n5 a_n2702_11550.n4 0.022
R13358 a_n2702_11550.n3 a_n2702_11550.n2 0.022
R13359 a_n2702_11550.n20 a_n2702_11550.n19 0.02
R13360 a_n2702_11550.n10 a_n2702_11550.n9 0.02
R13361 a_n2702_11550.n14 a_n2702_11550.n13 0.02
R13362 a_n2702_11550.n101 a_n2702_11550.n100 0.018
R13363 a_n2702_11550.n82 a_n2702_11550.n81 0.018
R13364 a_n2702_11550.n24 a_n2702_11550.n23 0.017
R13365 a_n2702_11550.n86 a_n2702_11550.n85 0.017
R13366 a_n2702_11550.n70 a_n2702_11550.n71 0.015
R13367 a_n2702_11550.n73 a_n2702_11550.n72 0.015
R13368 a_n2702_11550.n68 a_n2702_11550.n0 0.015
R13369 a_n2702_11550.n75 a_n2702_11550.n69 0.015
R13370 a_n2702_11550.n92 a_n2702_11550.n91 0.013
R13371 a_n2702_11550.n90 a_n2702_11550.n89 0.013
R13372 a_n2702_11550.n107 a_n2702_11550.n106 0.013
R13373 a_n2702_11550.n105 a_n2702_11550.n104 0.013
R13374 a_n2702_11550.n95 a_n2702_11550.n96 0.007
R13375 a_n2702_11550.n21 a_n2702_11550.n20 1.424
R13376 a_n2702_11550.n79 a_n2702_11550.n76 0.005
R13377 a_n2702_11550.n92 a_n2702_11550.n87 0.003
R13378 a_n2702_11550.n103 a_n2702_11550.n102 0.003
R13379 a_n2702_11550.n14 a_n2702_11550.n21 0.47
R13380 a_n4084_12278.n40 a_n4084_12278.t3 732.457
R13381 a_n4084_12278.n40 a_n4084_12278.t2 397.579
R13382 a_n4084_12278.n46 a_n4084_12278.n45 92.5
R13383 a_n4084_12278.n64 a_n4084_12278.n63 92.5
R13384 a_n4084_12278.n45 a_n4084_12278.t1 70.344
R13385 a_n4084_12278.n53 a_n4084_12278.n52 31.034
R13386 a_n4084_12278.n76 a_n4084_12278.n75 31.034
R13387 a_n4084_12278.n1 a_n4084_12278.n57 9.3
R13388 a_n4084_12278.n0 a_n4084_12278.n79 9.3
R13389 a_n4084_12278.n77 a_n4084_12278.n76 9.3
R13390 a_n4084_12278.n54 a_n4084_12278.n53 9.3
R13391 a_n4084_12278.n103 a_n4084_12278.n90 9.154
R13392 a_n4084_12278.n103 a_n4084_12278.n7 9.143
R13393 a_n4084_12278.n103 a_n4084_12278.n6 9.143
R13394 a_n4084_12278.n103 a_n4084_12278.n22 9.132
R13395 a_n4084_12278.n103 a_n4084_12278.n96 9.132
R13396 a_n4084_12278.n103 a_n4084_12278.n100 8.886
R13397 a_n4084_12278.n103 a_n4084_12278.n26 8.885
R13398 a_n4084_12278.n103 a_n4084_12278.n11 8.875
R13399 a_n4084_12278.n103 a_n4084_12278.n32 8.875
R13400 a_n4084_12278.n103 a_n4084_12278.n102 8.864
R13401 a_n4084_12278.n103 a_n4084_12278.n28 8.864
R13402 a_n4084_12278.n47 a_n4084_12278.n46 8.282
R13403 a_n4084_12278.n65 a_n4084_12278.n64 8.282
R13404 a_n4084_12278.t0 a_n4084_12278.n103 7.141
R13405 a_n4084_12278.n54 a_n4084_12278.n50 5.647
R13406 a_n4084_12278.n77 a_n4084_12278.n73 5.647
R13407 a_n4084_12278.n84 a_n4084_12278.n83 4.723
R13408 a_n4084_12278.n2 a_n4084_12278.n62 4.65
R13409 a_n4084_12278.n90 a_n4084_12278.n85 4.65
R13410 a_n4084_12278.n83 a_n4084_12278.n3 4.566
R13411 a_n4084_12278.n90 a_n4084_12278.n39 4.517
R13412 a_n4084_12278.n66 a_n4084_12278.n65 4.5
R13413 a_n4084_12278.n67 a_n4084_12278.n69 4.5
R13414 a_n4084_12278.n43 a_n4084_12278.n47 4.5
R13415 a_n4084_12278.n70 a_n4084_12278.n78 4.5
R13416 a_n4084_12278.n2 a_n4084_12278.n61 4.5
R13417 a_n4084_12278.n4 a_n4084_12278.n56 4.5
R13418 a_n4084_12278.n0 a_n4084_12278.n82 4.5
R13419 a_n4084_12278.n1 a_n4084_12278.n60 4.5
R13420 a_n4084_12278.n98 a_n4084_12278.n97 4.141
R13421 a_n4084_12278.n90 a_n4084_12278.n38 4.141
R13422 a_n4084_12278.n24 a_n4084_12278.n23 4.141
R13423 a_n4084_12278.n52 a_n4084_12278.n51 4.137
R13424 a_n4084_12278.n75 a_n4084_12278.n74 4.137
R13425 a_n4084_12278.n60 a_n4084_12278.n58 3.764
R13426 a_n4084_12278.n78 a_n4084_12278.n71 3.764
R13427 a_n4084_12278.n92 a_n4084_12278.n91 3.764
R13428 a_n4084_12278.n7 a_n4084_12278.n34 3.764
R13429 a_n4084_12278.n96 a_n4084_12278.n95 3.736
R13430 a_n4084_12278.n56 a_n4084_12278.n55 3.388
R13431 a_n4084_12278.n82 a_n4084_12278.n81 3.388
R13432 a_n4084_12278.n9 a_n4084_12278.n8 3.388
R13433 a_n4084_12278.n6 a_n4084_12278.n13 3.388
R13434 a_n4084_12278.n18 a_n4084_12278.n17 3.388
R13435 a_n4084_12278.n30 a_n4084_12278.n29 3.388
R13436 a_n4084_12278.n22 a_n4084_12278.n21 3.36
R13437 a_n4084_12278.n56 a_n4084_12278.n54 3.011
R13438 a_n4084_12278.n47 a_n4084_12278.n44 3.011
R13439 a_n4084_12278.n82 a_n4084_12278.n80 3.011
R13440 a_n4084_12278.n10 a_n4084_12278.n9 3.011
R13441 a_n4084_12278.n13 a_n4084_12278.n12 3.011
R13442 a_n4084_12278.n16 a_n4084_12278.n15 3.011
R13443 a_n4084_12278.n21 a_n4084_12278.n20 3.011
R13444 a_n4084_12278.n19 a_n4084_12278.n18 3.011
R13445 a_n4084_12278.n31 a_n4084_12278.n30 3.011
R13446 a_n4084_12278.n60 a_n4084_12278.n59 2.635
R13447 a_n4084_12278.n69 a_n4084_12278.n68 2.635
R13448 a_n4084_12278.n78 a_n4084_12278.n77 2.635
R13449 a_n4084_12278.n93 a_n4084_12278.n92 2.635
R13450 a_n4084_12278.n95 a_n4084_12278.n94 2.635
R13451 a_n4084_12278.n37 a_n4084_12278.n36 2.635
R13452 a_n4084_12278.n34 a_n4084_12278.n33 2.635
R13453 a_n4084_12278.n83 a_n4084_12278.n40 2.349
R13454 a_n4084_12278.n99 a_n4084_12278.n98 2.258
R13455 a_n4084_12278.n25 a_n4084_12278.n24 2.258
R13456 a_n4084_12278.n5 a_n4084_12278.n89 1.619
R13457 a_n4084_12278.n86 a_n4084_12278.n87 1.588
R13458 a_n4084_12278.n5 a_n4084_12278.n104 1.88
R13459 a_n4084_12278.n3 a_n4084_12278.n0 2.375
R13460 a_n4084_12278.n7 a_n4084_12278.n37 2.257
R13461 a_n4084_12278.n6 a_n4084_12278.n16 2.257
R13462 a_n4084_12278.n36 a_n4084_12278.n35 1.505
R13463 a_n4084_12278.n42 a_n4084_12278.n1 1.5
R13464 a_n4084_12278.n15 a_n4084_12278.n14 1.129
R13465 a_n4084_12278.n50 a_n4084_12278.n49 0.752
R13466 a_n4084_12278.n73 a_n4084_12278.n72 0.752
R13467 a_n4084_12278.n42 a_n4084_12278.n41 0.24
R13468 a_n4084_12278.n102 a_n4084_12278.n101 0.155
R13469 a_n4084_12278.n28 a_n4084_12278.n27 0.155
R13470 a_n4084_12278.n11 a_n4084_12278.n10 0.144
R13471 a_n4084_12278.n32 a_n4084_12278.n31 0.144
R13472 a_n4084_12278.n100 a_n4084_12278.n99 0.133
R13473 a_n4084_12278.n26 a_n4084_12278.n25 0.132
R13474 a_n4084_12278.n67 a_n4084_12278.n66 0.082
R13475 a_n4084_12278.n43 a_n4084_12278.n48 0.071
R13476 a_n4084_12278.n70 a_n4084_12278.n67 0.042
R13477 a_n4084_12278.n87 a_n4084_12278.n88 0.024
R13478 a_n4084_12278.n22 a_n4084_12278.n19 0.024
R13479 a_n4084_12278.n96 a_n4084_12278.n93 0.024
R13480 a_n4084_12278.n85 a_n4084_12278.n86 0.147
R13481 a_n4084_12278.n86 a_n4084_12278.n5 0.124
R13482 a_n4084_12278.n85 a_n4084_12278.n84 2.702
R13483 a_n4084_12278.n3 a_n4084_12278.n42 0.955
R13484 a_n4084_12278.n0 a_n4084_12278.n70 0.127
R13485 a_n4084_12278.n1 a_n4084_12278.n4 0.11
R13486 a_n4084_12278.n4 a_n4084_12278.n43 0.058
R13487 a_n4084_12278.n66 a_n4084_12278.n2 0.042
R13488 a_n11697_12356.n60 a_n11697_12356.t2 735.927
R13489 a_n11697_12356.n54 a_n11697_12356.t5 396.757
R13490 a_n11697_12356.n66 a_n11697_12356.t4 396.757
R13491 a_n11697_12356.n80 a_n11697_12356.n79 92.5
R13492 a_n11697_12356.n98 a_n11697_12356.n97 92.5
R13493 a_n11697_12356.n79 a_n11697_12356.t1 70.344
R13494 a_n11697_12356.n87 a_n11697_12356.n86 31.034
R13495 a_n11697_12356.n110 a_n11697_12356.n109 31.034
R13496 a_n11697_12356.n1 a_n11697_12356.n91 9.3
R13497 a_n11697_12356.n0 a_n11697_12356.n113 9.3
R13498 a_n11697_12356.n111 a_n11697_12356.n110 9.3
R13499 a_n11697_12356.n88 a_n11697_12356.n87 9.3
R13500 a_n11697_12356.n137 a_n11697_12356.n124 9.154
R13501 a_n11697_12356.n137 a_n11697_12356.n7 9.143
R13502 a_n11697_12356.n137 a_n11697_12356.n6 9.143
R13503 a_n11697_12356.n137 a_n11697_12356.n30 9.132
R13504 a_n11697_12356.n137 a_n11697_12356.n130 9.132
R13505 a_n11697_12356.n137 a_n11697_12356.n134 8.886
R13506 a_n11697_12356.n137 a_n11697_12356.n34 8.885
R13507 a_n11697_12356.n137 a_n11697_12356.n19 8.875
R13508 a_n11697_12356.n137 a_n11697_12356.n40 8.875
R13509 a_n11697_12356.n137 a_n11697_12356.n136 8.864
R13510 a_n11697_12356.n137 a_n11697_12356.n36 8.864
R13511 a_n11697_12356.n81 a_n11697_12356.n80 8.282
R13512 a_n11697_12356.n99 a_n11697_12356.n98 8.282
R13513 a_n11697_12356.t0 a_n11697_12356.n137 7.141
R13514 a_n11697_12356.n118 a_n11697_12356.n117 6.621
R13515 a_n11697_12356.n88 a_n11697_12356.n84 5.647
R13516 a_n11697_12356.n111 a_n11697_12356.n107 5.647
R13517 a_n11697_12356.n2 a_n11697_12356.n96 4.65
R13518 a_n11697_12356.n124 a_n11697_12356.n119 4.65
R13519 a_n11697_12356.n124 a_n11697_12356.n47 4.517
R13520 a_n11697_12356.n100 a_n11697_12356.n99 4.5
R13521 a_n11697_12356.n101 a_n11697_12356.n103 4.5
R13522 a_n11697_12356.n77 a_n11697_12356.n81 4.5
R13523 a_n11697_12356.n104 a_n11697_12356.n112 4.5
R13524 a_n11697_12356.n2 a_n11697_12356.n95 4.5
R13525 a_n11697_12356.n4 a_n11697_12356.n90 4.5
R13526 a_n11697_12356.n0 a_n11697_12356.n116 4.5
R13527 a_n11697_12356.n1 a_n11697_12356.n94 4.5
R13528 a_n11697_12356.n132 a_n11697_12356.n131 4.141
R13529 a_n11697_12356.n124 a_n11697_12356.n46 4.141
R13530 a_n11697_12356.n32 a_n11697_12356.n31 4.141
R13531 a_n11697_12356.n86 a_n11697_12356.n85 4.137
R13532 a_n11697_12356.n109 a_n11697_12356.n108 4.137
R13533 a_n11697_12356.n94 a_n11697_12356.n92 3.764
R13534 a_n11697_12356.n112 a_n11697_12356.n105 3.764
R13535 a_n11697_12356.n126 a_n11697_12356.n125 3.764
R13536 a_n11697_12356.n7 a_n11697_12356.n42 3.764
R13537 a_n11697_12356.n13 a_n11697_12356.n55 3.758
R13538 a_n11697_12356.n130 a_n11697_12356.n129 3.736
R13539 a_n11697_12356.n12 a_n11697_12356.n66 3.633
R13540 a_n11697_12356.n90 a_n11697_12356.n89 3.388
R13541 a_n11697_12356.n116 a_n11697_12356.n115 3.388
R13542 a_n11697_12356.n17 a_n11697_12356.n16 3.388
R13543 a_n11697_12356.n6 a_n11697_12356.n21 3.388
R13544 a_n11697_12356.n26 a_n11697_12356.n25 3.388
R13545 a_n11697_12356.n38 a_n11697_12356.n37 3.388
R13546 a_n11697_12356.n30 a_n11697_12356.n29 3.36
R13547 a_n11697_12356.n90 a_n11697_12356.n88 3.011
R13548 a_n11697_12356.n81 a_n11697_12356.n78 3.011
R13549 a_n11697_12356.n116 a_n11697_12356.n114 3.011
R13550 a_n11697_12356.n18 a_n11697_12356.n17 3.011
R13551 a_n11697_12356.n21 a_n11697_12356.n20 3.011
R13552 a_n11697_12356.n24 a_n11697_12356.n23 3.011
R13553 a_n11697_12356.n29 a_n11697_12356.n28 3.011
R13554 a_n11697_12356.n27 a_n11697_12356.n26 3.011
R13555 a_n11697_12356.n39 a_n11697_12356.n38 3.011
R13556 a_n11697_12356.n94 a_n11697_12356.n93 2.635
R13557 a_n11697_12356.n103 a_n11697_12356.n102 2.635
R13558 a_n11697_12356.n112 a_n11697_12356.n111 2.635
R13559 a_n11697_12356.n127 a_n11697_12356.n126 2.635
R13560 a_n11697_12356.n129 a_n11697_12356.n128 2.635
R13561 a_n11697_12356.n45 a_n11697_12356.n44 2.635
R13562 a_n11697_12356.n42 a_n11697_12356.n41 2.635
R13563 a_n11697_12356.n117 a_n11697_12356.n3 2.631
R13564 a_n11697_12356.n74 a_n11697_12356.n71 2.621
R13565 a_n11697_12356.n15 a_n11697_12356.n54 3.627
R13566 a_n11697_12356.n133 a_n11697_12356.n132 2.258
R13567 a_n11697_12356.n33 a_n11697_12356.n32 2.258
R13568 a_n11697_12356.n5 a_n11697_12356.n123 1.619
R13569 a_n11697_12356.n120 a_n11697_12356.n121 1.588
R13570 a_n11697_12356.n5 a_n11697_12356.n138 1.88
R13571 a_n11697_12356.n3 a_n11697_12356.n0 2.375
R13572 a_n11697_12356.n44 a_n11697_12356.n43 1.505
R13573 a_n11697_12356.n76 a_n11697_12356.n1 1.5
R13574 a_n11697_12356.n7 a_n11697_12356.n45 2.257
R13575 a_n11697_12356.n6 a_n11697_12356.n24 2.257
R13576 a_n11697_12356.n9 a_n11697_12356.n8 1.149
R13577 a_n11697_12356.n59 a_n11697_12356.n57 1.149
R13578 a_n11697_12356.n11 a_n11697_12356.n10 1.149
R13579 a_n11697_12356.n12 a_n11697_12356.n63 1.148
R13580 a_n11697_12356.n15 a_n11697_12356.n9 1.138
R13581 a_n11697_12356.n14 a_n11697_12356.t3 737.066
R13582 a_n11697_12356.n63 a_n11697_12356.n61 1.137
R13583 a_n11697_12356.n11 a_n11697_12356.n67 1.137
R13584 a_n11697_12356.n14 a_n11697_12356.n74 1.136
R13585 a_n11697_12356.n13 a_n11697_12356.n59 1.136
R13586 a_n11697_12356.n23 a_n11697_12356.n22 1.129
R13587 a_n11697_12356.n84 a_n11697_12356.n83 0.752
R13588 a_n11697_12356.n107 a_n11697_12356.n106 0.752
R13589 a_n11697_12356.n9 a_n11697_12356.n48 1.149
R13590 a_n11697_12356.n14 a_n11697_12356.n11 1.148
R13591 a_n11697_12356.n76 a_n11697_12356.n75 0.24
R13592 a_n11697_12356.n136 a_n11697_12356.n135 0.155
R13593 a_n11697_12356.n36 a_n11697_12356.n35 0.155
R13594 a_n11697_12356.n19 a_n11697_12356.n18 0.144
R13595 a_n11697_12356.n40 a_n11697_12356.n39 0.144
R13596 a_n11697_12356.n134 a_n11697_12356.n133 0.133
R13597 a_n11697_12356.n34 a_n11697_12356.n33 0.132
R13598 a_n11697_12356.n54 a_n11697_12356.n52 0.126
R13599 a_n11697_12356.n66 a_n11697_12356.n64 0.126
R13600 a_n11697_12356.n13 a_n11697_12356.n15 0.114
R13601 a_n11697_12356.n14 a_n11697_12356.n12 0.11
R13602 a_n11697_12356.n12 a_n11697_12356.n13 0.106
R13603 a_n11697_12356.n101 a_n11697_12356.n100 0.082
R13604 a_n11697_12356.n77 a_n11697_12356.n82 0.071
R13605 a_n11697_12356.n104 a_n11697_12356.n101 0.042
R13606 a_n11697_12356.n59 a_n11697_12356.n60 0.059
R13607 a_n11697_12356.n8 a_n11697_12356.n50 0.032
R13608 a_n11697_12356.n10 a_n11697_12356.n69 0.032
R13609 a_n11697_12356.n52 a_n11697_12356.n53 0.028
R13610 a_n11697_12356.n48 a_n11697_12356.n49 0.028
R13611 a_n11697_12356.n8 a_n11697_12356.n51 0.028
R13612 a_n11697_12356.n55 a_n11697_12356.n56 0.028
R13613 a_n11697_12356.n57 a_n11697_12356.n58 0.028
R13614 a_n11697_12356.n64 a_n11697_12356.n65 0.028
R13615 a_n11697_12356.n61 a_n11697_12356.n62 0.028
R13616 a_n11697_12356.n71 a_n11697_12356.n72 0.028
R13617 a_n11697_12356.n67 a_n11697_12356.n68 0.028
R13618 a_n11697_12356.n10 a_n11697_12356.n70 0.028
R13619 a_n11697_12356.n74 a_n11697_12356.n73 0.027
R13620 a_n11697_12356.n121 a_n11697_12356.n122 0.024
R13621 a_n11697_12356.n30 a_n11697_12356.n27 0.024
R13622 a_n11697_12356.n130 a_n11697_12356.n127 0.024
R13623 a_n11697_12356.n119 a_n11697_12356.n120 0.147
R13624 a_n11697_12356.n120 a_n11697_12356.n5 0.124
R13625 a_n11697_12356.n117 a_n11697_12356.n14 0.071
R13626 a_n11697_12356.n119 a_n11697_12356.n118 2.702
R13627 a_n11697_12356.n3 a_n11697_12356.n76 0.955
R13628 a_n11697_12356.n0 a_n11697_12356.n104 0.127
R13629 a_n11697_12356.n1 a_n11697_12356.n4 0.11
R13630 a_n11697_12356.n4 a_n11697_12356.n77 0.058
R13631 a_n11697_12356.n100 a_n11697_12356.n2 0.042
R13632 modi2.n261 modi2.t4 1037.92
R13633 modi2.n258 modi2.t2 1037.28
R13634 modi2.n258 modi2.t3 797.528
R13635 modi2.n261 modi2.t5 796.887
R13636 modi2.n31 modi2.n30 92.5
R13637 modi2.n59 modi2.n58 92.5
R13638 modi2.n58 modi2.t1 70.344
R13639 modi2.n19 modi2.n18 31.034
R13640 modi2.n50 modi2.n49 31.034
R13641 modi2.n114 modi2.n113 9.3
R13642 modi2.n191 modi2.n190 9.3
R13643 modi2.n3 modi2.n2 9.3
R13644 modi2.n51 modi2.n50 9.3
R13645 modi2.n20 modi2.n19 9.3
R13646 modi2.n78 modi2.n77 9.3
R13647 modi2.n230 modi2.n229 9.154
R13648 modi2.n32 modi2.n31 8.282
R13649 modi2.n60 modi2.n59 8.282
R13650 modi2.n229 modi2.t0 7.141
R13651 modi2.n150 modi2.n149 7.033
R13652 modi2.n93 modi2.n92 7.033
R13653 modi2.n259 modi2.n257 6.416
R13654 modi2.n20 modi2.n16 5.647
R13655 modi2.n51 modi2.n47 5.647
R13656 modi2.n231 modi2.n230 4.65
R13657 modi2.n57 modi2.n56 4.65
R13658 modi2.n177 modi2.n176 4.5
R13659 modi2.n197 modi2.n196 4.5
R13660 modi2.n210 modi2.n209 4.5
R13661 modi2.n217 modi2.n214 4.5
R13662 modi2.n226 modi2.n225 4.5
R13663 modi2.n232 modi2.n228 4.5
R13664 modi2.n101 modi2.n98 4.5
R13665 modi2.n108 modi2.n107 4.5
R13666 modi2.n120 modi2.n119 4.5
R13667 modi2.n130 modi2.n129 4.5
R13668 modi2.n140 modi2.n139 4.5
R13669 modi2.n164 modi2.n163 4.5
R13670 modi2.n84 modi2.n82 4.5
R13671 modi2.n55 modi2.n52 4.5
R13672 modi2.n70 modi2.n68 4.5
R13673 modi2.n33 modi2.n32 4.5
R13674 modi2.n40 modi2.n39 4.5
R13675 modi2.n61 modi2.n60 4.5
R13676 modi2.n23 modi2.n22 4.5
R13677 modi2.n8 modi2.n7 4.5
R13678 modi2.n129 modi2.n126 4.141
R13679 modi2.n163 modi2.n162 4.141
R13680 modi2.n18 modi2.n17 4.137
R13681 modi2.n49 modi2.n48 4.137
R13682 modi2.n302 modi2.n259 3.857
R13683 modi2.n119 modi2.n116 3.764
R13684 modi2.n209 modi2.n207 3.764
R13685 modi2.n7 modi2.n5 3.764
R13686 modi2.n52 modi2.n45 3.764
R13687 modi2.n264 modi2.n261 3.463
R13688 modi2.n139 modi2.n136 3.388
R13689 modi2.n107 modi2.n106 3.388
R13690 modi2.n196 modi2.n195 3.388
R13691 modi2.n176 modi2.n175 3.388
R13692 modi2.n22 modi2.n21 3.388
R13693 modi2.n82 modi2.n81 3.388
R13694 modi2.n139 modi2.n138 3.011
R13695 modi2.n107 modi2.n104 3.011
R13696 modi2.n98 modi2.n96 3.011
R13697 modi2.n190 modi2.n189 3.011
R13698 modi2.n196 modi2.n194 3.011
R13699 modi2.n176 modi2.n174 3.011
R13700 modi2.n22 modi2.n20 3.011
R13701 modi2.n32 modi2.n29 3.011
R13702 modi2.n82 modi2.n80 3.011
R13703 modi2.n119 modi2.n118 2.635
R13704 modi2.n113 modi2.n112 2.635
R13705 modi2.n214 modi2.n213 2.635
R13706 modi2.n209 modi2.n208 2.635
R13707 modi2.n7 modi2.n6 2.635
R13708 modi2.n68 modi2.n67 2.635
R13709 modi2.n52 modi2.n51 2.635
R13710 modi2.n129 modi2.n128 2.258
R13711 modi2.n163 modi2.n161 2.258
R13712 modi2.n259 modi2.n258 2.25
R13713 modi2.n26 modi2.n0 1.754
R13714 modi2.n180 modi2.n151 1.754
R13715 modi2.n26 modi2.n25 1.705
R13716 modi2.n43 modi2.n42 1.705
R13717 modi2.n73 modi2.n72 1.705
R13718 modi2.n87 modi2.n86 1.705
R13719 modi2.n256 modi2.n145 1.705
R13720 modi2.n200 modi2.n199 1.705
R13721 modi2.n220 modi2.n219 1.705
R13722 modi2.n249 modi2.n248 1.705
R13723 modi2.n255 modi2.n254 1.705
R13724 modi2.n243 modi2.n242 1.705
R13725 modi2.n237 modi2.n236 1.705
R13726 modi2.n186 modi2.n185 1.705
R13727 modi2.n180 modi2.n179 1.705
R13728 modi2.n214 modi2.n212 1.505
R13729 modi2.n198 modi2.n197 1.5
R13730 modi2.n211 modi2.n210 1.5
R13731 modi2.n218 modi2.n217 1.5
R13732 modi2.n227 modi2.n226 1.5
R13733 modi2.n233 modi2.n232 1.5
R13734 modi2.n85 modi2.n84 1.5
R13735 modi2.n72 modi2.n55 1.5
R13736 modi2.n34 modi2.n33 1.5
R13737 modi2.n71 modi2.n70 1.5
R13738 modi2.n41 modi2.n40 1.5
R13739 modi2.n62 modi2.n61 1.5
R13740 modi2.n24 modi2.n23 1.5
R13741 modi2.n9 modi2.n8 1.5
R13742 modi2.n298 modi2.n297 1.402
R13743 modi2.n265 modi2.n264 1.355
R13744 modi2.n257 modi2.n256 1.267
R13745 modi2.n299 modi2.n298 1.14
R13746 modi2.n277 modi2.n276 1.137
R13747 modi2.n288 modi2.n287 1.137
R13748 modi2.n281 modi2.n280 1.137
R13749 modi2.n271 modi2.n270 1.137
R13750 modi2.n266 modi2.n265 1.137
R13751 modi2.n98 modi2.n97 1.129
R13752 modi2.n151 modi2.n150 1.127
R13753 modi2.n145 modi2.n93 1.127
R13754 modi2.n141 modi2.n140 1.125
R13755 modi2.n178 modi2.n177 1.125
R13756 modi2.n16 modi2.n15 0.752
R13757 modi2.n47 modi2.n46 0.752
R13758 modi2.n257 modi2.n87 0.71
R13759 modi2.n300 modi2.n299 0.686
R13760 modi2.n92 modi2.n91 0.155
R13761 modi2.n149 modi2.n148 0.155
R13762 modi2.n138 modi2.n137 0.144
R13763 modi2.n174 modi2.n173 0.144
R13764 modi2.n128 modi2.n127 0.133
R13765 modi2.n161 modi2.n160 0.132
R13766 modi2.n134 modi2.n133 0.053
R13767 modi2.n124 modi2.n123 0.053
R13768 modi2.n114 modi2.n111 0.053
R13769 modi2.n158 modi2.n157 0.053
R13770 modi2.n168 modi2.n167 0.053
R13771 modi2.n171 modi2.n170 0.053
R13772 modi2.n78 modi2.n76 0.053
R13773 modi2.n43 modi2.n26 0.049
R13774 modi2.n73 modi2.n43 0.049
R13775 modi2.n87 modi2.n73 0.049
R13776 modi2.n256 modi2.n255 0.049
R13777 modi2.n255 modi2.n249 0.049
R13778 modi2.n249 modi2.n243 0.049
R13779 modi2.n243 modi2.n237 0.049
R13780 modi2.n237 modi2.n220 0.049
R13781 modi2.n220 modi2.n200 0.049
R13782 modi2.n200 modi2.n186 0.049
R13783 modi2.n186 modi2.n180 0.049
R13784 modi2.n264 modi2.n263 0.048
R13785 modi2.n40 modi2.n38 0.045
R13786 modi2.n70 modi2.n66 0.045
R13787 modi2.n101 modi2.n100 0.043
R13788 modi2.n226 modi2.n224 0.043
R13789 modi2.n294 modi2.n293 0.037
R13790 modi2.n89 modi2.n88 0.034
R13791 modi2.n167 modi2.n166 0.032
R13792 modi2.n135 modi2.n134 0.03
R13793 modi2.n133 modi2.n132 0.03
R13794 modi2.n157 modi2.n156 0.03
R13795 modi2.n10 modi2.n9 0.03
R13796 modi2.n85 modi2.n75 0.03
R13797 modi2.n123 modi2.n122 0.028
R13798 modi2.n169 modi2.n168 0.028
R13799 modi2.n172 modi2.n171 0.028
R13800 modi2.n95 modi2.n94 0.025
R13801 modi2.n125 modi2.n124 0.025
R13802 modi2.n61 modi2.n57 0.025
R13803 modi2.n118 modi2.n117 0.024
R13804 modi2.n194 modi2.n193 0.024
R13805 modi2.n232 modi2.n231 0.023
R13806 modi2.n159 modi2.n158 0.023
R13807 modi2.n121 modi2.n120 0.021
R13808 modi2.n115 modi2.n114 0.021
R13809 modi2.n204 modi2.n203 0.021
R13810 modi2.n8 modi2.n1 0.021
R13811 modi2.n4 modi2.n3 0.021
R13812 modi2.n55 modi2.n44 0.021
R13813 modi2.n280 modi2.n279 0.021
R13814 modi2.n140 modi2.n95 0.019
R13815 modi2.n111 modi2.n110 0.019
R13816 modi2.n110 modi2.n109 0.019
R13817 modi2.n108 modi2.n103 0.019
R13818 modi2.n205 modi2.n204 0.019
R13819 modi2.n192 modi2.n191 0.019
R13820 modi2.n177 modi2.n172 0.019
R13821 modi2.n199 modi2.n198 0.019
R13822 modi2.n13 modi2.n12 0.019
R13823 modi2.n14 modi2.n13 0.019
R13824 modi2.n54 modi2.n53 0.019
R13825 modi2.n79 modi2.n78 0.019
R13826 modi2.n84 modi2.n83 0.019
R13827 modi2.n93 modi2.n90 0.019
R13828 modi2.n150 modi2.n147 0.019
R13829 modi2.n287 modi2.n286 0.018
R13830 modi2.n276 modi2.n275 0.018
R13831 modi2.n140 modi2.n135 0.017
R13832 modi2.n131 modi2.n130 0.017
R13833 modi2.n109 modi2.n108 0.017
R13834 modi2.n102 modi2.n101 0.017
R13835 modi2.n197 modi2.n192 0.017
R13836 modi2.n165 modi2.n164 0.017
R13837 modi2.n177 modi2.n169 0.017
R13838 modi2.n23 modi2.n14 0.017
R13839 modi2.n33 modi2.n28 0.017
R13840 modi2.n84 modi2.n79 0.017
R13841 modi2.n143 modi2.n142 0.016
R13842 modi2.n253 modi2.n252 0.016
R13843 modi2.n247 modi2.n246 0.016
R13844 modi2.n182 modi2.n181 0.016
R13845 modi2.n154 modi2.n153 0.016
R13846 modi2.n297 modi2.n296 0.016
R13847 modi2.n295 modi2.n294 0.016
R13848 modi2.n293 modi2.n292 0.016
R13849 modi2.n263 modi2.n262 0.016
R13850 modi2.n120 modi2.n115 0.015
R13851 modi2.n217 modi2.n216 0.015
R13852 modi2.n210 modi2.n205 0.015
R13853 modi2.n239 modi2.n238 0.015
R13854 modi2.n233 modi2.n227 0.015
R13855 modi2.n218 modi2.n211 0.015
R13856 modi2.n8 modi2.n4 0.015
R13857 modi2.n70 modi2.n69 0.015
R13858 modi2.n55 modi2.n54 0.015
R13859 modi2.n41 modi2.n36 0.015
R13860 modi2.n71 modi2.n64 0.015
R13861 modi2.n72 modi2.n71 0.015
R13862 modi2.n178 modi2.n154 0.014
R13863 modi2.n35 modi2.n34 0.014
R13864 modi2.n63 modi2.n62 0.014
R13865 modi2.n142 modi2.n141 0.013
R13866 modi2.n234 modi2.n233 0.013
R13867 modi2.n227 modi2.n222 0.013
R13868 modi2.n106 modi2.n105 0.012
R13869 modi2.n207 modi2.n206 0.012
R13870 modi2.n130 modi2.n125 0.012
R13871 modi2.n103 modi2.n102 0.012
R13872 modi2.n216 modi2.n215 0.012
R13873 modi2.n164 modi2.n159 0.012
R13874 modi2.n28 modi2.n27 0.012
R13875 modi2.n144 modi2.n143 0.011
R13876 modi2.n252 modi2.n251 0.011
R13877 modi2.n240 modi2.n239 0.011
R13878 modi2.n219 modi2.n218 0.011
R13879 modi2.n185 modi2.n184 0.011
R13880 modi2.n183 modi2.n182 0.011
R13881 modi2.n153 modi2.n152 0.011
R13882 modi2.n298 modi2.n291 0.011
R13883 modi2.n287 modi2.n284 0.011
R13884 modi2.n270 modi2.n269 0.011
R13885 modi2.n265 modi2.n260 0.011
R13886 modi2.n242 modi2.n241 0.01
R13887 modi2.n211 modi2.n202 0.01
R13888 modi2.n25 modi2.n11 0.01
R13889 modi2.n286 modi2.n285 0.01
R13890 modi2.n275 modi2.n274 0.01
R13891 modi2.n254 modi2.n253 0.009
R13892 modi2.n188 modi2.n187 0.009
R13893 modi2.n283 modi2.n282 0.009
R13894 modi2.n273 modi2.n272 0.009
R13895 modi2.n100 modi2.n99 0.008
R13896 modi2.n224 modi2.n223 0.008
R13897 modi2.n246 modi2.n245 0.008
R13898 modi2.n245 modi2.n244 0.008
R13899 modi2.n38 modi2.n37 0.008
R13900 modi2.n66 modi2.n65 0.008
R13901 modi2.n296 modi2.n295 0.008
R13902 modi2.n198 modi2.n188 0.007
R13903 modi2.n42 modi2.n41 0.007
R13904 modi2.n75 modi2.n74 0.007
R13905 modi2.n86 modi2.n85 0.007
R13906 modi2.n290 modi2.n289 0.007
R13907 modi2.n281 modi2.n278 0.007
R13908 modi2.n278 modi2.n277 0.007
R13909 modi2.n268 modi2.n267 0.007
R13910 modi2.n132 modi2.n131 0.006
R13911 modi2.n122 modi2.n121 0.006
R13912 modi2.n156 modi2.n155 0.006
R13913 modi2.n166 modi2.n165 0.006
R13914 modi2.n202 modi2.n201 0.006
R13915 modi2.n11 modi2.n10 0.006
R13916 modi2.n282 modi2.n281 0.006
R13917 modi2.n277 modi2.n273 0.006
R13918 modi2.n145 modi2.n144 0.005
R13919 modi2.n251 modi2.n250 0.005
R13920 modi2.n241 modi2.n240 0.005
R13921 modi2.n184 modi2.n183 0.005
R13922 modi2.n179 modi2.n178 0.005
R13923 modi2.n90 modi2.n89 0.004
R13924 modi2.n147 modi2.n146 0.004
R13925 modi2.n289 modi2.n288 0.004
R13926 modi2.n271 modi2.n268 0.004
R13927 modi2.n267 modi2.n266 0.004
R13928 modi2.n302 modi2.n301 0.004
R13929 modi2.n303 modi2.n302 0.004
R13930 modi2.n305 modi2.n304 0.004
R13931 modi2.n306 modi2.n305 0.004
R13932 modi2 modi2.n306 0.004
R13933 modi2.n236 modi2.n235 0.003
R13934 modi2.n235 modi2.n234 0.002
R13935 modi2.n222 modi2.n221 0.002
R13936 modi2.n36 modi2.n35 0.002
R13937 modi2.n64 modi2.n63 0.002
R13938 modi2.n288 modi2.n283 0.002
R13939 modi2.n272 modi2.n271 0.002
R13940 modi2.n301 modi2.n300 0.002
R13941 modi2.n304 modi2.n303 0.002
R13942 modi2.n299 modi2.n290 0.001
R13943 modi2.n248 modi2.n247 0.001
R13944 modi2.n25 modi2.n24 0.001
R13945 a_n23348_12347.n60 a_n23348_12347.t3 735.927
R13946 a_n23348_12347.n54 a_n23348_12347.t2 396.757
R13947 a_n23348_12347.n66 a_n23348_12347.t4 396.757
R13948 a_n23348_12347.n80 a_n23348_12347.n79 92.5
R13949 a_n23348_12347.n98 a_n23348_12347.n97 92.5
R13950 a_n23348_12347.n79 a_n23348_12347.t1 70.344
R13951 a_n23348_12347.n87 a_n23348_12347.n86 31.034
R13952 a_n23348_12347.n110 a_n23348_12347.n109 31.034
R13953 a_n23348_12347.n1 a_n23348_12347.n91 9.3
R13954 a_n23348_12347.n0 a_n23348_12347.n113 9.3
R13955 a_n23348_12347.n111 a_n23348_12347.n110 9.3
R13956 a_n23348_12347.n88 a_n23348_12347.n87 9.3
R13957 a_n23348_12347.n137 a_n23348_12347.n124 9.154
R13958 a_n23348_12347.n137 a_n23348_12347.n7 9.143
R13959 a_n23348_12347.n137 a_n23348_12347.n6 9.143
R13960 a_n23348_12347.n137 a_n23348_12347.n30 9.132
R13961 a_n23348_12347.n137 a_n23348_12347.n130 9.132
R13962 a_n23348_12347.n137 a_n23348_12347.n134 8.886
R13963 a_n23348_12347.n137 a_n23348_12347.n34 8.885
R13964 a_n23348_12347.n137 a_n23348_12347.n19 8.875
R13965 a_n23348_12347.n137 a_n23348_12347.n40 8.875
R13966 a_n23348_12347.n137 a_n23348_12347.n136 8.864
R13967 a_n23348_12347.n137 a_n23348_12347.n36 8.864
R13968 a_n23348_12347.n81 a_n23348_12347.n80 8.282
R13969 a_n23348_12347.n99 a_n23348_12347.n98 8.282
R13970 a_n23348_12347.t0 a_n23348_12347.n137 7.141
R13971 a_n23348_12347.n118 a_n23348_12347.n117 6.622
R13972 a_n23348_12347.n88 a_n23348_12347.n84 5.647
R13973 a_n23348_12347.n111 a_n23348_12347.n107 5.647
R13974 a_n23348_12347.n2 a_n23348_12347.n96 4.65
R13975 a_n23348_12347.n124 a_n23348_12347.n119 4.65
R13976 a_n23348_12347.n124 a_n23348_12347.n47 4.517
R13977 a_n23348_12347.n100 a_n23348_12347.n99 4.5
R13978 a_n23348_12347.n101 a_n23348_12347.n103 4.5
R13979 a_n23348_12347.n77 a_n23348_12347.n81 4.5
R13980 a_n23348_12347.n104 a_n23348_12347.n112 4.5
R13981 a_n23348_12347.n2 a_n23348_12347.n95 4.5
R13982 a_n23348_12347.n4 a_n23348_12347.n90 4.5
R13983 a_n23348_12347.n0 a_n23348_12347.n116 4.5
R13984 a_n23348_12347.n1 a_n23348_12347.n94 4.5
R13985 a_n23348_12347.n132 a_n23348_12347.n131 4.141
R13986 a_n23348_12347.n124 a_n23348_12347.n46 4.141
R13987 a_n23348_12347.n32 a_n23348_12347.n31 4.141
R13988 a_n23348_12347.n86 a_n23348_12347.n85 4.137
R13989 a_n23348_12347.n109 a_n23348_12347.n108 4.137
R13990 a_n23348_12347.n94 a_n23348_12347.n92 3.764
R13991 a_n23348_12347.n112 a_n23348_12347.n105 3.764
R13992 a_n23348_12347.n126 a_n23348_12347.n125 3.764
R13993 a_n23348_12347.n7 a_n23348_12347.n42 3.764
R13994 a_n23348_12347.n13 a_n23348_12347.n55 3.758
R13995 a_n23348_12347.n130 a_n23348_12347.n129 3.736
R13996 a_n23348_12347.n12 a_n23348_12347.n66 3.633
R13997 a_n23348_12347.n90 a_n23348_12347.n89 3.388
R13998 a_n23348_12347.n116 a_n23348_12347.n115 3.388
R13999 a_n23348_12347.n17 a_n23348_12347.n16 3.388
R14000 a_n23348_12347.n6 a_n23348_12347.n21 3.388
R14001 a_n23348_12347.n26 a_n23348_12347.n25 3.388
R14002 a_n23348_12347.n38 a_n23348_12347.n37 3.388
R14003 a_n23348_12347.n30 a_n23348_12347.n29 3.36
R14004 a_n23348_12347.n90 a_n23348_12347.n88 3.011
R14005 a_n23348_12347.n81 a_n23348_12347.n78 3.011
R14006 a_n23348_12347.n116 a_n23348_12347.n114 3.011
R14007 a_n23348_12347.n18 a_n23348_12347.n17 3.011
R14008 a_n23348_12347.n21 a_n23348_12347.n20 3.011
R14009 a_n23348_12347.n24 a_n23348_12347.n23 3.011
R14010 a_n23348_12347.n29 a_n23348_12347.n28 3.011
R14011 a_n23348_12347.n27 a_n23348_12347.n26 3.011
R14012 a_n23348_12347.n39 a_n23348_12347.n38 3.011
R14013 a_n23348_12347.n94 a_n23348_12347.n93 2.635
R14014 a_n23348_12347.n103 a_n23348_12347.n102 2.635
R14015 a_n23348_12347.n112 a_n23348_12347.n111 2.635
R14016 a_n23348_12347.n127 a_n23348_12347.n126 2.635
R14017 a_n23348_12347.n129 a_n23348_12347.n128 2.635
R14018 a_n23348_12347.n45 a_n23348_12347.n44 2.635
R14019 a_n23348_12347.n42 a_n23348_12347.n41 2.635
R14020 a_n23348_12347.n117 a_n23348_12347.n3 2.631
R14021 a_n23348_12347.n74 a_n23348_12347.n71 2.621
R14022 a_n23348_12347.n15 a_n23348_12347.n54 3.627
R14023 a_n23348_12347.n133 a_n23348_12347.n132 2.258
R14024 a_n23348_12347.n33 a_n23348_12347.n32 2.258
R14025 a_n23348_12347.n5 a_n23348_12347.n123 1.619
R14026 a_n23348_12347.n120 a_n23348_12347.n121 1.588
R14027 a_n23348_12347.n5 a_n23348_12347.n138 1.88
R14028 a_n23348_12347.n3 a_n23348_12347.n0 2.375
R14029 a_n23348_12347.n44 a_n23348_12347.n43 1.505
R14030 a_n23348_12347.n76 a_n23348_12347.n1 1.5
R14031 a_n23348_12347.n7 a_n23348_12347.n45 2.257
R14032 a_n23348_12347.n6 a_n23348_12347.n24 2.257
R14033 a_n23348_12347.n9 a_n23348_12347.n8 1.149
R14034 a_n23348_12347.n59 a_n23348_12347.n57 1.149
R14035 a_n23348_12347.n11 a_n23348_12347.n10 1.149
R14036 a_n23348_12347.n12 a_n23348_12347.n63 1.148
R14037 a_n23348_12347.n15 a_n23348_12347.n9 1.138
R14038 a_n23348_12347.n14 a_n23348_12347.t5 737.066
R14039 a_n23348_12347.n63 a_n23348_12347.n61 1.137
R14040 a_n23348_12347.n11 a_n23348_12347.n67 1.137
R14041 a_n23348_12347.n14 a_n23348_12347.n74 1.136
R14042 a_n23348_12347.n13 a_n23348_12347.n59 1.136
R14043 a_n23348_12347.n23 a_n23348_12347.n22 1.129
R14044 a_n23348_12347.n84 a_n23348_12347.n83 0.752
R14045 a_n23348_12347.n107 a_n23348_12347.n106 0.752
R14046 a_n23348_12347.n9 a_n23348_12347.n48 1.149
R14047 a_n23348_12347.n14 a_n23348_12347.n11 1.148
R14048 a_n23348_12347.n76 a_n23348_12347.n75 0.24
R14049 a_n23348_12347.n136 a_n23348_12347.n135 0.155
R14050 a_n23348_12347.n36 a_n23348_12347.n35 0.155
R14051 a_n23348_12347.n19 a_n23348_12347.n18 0.144
R14052 a_n23348_12347.n40 a_n23348_12347.n39 0.144
R14053 a_n23348_12347.n134 a_n23348_12347.n133 0.133
R14054 a_n23348_12347.n34 a_n23348_12347.n33 0.132
R14055 a_n23348_12347.n54 a_n23348_12347.n52 0.126
R14056 a_n23348_12347.n66 a_n23348_12347.n64 0.126
R14057 a_n23348_12347.n13 a_n23348_12347.n15 0.114
R14058 a_n23348_12347.n14 a_n23348_12347.n12 0.11
R14059 a_n23348_12347.n12 a_n23348_12347.n13 0.106
R14060 a_n23348_12347.n101 a_n23348_12347.n100 0.082
R14061 a_n23348_12347.n77 a_n23348_12347.n82 0.071
R14062 a_n23348_12347.n104 a_n23348_12347.n101 0.042
R14063 a_n23348_12347.n59 a_n23348_12347.n60 0.059
R14064 a_n23348_12347.n8 a_n23348_12347.n50 0.032
R14065 a_n23348_12347.n10 a_n23348_12347.n69 0.032
R14066 a_n23348_12347.n52 a_n23348_12347.n53 0.028
R14067 a_n23348_12347.n48 a_n23348_12347.n49 0.028
R14068 a_n23348_12347.n8 a_n23348_12347.n51 0.028
R14069 a_n23348_12347.n55 a_n23348_12347.n56 0.028
R14070 a_n23348_12347.n57 a_n23348_12347.n58 0.028
R14071 a_n23348_12347.n64 a_n23348_12347.n65 0.028
R14072 a_n23348_12347.n61 a_n23348_12347.n62 0.028
R14073 a_n23348_12347.n71 a_n23348_12347.n72 0.028
R14074 a_n23348_12347.n67 a_n23348_12347.n68 0.028
R14075 a_n23348_12347.n10 a_n23348_12347.n70 0.028
R14076 a_n23348_12347.n74 a_n23348_12347.n73 0.027
R14077 a_n23348_12347.n121 a_n23348_12347.n122 0.024
R14078 a_n23348_12347.n30 a_n23348_12347.n27 0.024
R14079 a_n23348_12347.n130 a_n23348_12347.n127 0.024
R14080 a_n23348_12347.n119 a_n23348_12347.n120 0.147
R14081 a_n23348_12347.n120 a_n23348_12347.n5 0.124
R14082 a_n23348_12347.n117 a_n23348_12347.n14 0.071
R14083 a_n23348_12347.n119 a_n23348_12347.n118 2.702
R14084 a_n23348_12347.n3 a_n23348_12347.n76 0.955
R14085 a_n23348_12347.n0 a_n23348_12347.n104 0.127
R14086 a_n23348_12347.n1 a_n23348_12347.n4 0.11
R14087 a_n23348_12347.n4 a_n23348_12347.n77 0.058
R14088 a_n23348_12347.n100 a_n23348_12347.n2 0.042
R14089 modi5.n6 modi5.t3 1037.94
R14090 modi5.n43 modi5.t4 1037.28
R14091 modi5.n43 modi5.t5 797.53
R14092 modi5.n6 modi5.t2 796.922
R14093 modi5.n291 modi5.n290 92.5
R14094 modi5.n263 modi5.n262 92.5
R14095 modi5.n290 modi5.t0 70.344
R14096 modi5.n277 modi5.n276 31.034
R14097 modi5.n243 modi5.n242 31.034
R14098 modi5.n218 modi5.n217 9.3
R14099 modi5.n278 modi5.n277 9.3
R14100 modi5.n244 modi5.n243 9.3
R14101 modi5.n228 modi5.n227 9.3
R14102 modi5.n90 modi5.n89 9.3
R14103 modi5.n172 modi5.n171 9.3
R14104 modi5.n128 modi5.n127 9.154
R14105 modi5.n292 modi5.n291 8.282
R14106 modi5.n264 modi5.n263 8.282
R14107 modi5.n127 modi5.t1 7.141
R14108 modi5.n48 modi5.n47 7.033
R14109 modi5.n210 modi5.n209 7.032
R14110 modi5.n301 modi5.n300 6.465
R14111 modi5.n278 modi5.n274 5.647
R14112 modi5.n244 modi5.n240 5.647
R14113 modi5.n284 modi5.n283 4.65
R14114 modi5.n129 modi5.n128 4.65
R14115 modi5.n234 modi5.n232 4.5
R14116 modi5.n249 modi5.n245 4.5
R14117 modi5.n256 modi5.n253 4.5
R14118 modi5.n281 modi5.n280 4.5
R14119 modi5.n295 modi5.n292 4.5
R14120 modi5.n285 modi5.n282 4.5
R14121 modi5.n265 modi5.n264 4.5
R14122 modi5.n223 modi5.n222 4.5
R14123 modi5.n200 modi5.n199 4.5
R14124 modi5.n188 modi5.n187 4.5
R14125 modi5.n178 modi5.n177 4.5
R14126 modi5.n166 modi5.n165 4.5
R14127 modi5.n159 modi5.n158 4.5
R14128 modi5.n131 modi5.n130 4.5
R14129 modi5.n125 modi5.n124 4.5
R14130 modi5.n116 modi5.n115 4.5
R14131 modi5.n109 modi5.n108 4.5
R14132 modi5.n96 modi5.n95 4.5
R14133 modi5.n65 modi5.n64 4.5
R14134 modi5.n75 modi5.n74 4.5
R14135 modi5.n64 modi5.n61 4.141
R14136 modi5.n187 modi5.n186 4.141
R14137 modi5.n276 modi5.n275 4.137
R14138 modi5.n242 modi5.n241 4.137
R14139 modi5.n222 modi5.n220 3.764
R14140 modi5.n245 modi5.n238 3.764
R14141 modi5.n95 modi5.n92 3.764
R14142 modi5.n165 modi5.n163 3.764
R14143 modi5.n11 modi5.n6 3.464
R14144 modi5.n280 modi5.n279 3.388
R14145 modi5.n232 modi5.n231 3.388
R14146 modi5.n74 modi5.n71 3.388
R14147 modi5.n108 modi5.n107 3.388
R14148 modi5.n177 modi5.n176 3.388
R14149 modi5.n199 modi5.n198 3.388
R14150 modi5.n280 modi5.n278 3.011
R14151 modi5.n292 modi5.n289 3.011
R14152 modi5.n232 modi5.n230 3.011
R14153 modi5.n74 modi5.n73 3.011
R14154 modi5.n108 modi5.n105 3.011
R14155 modi5.n115 modi5.n113 3.011
R14156 modi5.n171 modi5.n170 3.011
R14157 modi5.n177 modi5.n175 3.011
R14158 modi5.n199 modi5.n197 3.011
R14159 modi5 modi5.n301 3.01
R14160 modi5.n222 modi5.n221 2.635
R14161 modi5.n253 modi5.n252 2.635
R14162 modi5.n245 modi5.n244 2.635
R14163 modi5.n95 modi5.n94 2.635
R14164 modi5.n89 modi5.n88 2.635
R14165 modi5.n158 modi5.n157 2.635
R14166 modi5.n165 modi5.n164 2.635
R14167 modi5.n64 modi5.n63 2.258
R14168 modi5.n187 modi5.n185 2.258
R14169 modi5.n301 modi5.n43 2.25
R14170 modi5.n78 modi5.n49 1.754
R14171 modi5.n251 modi5.n226 1.754
R14172 modi5.n78 modi5.n77 1.705
R14173 modi5.n153 modi5.n152 1.705
R14174 modi5.n147 modi5.n146 1.705
R14175 modi5.n142 modi5.n141 1.705
R14176 modi5.n136 modi5.n135 1.705
R14177 modi5.n119 modi5.n118 1.705
R14178 modi5.n99 modi5.n98 1.705
R14179 modi5.n84 modi5.n83 1.705
R14180 modi5.n299 modi5.n225 1.705
R14181 modi5.n298 modi5.n297 1.705
R14182 modi5.n268 modi5.n267 1.705
R14183 modi5.n251 modi5.n250 1.705
R14184 modi5.n212 modi5.n211 1.705
R14185 modi5.n158 modi5.n156 1.505
R14186 modi5.n235 modi5.n234 1.5
R14187 modi5.n250 modi5.n249 1.5
R14188 modi5.n297 modi5.n281 1.5
R14189 modi5.n296 modi5.n295 1.5
R14190 modi5.n257 modi5.n256 1.5
R14191 modi5.n286 modi5.n285 1.5
R14192 modi5.n266 modi5.n265 1.5
R14193 modi5.n224 modi5.n223 1.5
R14194 modi5.n132 modi5.n131 1.5
R14195 modi5.n126 modi5.n125 1.5
R14196 modi5.n117 modi5.n116 1.5
R14197 modi5.n110 modi5.n109 1.5
R14198 modi5.n97 modi5.n96 1.5
R14199 modi5.n38 modi5.n37 1.402
R14200 modi5.n13 modi5.n11 1.355
R14201 modi5.n300 modi5.n212 1.268
R14202 modi5.n14 modi5.n13 1.141
R14203 modi5.n26 modi5.n14 1.137
R14204 modi5.n3 modi5.n2 1.137
R14205 modi5.n20 modi5.n19 1.137
R14206 modi5.n39 modi5.n38 1.137
R14207 modi5.n31 modi5.n30 1.137
R14208 modi5.n23 modi5.n22 1.137
R14209 modi5.n25 modi5.n24 1.136
R14210 modi5.n41 modi5.n40 1.136
R14211 modi5.n211 modi5.n210 1.129
R14212 modi5.n115 modi5.n114 1.129
R14213 modi5.n49 modi5.n48 1.127
R14214 modi5.n201 modi5.n200 1.125
R14215 modi5.n76 modi5.n75 1.125
R14216 modi5.n274 modi5.n273 0.752
R14217 modi5.n240 modi5.n239 0.752
R14218 modi5.n300 modi5.n299 0.709
R14219 modi5.n47 modi5.n46 0.155
R14220 modi5.n209 modi5.n208 0.155
R14221 modi5.n73 modi5.n72 0.144
R14222 modi5.n197 modi5.n196 0.144
R14223 modi5.n63 modi5.n62 0.133
R14224 modi5.n185 modi5.n184 0.132
R14225 modi5.n218 modi5.n216 0.053
R14226 modi5.n54 modi5.n53 0.053
R14227 modi5.n69 modi5.n68 0.053
R14228 modi5.n59 modi5.n58 0.053
R14229 modi5.n172 modi5.n169 0.053
R14230 modi5.n182 modi5.n181 0.053
R14231 modi5.n192 modi5.n191 0.053
R14232 modi5.n84 modi5.n78 0.049
R14233 modi5.n99 modi5.n84 0.049
R14234 modi5.n119 modi5.n99 0.049
R14235 modi5.n136 modi5.n119 0.049
R14236 modi5.n142 modi5.n136 0.049
R14237 modi5.n147 modi5.n142 0.049
R14238 modi5.n153 modi5.n147 0.049
R14239 modi5.n212 modi5.n153 0.049
R14240 modi5.n299 modi5.n298 0.049
R14241 modi5.n298 modi5.n268 0.049
R14242 modi5.n268 modi5.n251 0.049
R14243 modi5.n11 modi5.n10 0.048
R14244 modi5.n125 modi5.n123 0.045
R14245 modi5.n159 modi5.n155 0.045
R14246 modi5.n295 modi5.n294 0.043
R14247 modi5.n265 modi5.n261 0.043
R14248 modi5.n191 modi5.n190 0.032
R14249 modi5.n206 modi5.n205 0.032
R14250 modi5.n224 modi5.n214 0.03
R14251 modi5.n236 modi5.n235 0.03
R14252 modi5.n70 modi5.n69 0.03
R14253 modi5.n68 modi5.n67 0.03
R14254 modi5.n181 modi5.n180 0.03
R14255 modi5.n58 modi5.n57 0.028
R14256 modi5.n193 modi5.n192 0.028
R14257 modi5.n195 modi5.n194 0.028
R14258 modi5.n55 modi5.n54 0.025
R14259 modi5.n60 modi5.n59 0.025
R14260 modi5.n131 modi5.n129 0.025
R14261 modi5.n94 modi5.n93 0.024
R14262 modi5.n175 modi5.n174 0.024
R14263 modi5.n285 modi5.n284 0.023
R14264 modi5.n183 modi5.n182 0.023
R14265 modi5.n223 modi5.n215 0.021
R14266 modi5.n219 modi5.n218 0.021
R14267 modi5.n247 modi5.n246 0.021
R14268 modi5.n91 modi5.n90 0.021
R14269 modi5.n166 modi5.n161 0.021
R14270 modi5.n169 modi5.n168 0.021
R14271 modi5.n19 modi5.n18 0.021
R14272 modi5.n270 modi5.n269 0.019
R14273 modi5.n281 modi5.n272 0.019
R14274 modi5.n248 modi5.n247 0.019
R14275 modi5.n229 modi5.n228 0.019
R14276 modi5.n234 modi5.n233 0.019
R14277 modi5.n75 modi5.n55 0.019
R14278 modi5.n103 modi5.n102 0.019
R14279 modi5.n104 modi5.n103 0.019
R14280 modi5.n168 modi5.n167 0.019
R14281 modi5.n173 modi5.n172 0.019
R14282 modi5.n179 modi5.n178 0.019
R14283 modi5.n200 modi5.n195 0.019
R14284 modi5.n210 modi5.n207 0.019
R14285 modi5.n48 modi5.n45 0.019
R14286 modi5.n2 modi5.n1 0.018
R14287 modi5.n19 modi5.n17 0.018
R14288 modi5.n22 modi5.n21 0.018
R14289 modi5.n30 modi5.n28 0.018
R14290 modi5.n281 modi5.n270 0.017
R14291 modi5.n234 modi5.n229 0.017
R14292 modi5.n75 modi5.n70 0.017
R14293 modi5.n66 modi5.n65 0.017
R14294 modi5.n109 modi5.n104 0.017
R14295 modi5.n116 modi5.n112 0.017
R14296 modi5.n178 modi5.n173 0.017
R14297 modi5.n189 modi5.n188 0.017
R14298 modi5.n200 modi5.n193 0.017
R14299 modi5.n98 modi5.n97 0.017
R14300 modi5.n297 modi5.n296 0.016
R14301 modi5.n52 modi5.n51 0.016
R14302 modi5.n80 modi5.n79 0.016
R14303 modi5.n86 modi5.n85 0.016
R14304 modi5.n146 modi5.n145 0.016
R14305 modi5.n151 modi5.n150 0.016
R14306 modi5.n203 modi5.n202 0.016
R14307 modi5.n10 modi5.n9 0.016
R14308 modi5.n8 modi5.n7 0.016
R14309 modi5.n35 modi5.n34 0.016
R14310 modi5.n37 modi5.n36 0.016
R14311 modi5.n223 modi5.n219 0.015
R14312 modi5.n256 modi5.n255 0.015
R14313 modi5.n249 modi5.n248 0.015
R14314 modi5.n287 modi5.n286 0.015
R14315 modi5.n258 modi5.n257 0.015
R14316 modi5.n96 modi5.n91 0.015
R14317 modi5.n160 modi5.n159 0.015
R14318 modi5.n167 modi5.n166 0.015
R14319 modi5.n117 modi5.n110 0.015
R14320 modi5.n132 modi5.n126 0.015
R14321 modi5.n138 modi5.n137 0.015
R14322 modi5.n296 modi5.n288 0.014
R14323 modi5.n266 modi5.n259 0.014
R14324 modi5.n202 modi5.n201 0.014
R14325 modi5 modi5.n42 0.014
R14326 modi5.n76 modi5.n52 0.013
R14327 modi5.n126 modi5.n121 0.013
R14328 modi5.n133 modi5.n132 0.013
R14329 modi5.n107 modi5.n106 0.012
R14330 modi5.n163 modi5.n162 0.012
R14331 modi5.n272 modi5.n271 0.012
R14332 modi5.n255 modi5.n254 0.012
R14333 modi5.n65 modi5.n60 0.012
R14334 modi5.n112 modi5.n111 0.012
R14335 modi5.n161 modi5.n160 0.012
R14336 modi5.n188 modi5.n183 0.012
R14337 modi5.n250 modi5.n237 0.011
R14338 modi5.n51 modi5.n50 0.011
R14339 modi5.n81 modi5.n80 0.011
R14340 modi5.n110 modi5.n101 0.011
R14341 modi5.n150 modi5.n149 0.011
R14342 modi5.n204 modi5.n203 0.011
R14343 modi5.n13 modi5.n12 0.011
R14344 modi5.n2 modi5.n0 0.011
R14345 modi5.n30 modi5.n29 0.011
R14346 modi5.n38 modi5.n33 0.011
R14347 modi5.n20 modi5.n16 0.011
R14348 modi5.n83 modi5.n82 0.01
R14349 modi5.n118 modi5.n117 0.01
R14350 modi5.n139 modi5.n138 0.01
R14351 modi5.n225 modi5.n224 0.009
R14352 modi5.n141 modi5.n140 0.009
R14353 modi5.n145 modi5.n144 0.009
R14354 modi5.n294 modi5.n293 0.008
R14355 modi5.n261 modi5.n260 0.008
R14356 modi5.n267 modi5.n266 0.008
R14357 modi5.n123 modi5.n122 0.008
R14358 modi5.n155 modi5.n154 0.008
R14359 modi5.n87 modi5.n86 0.008
R14360 modi5.n97 modi5.n87 0.008
R14361 modi5.n152 modi5.n151 0.008
R14362 modi5.n9 modi5.n8 0.008
R14363 modi5.n36 modi5.n35 0.008
R14364 modi5.n237 modi5.n236 0.007
R14365 modi5.n144 modi5.n143 0.007
R14366 modi5.n5 modi5.n4 0.007
R14367 modi5.n24 modi5.n20 0.007
R14368 modi5.n24 modi5.n23 0.007
R14369 modi5.n40 modi5.n32 0.007
R14370 modi5.n31 modi5.n27 0.007
R14371 modi5.n214 modi5.n213 0.006
R14372 modi5.n67 modi5.n66 0.006
R14373 modi5.n57 modi5.n56 0.006
R14374 modi5.n180 modi5.n179 0.006
R14375 modi5.n190 modi5.n189 0.006
R14376 modi5.n140 modi5.n139 0.006
R14377 modi5.n77 modi5.n76 0.005
R14378 modi5.n82 modi5.n81 0.005
R14379 modi5.n101 modi5.n100 0.005
R14380 modi5.n149 modi5.n148 0.005
R14381 modi5.n211 modi5.n204 0.005
R14382 modi5.n45 modi5.n44 0.004
R14383 modi5.n207 modi5.n206 0.004
R14384 modi5.n4 modi5.n3 0.004
R14385 modi5.n32 modi5.n31 0.004
R14386 modi5.n40 modi5.n39 0.004
R14387 modi5.n25 modi5.n15 0.004
R14388 modi5.n42 modi5.n41 0.003
R14389 modi5.n26 modi5.n25 0.002
R14390 modi5.n14 modi5.n5 0.002
R14391 modi5.n288 modi5.n287 0.002
R14392 modi5.n259 modi5.n258 0.002
R14393 modi5.n121 modi5.n120 0.002
R14394 modi5.n134 modi5.n133 0.002
R14395 modi5.n135 modi5.n134 0.002
R14396 modi5.n41 modi5.n26 0.002
R14397 a_n12857_2907.n95 a_n12857_2907.t4 730.681
R14398 a_n12857_2907.n95 a_n12857_2907.t3 395.834
R14399 a_n12857_2907.n41 a_n12857_2907.n40 13.176
R14400 a_n12857_2907.n96 a_n12857_2907.t0 11.721
R14401 a_n12857_2907.n96 a_n12857_2907.t2 10.994
R14402 a_n12857_2907.n150 a_n12857_2907.n34 9.3
R14403 a_n12857_2907.n150 a_n12857_2907.n141 9.3
R14404 a_n12857_2907.n150 a_n12857_2907.n135 9.3
R14405 a_n12857_2907.n150 a_n12857_2907.n49 9.3
R14406 a_n12857_2907.n150 a_n12857_2907.n54 9.3
R14407 a_n12857_2907.n150 a_n12857_2907.n123 9.3
R14408 a_n12857_2907.n150 a_n12857_2907.n149 8.469
R14409 a_n12857_2907.n150 a_n12857_2907.n113 8.469
R14410 a_n12857_2907.n150 a_n12857_2907.n118 8.125
R14411 a_n12857_2907.n150 a_n12857_2907.n29 8.124
R14412 a_n12857_2907.n150 a_n12857_2907.n110 8.097
R14413 a_n12857_2907.n150 a_n12857_2907.n146 8.096
R14414 a_n12857_2907.n150 a_n12857_2907.n126 8.016
R14415 a_n12857_2907.n150 a_n12857_2907.n39 8.016
R14416 a_n12857_2907.n150 a_n12857_2907.n130 7.964
R14417 a_n12857_2907.n150 a_n12857_2907.n44 7.964
R14418 a_n12857_2907.n125 a_n12857_2907.n124 6.4
R14419 a_n12857_2907.n109 a_n12857_2907.n55 6.4
R14420 a_n12857_2907.n144 a_n12857_2907.n143 6.023
R14421 a_n12857_2907.n37 a_n12857_2907.n36 6.023
R14422 a_n12857_2907.n135 a_n12857_2907.n134 6.023
R14423 a_n12857_2907.n43 a_n12857_2907.n42 6.023
R14424 a_n12857_2907.n129 a_n12857_2907.n128 6.023
R14425 a_n12857_2907.n148 a_n12857_2907.n147 5.647
R14426 a_n12857_2907.n49 a_n12857_2907.n46 5.647
R14427 a_n12857_2907.n116 a_n12857_2907.n115 5.647
R14428 a_n12857_2907.n112 a_n12857_2907.n111 5.647
R14429 a_n12857_2907.n132 a_n12857_2907.n131 5.457
R14430 a_n12857_2907.n27 a_n12857_2907.n26 5.27
R14431 a_n12857_2907.n48 a_n12857_2907.n47 5.08
R14432 a_n12857_2907.n34 a_n12857_2907.n33 4.517
R14433 a_n12857_2907.n123 a_n12857_2907.n120 4.517
R14434 a_n12857_2907.n63 a_n12857_2907.n62 4.5
R14435 a_n12857_2907.n2 a_n12857_2907.n1 4.5
R14436 a_n12857_2907.n31 a_n12857_2907.n30 4.314
R14437 a_n12857_2907.n140 a_n12857_2907.n139 4.141
R14438 a_n12857_2907.n51 a_n12857_2907.n50 4.141
R14439 a_n12857_2907.n137 a_n12857_2907.n136 3.944
R14440 a_n12857_2907.n122 a_n12857_2907.n121 3.937
R14441 a_n12857_2907.n53 a_n12857_2907.n52 3.567
R14442 a_n12857_2907.n109 a_n12857_2907.n108 3.033
R14443 a_n12857_2907.t1 a_n12857_2907.n150 2.9
R14444 a_n12857_2907.n141 a_n12857_2907.n140 2.258
R14445 a_n12857_2907.n54 a_n12857_2907.n51 2.258
R14446 a_n12857_2907.n33 a_n12857_2907.n32 1.882
R14447 a_n12857_2907.n120 a_n12857_2907.n119 1.882
R14448 a_n12857_2907.n98 a_n12857_2907.n97 1.672
R14449 a_n12857_2907.n54 a_n12857_2907.n53 1.505
R14450 a_n12857_2907.n82 a_n12857_2907.n102 1.5
R14451 a_n12857_2907.n64 a_n12857_2907.n66 1.5
R14452 a_n12857_2907.n63 a_n12857_2907.n61 1.5
R14453 a_n12857_2907.n21 a_n12857_2907.n24 1.5
R14454 a_n12857_2907.n12 a_n12857_2907.n11 1.5
R14455 a_n12857_2907.n108 a_n12857_2907.n80 1.5
R14456 a_n12857_2907.n97 a_n12857_2907.n96 1.221
R14457 a_n12857_2907.n28 a_n12857_2907.n27 1.129
R14458 a_n12857_2907.n26 a_n12857_2907.n25 1.129
R14459 a_n12857_2907.n141 a_n12857_2907.n137 1.129
R14460 a_n12857_2907.n139 a_n12857_2907.n138 1.129
R14461 a_n12857_2907.n101 a_n12857_2907.n100 0.853
R14462 a_n12857_2907.n149 a_n12857_2907.n148 0.752
R14463 a_n12857_2907.n46 a_n12857_2907.n45 0.752
R14464 a_n12857_2907.n49 a_n12857_2907.n48 0.752
R14465 a_n12857_2907.n123 a_n12857_2907.n122 0.752
R14466 a_n12857_2907.n115 a_n12857_2907.n114 0.752
R14467 a_n12857_2907.n117 a_n12857_2907.n116 0.752
R14468 a_n12857_2907.n113 a_n12857_2907.n112 0.752
R14469 a_n12857_2907.n89 a_n12857_2907.n88 0.716
R14470 a_n12857_2907.n97 a_n12857_2907.n95 0.637
R14471 a_n12857_2907.n130 a_n12857_2907.n129 0.536
R14472 a_n12857_2907.n44 a_n12857_2907.n43 0.536
R14473 a_n12857_2907.n126 a_n12857_2907.n125 0.476
R14474 a_n12857_2907.n39 a_n12857_2907.n38 0.475
R14475 a_n12857_2907.n110 a_n12857_2907.n109 0.382
R14476 a_n12857_2907.n146 a_n12857_2907.n145 0.382
R14477 a_n12857_2907.n145 a_n12857_2907.n144 0.376
R14478 a_n12857_2907.n143 a_n12857_2907.n142 0.376
R14479 a_n12857_2907.n34 a_n12857_2907.n31 0.376
R14480 a_n12857_2907.n38 a_n12857_2907.n37 0.376
R14481 a_n12857_2907.n36 a_n12857_2907.n35 0.376
R14482 a_n12857_2907.n135 a_n12857_2907.n132 0.376
R14483 a_n12857_2907.n134 a_n12857_2907.n133 0.376
R14484 a_n12857_2907.n42 a_n12857_2907.n41 0.376
R14485 a_n12857_2907.n128 a_n12857_2907.n127 0.376
R14486 a_n12857_2907.n118 a_n12857_2907.n117 0.35
R14487 a_n12857_2907.n29 a_n12857_2907.n28 0.349
R14488 a_n12857_2907.n2 a_n12857_2907.n0 0.066
R14489 a_n12857_2907.n87 a_n12857_2907.n86 0.047
R14490 a_n12857_2907.n72 a_n12857_2907.n71 0.043
R14491 a_n12857_2907.n68 a_n12857_2907.n67 0.043
R14492 a_n12857_2907.n64 a_n12857_2907.n63 0.041
R14493 a_n12857_2907.n79 a_n12857_2907.n78 0.035
R14494 a_n12857_2907.n107 a_n12857_2907.n106 0.035
R14495 a_n12857_2907.n19 a_n12857_2907.n18 0.034
R14496 a_n12857_2907.n23 a_n12857_2907.n22 0.034
R14497 a_n12857_2907.n8 a_n12857_2907.n7 0.034
R14498 a_n12857_2907.n77 a_n12857_2907.n76 0.034
R14499 a_n12857_2907.n105 a_n12857_2907.n104 0.034
R14500 a_n12857_2907.n12 a_n12857_2907.n6 0.032
R14501 a_n12857_2907.n108 a_n12857_2907.n70 0.032
R14502 a_n12857_2907.n99 a_n12857_2907.n98 0.031
R14503 a_n12857_2907.n9 a_n12857_2907.n8 0.03
R14504 a_n12857_2907.n75 a_n12857_2907.n74 0.03
R14505 a_n12857_2907.n101 a_n12857_2907.n94 0.03
R14506 a_n12857_2907.n81 a_n12857_2907.n87 0.03
R14507 a_n12857_2907.n11 a_n12857_2907.n10 0.028
R14508 a_n12857_2907.n60 a_n12857_2907.n58 0.028
R14509 a_n12857_2907.n73 a_n12857_2907.n72 0.028
R14510 a_n12857_2907.n91 a_n12857_2907.n90 0.028
R14511 a_n12857_2907.n13 a_n12857_2907.n12 0.028
R14512 a_n12857_2907.n57 a_n12857_2907.n56 0.028
R14513 a_n12857_2907.n69 a_n12857_2907.n68 0.028
R14514 a_n12857_2907.n103 a_n12857_2907.n82 0.028
R14515 a_n12857_2907.n85 a_n12857_2907.n83 0.028
R14516 a_n12857_2907.n17 a_n12857_2907.n15 0.026
R14517 a_n12857_2907.n66 a_n12857_2907.n65 0.026
R14518 a_n12857_2907.n93 a_n12857_2907.n92 0.026
R14519 a_n12857_2907.n4 a_n12857_2907.n3 0.026
R14520 a_n12857_2907.n90 a_n12857_2907.n89 0.024
R14521 a_n12857_2907.n18 a_n12857_2907.n17 0.024
R14522 a_n12857_2907.n6 a_n12857_2907.n5 0.024
R14523 a_n12857_2907.n15 a_n12857_2907.n16 0.022
R14524 a_n12857_2907.n5 a_n12857_2907.n4 0.022
R14525 a_n12857_2907.n3 a_n12857_2907.n2 0.022
R14526 a_n12857_2907.n20 a_n12857_2907.n19 0.02
R14527 a_n12857_2907.n10 a_n12857_2907.n9 0.02
R14528 a_n12857_2907.n94 a_n12857_2907.n93 0.02
R14529 a_n12857_2907.n14 a_n12857_2907.n13 0.02
R14530 a_n12857_2907.n100 a_n12857_2907.n99 0.019
R14531 a_n12857_2907.n82 a_n12857_2907.n81 0.018
R14532 a_n12857_2907.n102 a_n12857_2907.n101 0.018
R14533 a_n12857_2907.n70 a_n12857_2907.n69 0.018
R14534 a_n12857_2907.n24 a_n12857_2907.n23 0.017
R14535 a_n12857_2907.n74 a_n12857_2907.n73 0.017
R14536 a_n12857_2907.n58 a_n12857_2907.n59 0.015
R14537 a_n12857_2907.n61 a_n12857_2907.n60 0.015
R14538 a_n12857_2907.n56 a_n12857_2907.n0 0.015
R14539 a_n12857_2907.n63 a_n12857_2907.n57 0.015
R14540 a_n12857_2907.n80 a_n12857_2907.n79 0.013
R14541 a_n12857_2907.n78 a_n12857_2907.n77 0.013
R14542 a_n12857_2907.n108 a_n12857_2907.n107 0.013
R14543 a_n12857_2907.n106 a_n12857_2907.n105 0.013
R14544 a_n12857_2907.n92 a_n12857_2907.n91 0.007
R14545 a_n12857_2907.n86 a_n12857_2907.n85 0.007
R14546 a_n12857_2907.n21 a_n12857_2907.n20 1.424
R14547 a_n12857_2907.n67 a_n12857_2907.n64 0.005
R14548 a_n12857_2907.n80 a_n12857_2907.n75 0.003
R14549 a_n12857_2907.n104 a_n12857_2907.n103 0.003
R14550 a_n12857_2907.n83 a_n12857_2907.n84 0.003
R14551 a_n12857_2907.n14 a_n12857_2907.n21 0.47
R14552 a_n24474_2912.n95 a_n24474_2912.t4 730.681
R14553 a_n24474_2912.n95 a_n24474_2912.t3 395.834
R14554 a_n24474_2912.n41 a_n24474_2912.n40 13.176
R14555 a_n24474_2912.n96 a_n24474_2912.t0 11.722
R14556 a_n24474_2912.n96 a_n24474_2912.t1 10.994
R14557 a_n24474_2912.n150 a_n24474_2912.n34 9.3
R14558 a_n24474_2912.n150 a_n24474_2912.n141 9.3
R14559 a_n24474_2912.n150 a_n24474_2912.n135 9.3
R14560 a_n24474_2912.n150 a_n24474_2912.n49 9.3
R14561 a_n24474_2912.n150 a_n24474_2912.n54 9.3
R14562 a_n24474_2912.n150 a_n24474_2912.n123 9.3
R14563 a_n24474_2912.n150 a_n24474_2912.n149 8.469
R14564 a_n24474_2912.n150 a_n24474_2912.n113 8.469
R14565 a_n24474_2912.n150 a_n24474_2912.n118 8.125
R14566 a_n24474_2912.n150 a_n24474_2912.n29 8.124
R14567 a_n24474_2912.n150 a_n24474_2912.n110 8.097
R14568 a_n24474_2912.n150 a_n24474_2912.n146 8.096
R14569 a_n24474_2912.n150 a_n24474_2912.n126 8.016
R14570 a_n24474_2912.n150 a_n24474_2912.n39 8.016
R14571 a_n24474_2912.n150 a_n24474_2912.n130 7.964
R14572 a_n24474_2912.n150 a_n24474_2912.n44 7.964
R14573 a_n24474_2912.n125 a_n24474_2912.n124 6.4
R14574 a_n24474_2912.n109 a_n24474_2912.n55 6.4
R14575 a_n24474_2912.n144 a_n24474_2912.n143 6.023
R14576 a_n24474_2912.n37 a_n24474_2912.n36 6.023
R14577 a_n24474_2912.n135 a_n24474_2912.n134 6.023
R14578 a_n24474_2912.n43 a_n24474_2912.n42 6.023
R14579 a_n24474_2912.n129 a_n24474_2912.n128 6.023
R14580 a_n24474_2912.n148 a_n24474_2912.n147 5.647
R14581 a_n24474_2912.n49 a_n24474_2912.n46 5.647
R14582 a_n24474_2912.n116 a_n24474_2912.n115 5.647
R14583 a_n24474_2912.n112 a_n24474_2912.n111 5.647
R14584 a_n24474_2912.n132 a_n24474_2912.n131 5.457
R14585 a_n24474_2912.n27 a_n24474_2912.n26 5.27
R14586 a_n24474_2912.n48 a_n24474_2912.n47 5.08
R14587 a_n24474_2912.n34 a_n24474_2912.n33 4.517
R14588 a_n24474_2912.n123 a_n24474_2912.n120 4.517
R14589 a_n24474_2912.n63 a_n24474_2912.n62 4.5
R14590 a_n24474_2912.n2 a_n24474_2912.n1 4.5
R14591 a_n24474_2912.n31 a_n24474_2912.n30 4.314
R14592 a_n24474_2912.n140 a_n24474_2912.n139 4.141
R14593 a_n24474_2912.n51 a_n24474_2912.n50 4.141
R14594 a_n24474_2912.n137 a_n24474_2912.n136 3.944
R14595 a_n24474_2912.n122 a_n24474_2912.n121 3.937
R14596 a_n24474_2912.n53 a_n24474_2912.n52 3.567
R14597 a_n24474_2912.n109 a_n24474_2912.n108 3.033
R14598 a_n24474_2912.t2 a_n24474_2912.n150 2.9
R14599 a_n24474_2912.n141 a_n24474_2912.n140 2.258
R14600 a_n24474_2912.n54 a_n24474_2912.n51 2.258
R14601 a_n24474_2912.n33 a_n24474_2912.n32 1.882
R14602 a_n24474_2912.n120 a_n24474_2912.n119 1.882
R14603 a_n24474_2912.n98 a_n24474_2912.n97 1.672
R14604 a_n24474_2912.n54 a_n24474_2912.n53 1.505
R14605 a_n24474_2912.n82 a_n24474_2912.n102 1.5
R14606 a_n24474_2912.n64 a_n24474_2912.n66 1.5
R14607 a_n24474_2912.n63 a_n24474_2912.n61 1.5
R14608 a_n24474_2912.n21 a_n24474_2912.n24 1.5
R14609 a_n24474_2912.n12 a_n24474_2912.n11 1.5
R14610 a_n24474_2912.n108 a_n24474_2912.n80 1.5
R14611 a_n24474_2912.n97 a_n24474_2912.n96 1.222
R14612 a_n24474_2912.n28 a_n24474_2912.n27 1.129
R14613 a_n24474_2912.n26 a_n24474_2912.n25 1.129
R14614 a_n24474_2912.n141 a_n24474_2912.n137 1.129
R14615 a_n24474_2912.n139 a_n24474_2912.n138 1.129
R14616 a_n24474_2912.n101 a_n24474_2912.n100 0.853
R14617 a_n24474_2912.n149 a_n24474_2912.n148 0.752
R14618 a_n24474_2912.n46 a_n24474_2912.n45 0.752
R14619 a_n24474_2912.n49 a_n24474_2912.n48 0.752
R14620 a_n24474_2912.n123 a_n24474_2912.n122 0.752
R14621 a_n24474_2912.n115 a_n24474_2912.n114 0.752
R14622 a_n24474_2912.n117 a_n24474_2912.n116 0.752
R14623 a_n24474_2912.n113 a_n24474_2912.n112 0.752
R14624 a_n24474_2912.n89 a_n24474_2912.n88 0.716
R14625 a_n24474_2912.n97 a_n24474_2912.n95 0.637
R14626 a_n24474_2912.n130 a_n24474_2912.n129 0.536
R14627 a_n24474_2912.n44 a_n24474_2912.n43 0.536
R14628 a_n24474_2912.n126 a_n24474_2912.n125 0.476
R14629 a_n24474_2912.n39 a_n24474_2912.n38 0.475
R14630 a_n24474_2912.n110 a_n24474_2912.n109 0.382
R14631 a_n24474_2912.n146 a_n24474_2912.n145 0.382
R14632 a_n24474_2912.n145 a_n24474_2912.n144 0.376
R14633 a_n24474_2912.n143 a_n24474_2912.n142 0.376
R14634 a_n24474_2912.n34 a_n24474_2912.n31 0.376
R14635 a_n24474_2912.n38 a_n24474_2912.n37 0.376
R14636 a_n24474_2912.n36 a_n24474_2912.n35 0.376
R14637 a_n24474_2912.n135 a_n24474_2912.n132 0.376
R14638 a_n24474_2912.n134 a_n24474_2912.n133 0.376
R14639 a_n24474_2912.n42 a_n24474_2912.n41 0.376
R14640 a_n24474_2912.n128 a_n24474_2912.n127 0.376
R14641 a_n24474_2912.n118 a_n24474_2912.n117 0.35
R14642 a_n24474_2912.n29 a_n24474_2912.n28 0.349
R14643 a_n24474_2912.n2 a_n24474_2912.n0 0.066
R14644 a_n24474_2912.n87 a_n24474_2912.n86 0.047
R14645 a_n24474_2912.n72 a_n24474_2912.n71 0.043
R14646 a_n24474_2912.n68 a_n24474_2912.n67 0.043
R14647 a_n24474_2912.n64 a_n24474_2912.n63 0.041
R14648 a_n24474_2912.n79 a_n24474_2912.n78 0.035
R14649 a_n24474_2912.n107 a_n24474_2912.n106 0.035
R14650 a_n24474_2912.n19 a_n24474_2912.n18 0.034
R14651 a_n24474_2912.n23 a_n24474_2912.n22 0.034
R14652 a_n24474_2912.n8 a_n24474_2912.n7 0.034
R14653 a_n24474_2912.n77 a_n24474_2912.n76 0.034
R14654 a_n24474_2912.n105 a_n24474_2912.n104 0.034
R14655 a_n24474_2912.n12 a_n24474_2912.n6 0.032
R14656 a_n24474_2912.n108 a_n24474_2912.n70 0.032
R14657 a_n24474_2912.n99 a_n24474_2912.n98 0.031
R14658 a_n24474_2912.n9 a_n24474_2912.n8 0.03
R14659 a_n24474_2912.n75 a_n24474_2912.n74 0.03
R14660 a_n24474_2912.n101 a_n24474_2912.n94 0.03
R14661 a_n24474_2912.n81 a_n24474_2912.n87 0.03
R14662 a_n24474_2912.n11 a_n24474_2912.n10 0.028
R14663 a_n24474_2912.n60 a_n24474_2912.n58 0.028
R14664 a_n24474_2912.n73 a_n24474_2912.n72 0.028
R14665 a_n24474_2912.n91 a_n24474_2912.n90 0.028
R14666 a_n24474_2912.n13 a_n24474_2912.n12 0.028
R14667 a_n24474_2912.n57 a_n24474_2912.n56 0.028
R14668 a_n24474_2912.n69 a_n24474_2912.n68 0.028
R14669 a_n24474_2912.n103 a_n24474_2912.n82 0.028
R14670 a_n24474_2912.n85 a_n24474_2912.n83 0.028
R14671 a_n24474_2912.n17 a_n24474_2912.n15 0.026
R14672 a_n24474_2912.n66 a_n24474_2912.n65 0.026
R14673 a_n24474_2912.n93 a_n24474_2912.n92 0.026
R14674 a_n24474_2912.n4 a_n24474_2912.n3 0.026
R14675 a_n24474_2912.n90 a_n24474_2912.n89 0.024
R14676 a_n24474_2912.n18 a_n24474_2912.n17 0.024
R14677 a_n24474_2912.n6 a_n24474_2912.n5 0.024
R14678 a_n24474_2912.n15 a_n24474_2912.n16 0.022
R14679 a_n24474_2912.n5 a_n24474_2912.n4 0.022
R14680 a_n24474_2912.n3 a_n24474_2912.n2 0.022
R14681 a_n24474_2912.n20 a_n24474_2912.n19 0.02
R14682 a_n24474_2912.n10 a_n24474_2912.n9 0.02
R14683 a_n24474_2912.n94 a_n24474_2912.n93 0.02
R14684 a_n24474_2912.n14 a_n24474_2912.n13 0.02
R14685 a_n24474_2912.n100 a_n24474_2912.n99 0.019
R14686 a_n24474_2912.n82 a_n24474_2912.n81 0.018
R14687 a_n24474_2912.n102 a_n24474_2912.n101 0.018
R14688 a_n24474_2912.n70 a_n24474_2912.n69 0.018
R14689 a_n24474_2912.n24 a_n24474_2912.n23 0.017
R14690 a_n24474_2912.n74 a_n24474_2912.n73 0.017
R14691 a_n24474_2912.n58 a_n24474_2912.n59 0.015
R14692 a_n24474_2912.n61 a_n24474_2912.n60 0.015
R14693 a_n24474_2912.n56 a_n24474_2912.n0 0.015
R14694 a_n24474_2912.n63 a_n24474_2912.n57 0.015
R14695 a_n24474_2912.n80 a_n24474_2912.n79 0.013
R14696 a_n24474_2912.n78 a_n24474_2912.n77 0.013
R14697 a_n24474_2912.n108 a_n24474_2912.n107 0.013
R14698 a_n24474_2912.n106 a_n24474_2912.n105 0.013
R14699 a_n24474_2912.n92 a_n24474_2912.n91 0.007
R14700 a_n24474_2912.n86 a_n24474_2912.n85 0.007
R14701 a_n24474_2912.n21 a_n24474_2912.n20 1.424
R14702 a_n24474_2912.n67 a_n24474_2912.n64 0.005
R14703 a_n24474_2912.n80 a_n24474_2912.n75 0.003
R14704 a_n24474_2912.n104 a_n24474_2912.n103 0.003
R14705 a_n24474_2912.n83 a_n24474_2912.n84 0.003
R14706 a_n24474_2912.n14 a_n24474_2912.n21 0.47
R14707 a_n24497_6006.n13 a_n24497_6006.t2 732.458
R14708 a_n24497_6006.n13 a_n24497_6006.t3 397.578
R14709 a_n24497_6006.n51 a_n24497_6006.n50 92.5
R14710 a_n24497_6006.n9 a_n24497_6006.n8 92.5
R14711 a_n24497_6006.n50 a_n24497_6006.t1 70.344
R14712 a_n24497_6006.n45 a_n24497_6006.n44 31.034
R14713 a_n24497_6006.n24 a_n24497_6006.n23 31.034
R14714 a_n24497_6006.n27 a_n24497_6006.n28 9.3
R14715 a_n24497_6006.n38 a_n24497_6006.n39 9.3
R14716 a_n24497_6006.n46 a_n24497_6006.n45 9.3
R14717 a_n24497_6006.n25 a_n24497_6006.n24 9.3
R14718 a_n24497_6006.n105 a_n24497_6006.n98 9.154
R14719 a_n24497_6006.n105 a_n24497_6006.n4 9.143
R14720 a_n24497_6006.n105 a_n24497_6006.n3 9.143
R14721 a_n24497_6006.n105 a_n24497_6006.n78 9.132
R14722 a_n24497_6006.n105 a_n24497_6006.n62 9.132
R14723 a_n24497_6006.n105 a_n24497_6006.n102 8.885
R14724 a_n24497_6006.n105 a_n24497_6006.n82 8.885
R14725 a_n24497_6006.n105 a_n24497_6006.n86 8.875
R14726 a_n24497_6006.n105 a_n24497_6006.n56 8.875
R14727 a_n24497_6006.n105 a_n24497_6006.n104 8.864
R14728 a_n24497_6006.n105 a_n24497_6006.n88 8.864
R14729 a_n24497_6006.n52 a_n24497_6006.n51 8.282
R14730 a_n24497_6006.n10 a_n24497_6006.n9 8.282
R14731 a_n24497_6006.t0 a_n24497_6006.n105 7.141
R14732 a_n24497_6006.n46 a_n24497_6006.n42 5.647
R14733 a_n24497_6006.n25 a_n24497_6006.n21 5.647
R14734 a_n24497_6006.n1 a_n24497_6006.n11 4.65
R14735 a_n24497_6006.n16 a_n24497_6006.n15 4.566
R14736 a_n24497_6006.n98 a_n24497_6006.n90 4.517
R14737 a_n24497_6006.n0 a_n24497_6006.n10 4.5
R14738 a_n24497_6006.n1 a_n24497_6006.n7 4.5
R14739 a_n24497_6006.n6 a_n24497_6006.n52 4.5
R14740 a_n24497_6006.n40 a_n24497_6006.n48 4.5
R14741 a_n24497_6006.n12 a_n24497_6006.n37 4.5
R14742 a_n24497_6006.n17 a_n24497_6006.n32 4.5
R14743 a_n24497_6006.n15 a_n24497_6006.n14 4.481
R14744 a_n24497_6006.n100 a_n24497_6006.n99 4.141
R14745 a_n24497_6006.n98 a_n24497_6006.n89 4.141
R14746 a_n24497_6006.n80 a_n24497_6006.n79 4.141
R14747 a_n24497_6006.n44 a_n24497_6006.n43 4.137
R14748 a_n24497_6006.n23 a_n24497_6006.n22 4.137
R14749 a_n24497_6006.n37 a_n24497_6006.n35 3.764
R14750 a_n24497_6006.n26 a_n24497_6006.n19 3.764
R14751 a_n24497_6006.n58 a_n24497_6006.n57 3.764
R14752 a_n24497_6006.n3 a_n24497_6006.n69 3.764
R14753 a_n24497_6006.n62 a_n24497_6006.n61 3.736
R14754 a_n24497_6006.n48 a_n24497_6006.n47 3.388
R14755 a_n24497_6006.n32 a_n24497_6006.n31 3.388
R14756 a_n24497_6006.n54 a_n24497_6006.n53 3.388
R14757 a_n24497_6006.n4 a_n24497_6006.n67 3.388
R14758 a_n24497_6006.n76 a_n24497_6006.n75 3.388
R14759 a_n24497_6006.n84 a_n24497_6006.n83 3.388
R14760 a_n24497_6006.n78 a_n24497_6006.n74 3.36
R14761 a_n24497_6006.n48 a_n24497_6006.n46 3.011
R14762 a_n24497_6006.n52 a_n24497_6006.n49 3.011
R14763 a_n24497_6006.n32 a_n24497_6006.n30 3.011
R14764 a_n24497_6006.n55 a_n24497_6006.n54 3.011
R14765 a_n24497_6006.n67 a_n24497_6006.n66 3.011
R14766 a_n24497_6006.n65 a_n24497_6006.n64 3.011
R14767 a_n24497_6006.n74 a_n24497_6006.n73 3.011
R14768 a_n24497_6006.n77 a_n24497_6006.n76 3.011
R14769 a_n24497_6006.n85 a_n24497_6006.n84 3.011
R14770 a_n24497_6006.n91 a_n24497_6006.n14 2.921
R14771 a_n24497_6006.n37 a_n24497_6006.n36 2.635
R14772 a_n24497_6006.n26 a_n24497_6006.n25 2.635
R14773 a_n24497_6006.n59 a_n24497_6006.n58 2.635
R14774 a_n24497_6006.n61 a_n24497_6006.n60 2.635
R14775 a_n24497_6006.n72 a_n24497_6006.n71 2.635
R14776 a_n24497_6006.n69 a_n24497_6006.n68 2.635
R14777 a_n24497_6006.n15 a_n24497_6006.n13 2.349
R14778 a_n24497_6006.n101 a_n24497_6006.n100 2.258
R14779 a_n24497_6006.n81 a_n24497_6006.n80 2.258
R14780 a_n24497_6006.n5 a_n24497_6006.n96 1.633
R14781 a_n24497_6006.n2 a_n24497_6006.n95 1.619
R14782 a_n24497_6006.n92 a_n24497_6006.n93 1.588
R14783 a_n24497_6006.n5 a_n24497_6006.n106 1.587
R14784 a_n24497_6006.n71 a_n24497_6006.n70 1.505
R14785 a_n24497_6006.n12 a_n24497_6006.n34 1.5
R14786 a_n24497_6006.n64 a_n24497_6006.n63 1.129
R14787 a_n24497_6006.n42 a_n24497_6006.n41 0.752
R14788 a_n24497_6006.n21 a_n24497_6006.n20 0.752
R14789 a_n24497_6006.n104 a_n24497_6006.n103 0.155
R14790 a_n24497_6006.n88 a_n24497_6006.n87 0.155
R14791 a_n24497_6006.n56 a_n24497_6006.n55 0.144
R14792 a_n24497_6006.n86 a_n24497_6006.n85 0.144
R14793 a_n24497_6006.n102 a_n24497_6006.n101 0.132
R14794 a_n24497_6006.n82 a_n24497_6006.n81 0.132
R14795 a_n24497_6006.n91 a_n24497_6006.n92 0.125
R14796 a_n24497_6006.n106 a_n24497_6006.n107 0.037
R14797 a_n24497_6006.n96 a_n24497_6006.n97 0.034
R14798 a_n24497_6006.n40 a_n24497_6006.n38 0.094
R14799 a_n24497_6006.n34 a_n24497_6006.n33 0.293
R14800 a_n24497_6006.n34 a_n24497_6006.n18 0.877
R14801 a_n24497_6006.n93 a_n24497_6006.n94 0.024
R14802 a_n24497_6006.n62 a_n24497_6006.n59 0.024
R14803 a_n24497_6006.n78 a_n24497_6006.n77 0.024
R14804 a_n24497_6006.n98 a_n24497_6006.n91 4.672
R14805 a_n24497_6006.n18 a_n24497_6006.n16 0.019
R14806 a_n24497_6006.n18 a_n24497_6006.n17 2.433
R14807 a_n24497_6006.n6 a_n24497_6006.n40 0.044
R14808 a_n24497_6006.n17 a_n24497_6006.n27 0.032
R14809 a_n24497_6006.n38 a_n24497_6006.n12 0.031
R14810 a_n24497_6006.n17 a_n24497_6006.n29 0.017
R14811 a_n24497_6006.n27 a_n24497_6006.n26 4.595
R14812 a_n24497_6006.n4 a_n24497_6006.n65 2.257
R14813 a_n24497_6006.n3 a_n24497_6006.n72 2.257
R14814 a_n24497_6006.n2 a_n24497_6006.n5 0.256
R14815 a_n24497_6006.n92 a_n24497_6006.n2 0.124
R14816 a_n24497_6006.n6 a_n24497_6006.n1 0.07
R14817 a_n24497_6006.n1 a_n24497_6006.n0 0.053
R14818 a_n7023_6002.n13 a_n7023_6002.t3 732.458
R14819 a_n7023_6002.n13 a_n7023_6002.t2 397.578
R14820 a_n7023_6002.n51 a_n7023_6002.n50 92.5
R14821 a_n7023_6002.n9 a_n7023_6002.n8 92.5
R14822 a_n7023_6002.n50 a_n7023_6002.t1 70.344
R14823 a_n7023_6002.n45 a_n7023_6002.n44 31.034
R14824 a_n7023_6002.n24 a_n7023_6002.n23 31.034
R14825 a_n7023_6002.n27 a_n7023_6002.n28 9.3
R14826 a_n7023_6002.n38 a_n7023_6002.n39 9.3
R14827 a_n7023_6002.n46 a_n7023_6002.n45 9.3
R14828 a_n7023_6002.n25 a_n7023_6002.n24 9.3
R14829 a_n7023_6002.n105 a_n7023_6002.n98 9.154
R14830 a_n7023_6002.n105 a_n7023_6002.n4 9.143
R14831 a_n7023_6002.n105 a_n7023_6002.n3 9.143
R14832 a_n7023_6002.n105 a_n7023_6002.n78 9.132
R14833 a_n7023_6002.n105 a_n7023_6002.n62 9.132
R14834 a_n7023_6002.n105 a_n7023_6002.n102 8.885
R14835 a_n7023_6002.n105 a_n7023_6002.n82 8.885
R14836 a_n7023_6002.n105 a_n7023_6002.n86 8.875
R14837 a_n7023_6002.n105 a_n7023_6002.n56 8.875
R14838 a_n7023_6002.n105 a_n7023_6002.n104 8.864
R14839 a_n7023_6002.n105 a_n7023_6002.n88 8.864
R14840 a_n7023_6002.n52 a_n7023_6002.n51 8.282
R14841 a_n7023_6002.n10 a_n7023_6002.n9 8.282
R14842 a_n7023_6002.t0 a_n7023_6002.n105 7.141
R14843 a_n7023_6002.n46 a_n7023_6002.n42 5.647
R14844 a_n7023_6002.n25 a_n7023_6002.n21 5.647
R14845 a_n7023_6002.n1 a_n7023_6002.n11 4.65
R14846 a_n7023_6002.n16 a_n7023_6002.n15 4.566
R14847 a_n7023_6002.n98 a_n7023_6002.n90 4.517
R14848 a_n7023_6002.n0 a_n7023_6002.n10 4.5
R14849 a_n7023_6002.n1 a_n7023_6002.n7 4.5
R14850 a_n7023_6002.n6 a_n7023_6002.n52 4.5
R14851 a_n7023_6002.n40 a_n7023_6002.n48 4.5
R14852 a_n7023_6002.n12 a_n7023_6002.n37 4.5
R14853 a_n7023_6002.n17 a_n7023_6002.n32 4.5
R14854 a_n7023_6002.n15 a_n7023_6002.n14 4.482
R14855 a_n7023_6002.n100 a_n7023_6002.n99 4.141
R14856 a_n7023_6002.n98 a_n7023_6002.n89 4.141
R14857 a_n7023_6002.n80 a_n7023_6002.n79 4.141
R14858 a_n7023_6002.n44 a_n7023_6002.n43 4.137
R14859 a_n7023_6002.n23 a_n7023_6002.n22 4.137
R14860 a_n7023_6002.n37 a_n7023_6002.n35 3.764
R14861 a_n7023_6002.n26 a_n7023_6002.n19 3.764
R14862 a_n7023_6002.n58 a_n7023_6002.n57 3.764
R14863 a_n7023_6002.n3 a_n7023_6002.n69 3.764
R14864 a_n7023_6002.n62 a_n7023_6002.n61 3.736
R14865 a_n7023_6002.n48 a_n7023_6002.n47 3.388
R14866 a_n7023_6002.n32 a_n7023_6002.n31 3.388
R14867 a_n7023_6002.n54 a_n7023_6002.n53 3.388
R14868 a_n7023_6002.n4 a_n7023_6002.n67 3.388
R14869 a_n7023_6002.n76 a_n7023_6002.n75 3.388
R14870 a_n7023_6002.n84 a_n7023_6002.n83 3.388
R14871 a_n7023_6002.n78 a_n7023_6002.n74 3.36
R14872 a_n7023_6002.n48 a_n7023_6002.n46 3.011
R14873 a_n7023_6002.n52 a_n7023_6002.n49 3.011
R14874 a_n7023_6002.n32 a_n7023_6002.n30 3.011
R14875 a_n7023_6002.n55 a_n7023_6002.n54 3.011
R14876 a_n7023_6002.n67 a_n7023_6002.n66 3.011
R14877 a_n7023_6002.n65 a_n7023_6002.n64 3.011
R14878 a_n7023_6002.n74 a_n7023_6002.n73 3.011
R14879 a_n7023_6002.n77 a_n7023_6002.n76 3.011
R14880 a_n7023_6002.n85 a_n7023_6002.n84 3.011
R14881 a_n7023_6002.n91 a_n7023_6002.n14 2.921
R14882 a_n7023_6002.n37 a_n7023_6002.n36 2.635
R14883 a_n7023_6002.n26 a_n7023_6002.n25 2.635
R14884 a_n7023_6002.n59 a_n7023_6002.n58 2.635
R14885 a_n7023_6002.n61 a_n7023_6002.n60 2.635
R14886 a_n7023_6002.n72 a_n7023_6002.n71 2.635
R14887 a_n7023_6002.n69 a_n7023_6002.n68 2.635
R14888 a_n7023_6002.n15 a_n7023_6002.n13 2.354
R14889 a_n7023_6002.n101 a_n7023_6002.n100 2.258
R14890 a_n7023_6002.n81 a_n7023_6002.n80 2.258
R14891 a_n7023_6002.n5 a_n7023_6002.n96 1.633
R14892 a_n7023_6002.n2 a_n7023_6002.n95 1.619
R14893 a_n7023_6002.n92 a_n7023_6002.n93 1.588
R14894 a_n7023_6002.n5 a_n7023_6002.n106 1.587
R14895 a_n7023_6002.n71 a_n7023_6002.n70 1.505
R14896 a_n7023_6002.n12 a_n7023_6002.n34 1.5
R14897 a_n7023_6002.n64 a_n7023_6002.n63 1.129
R14898 a_n7023_6002.n42 a_n7023_6002.n41 0.752
R14899 a_n7023_6002.n21 a_n7023_6002.n20 0.752
R14900 a_n7023_6002.n104 a_n7023_6002.n103 0.155
R14901 a_n7023_6002.n88 a_n7023_6002.n87 0.155
R14902 a_n7023_6002.n56 a_n7023_6002.n55 0.144
R14903 a_n7023_6002.n86 a_n7023_6002.n85 0.144
R14904 a_n7023_6002.n102 a_n7023_6002.n101 0.132
R14905 a_n7023_6002.n82 a_n7023_6002.n81 0.132
R14906 a_n7023_6002.n91 a_n7023_6002.n92 0.125
R14907 a_n7023_6002.n106 a_n7023_6002.n107 0.037
R14908 a_n7023_6002.n96 a_n7023_6002.n97 0.034
R14909 a_n7023_6002.n40 a_n7023_6002.n38 0.094
R14910 a_n7023_6002.n34 a_n7023_6002.n33 0.293
R14911 a_n7023_6002.n34 a_n7023_6002.n18 0.877
R14912 a_n7023_6002.n93 a_n7023_6002.n94 0.024
R14913 a_n7023_6002.n62 a_n7023_6002.n59 0.024
R14914 a_n7023_6002.n78 a_n7023_6002.n77 0.024
R14915 a_n7023_6002.n98 a_n7023_6002.n91 4.672
R14916 a_n7023_6002.n18 a_n7023_6002.n16 0.019
R14917 a_n7023_6002.n18 a_n7023_6002.n17 2.433
R14918 a_n7023_6002.n6 a_n7023_6002.n40 0.044
R14919 a_n7023_6002.n17 a_n7023_6002.n27 0.032
R14920 a_n7023_6002.n38 a_n7023_6002.n12 0.031
R14921 a_n7023_6002.n17 a_n7023_6002.n29 0.017
R14922 a_n7023_6002.n27 a_n7023_6002.n26 4.595
R14923 a_n7023_6002.n4 a_n7023_6002.n65 2.257
R14924 a_n7023_6002.n3 a_n7023_6002.n72 2.257
R14925 a_n7023_6002.n2 a_n7023_6002.n5 0.256
R14926 a_n7023_6002.n92 a_n7023_6002.n2 0.124
R14927 a_n7023_6002.n6 a_n7023_6002.n1 0.07
R14928 a_n7023_6002.n1 a_n7023_6002.n0 0.053
R14929 fout3.n536 fout3.t5 1038.95
R14930 fout3.n8 fout3.t6 1037.29
R14931 fout3.n9 fout3.t12 797.225
R14932 fout3.n520 fout3.t7 797.172
R14933 fout3.n378 fout3.t11 732.331
R14934 fout3.n460 fout3.t9 731.671
R14935 fout3.n440 fout3.t13 731.671
R14936 fout3.n497 fout3.t8 730.672
R14937 fout3.n453 fout3.t10 400.616
R14938 fout3.n496 fout3.t3 400.614
R14939 fout3.n393 fout3.t14 397.311
R14940 fout3.n497 fout3.t4 395.84
R14941 fout3.n218 fout3.n217 13.176
R14942 fout3.n30 fout3.t0 11.73
R14943 fout3.n30 fout3.t2 10.985
R14944 fout3.n38 fout3.n36 9.3
R14945 fout3.n340 fout3.n339 9.3
R14946 fout3.n86 fout3.n85 9.3
R14947 fout3.n88 fout3.n87 9.3
R14948 fout3.n146 fout3.n145 9.3
R14949 fout3.n143 fout3.n142 9.3
R14950 fout3.n100 fout3.n99 9.3
R14951 fout3.n98 fout3.n97 9.3
R14952 fout3.n224 fout3.n223 9.3
R14953 fout3.n124 fout3.n123 9.3
R14954 fout3.n132 fout3.n131 9.3
R14955 fout3.n135 fout3.n134 9.3
R14956 fout3.n254 fout3.n253 9.3
R14957 fout3.n251 fout3.n250 9.3
R14958 fout3.n335 fout3.n334 9.3
R14959 fout3.n333 fout3.n332 9.3
R14960 fout3.n326 fout3.n325 8.097
R14961 fout3.n134 fout3.n133 5.457
R14962 fout3.n253 fout3.n252 5.08
R14963 fout3.n324 fout3.n323 4.65
R14964 fout3.n263 fout3.n262 4.65
R14965 fout3.n345 fout3.n338 4.5
R14966 fout3.n319 fout3.n318 4.5
R14967 fout3.n312 fout3.n311 4.5
R14968 fout3.n243 fout3.n242 4.5
R14969 fout3.n233 fout3.n232 4.5
R14970 fout3.n220 fout3.n219 4.5
R14971 fout3.n196 fout3.n195 4.5
R14972 fout3.n129 fout3.n120 4.5
R14973 fout3.n152 fout3.n151 4.5
R14974 fout3.n96 fout3.n95 4.5
R14975 fout3.n108 fout3.n107 4.5
R14976 fout3.n115 fout3.n114 4.5
R14977 fout3.n160 fout3.n159 4.5
R14978 fout3.n140 fout3.n139 4.5
R14979 fout3.n305 fout3.n304 4.5
R14980 fout3.n84 fout3.n83 4.5
R14981 fout3.n354 fout3.n351 4.5
R14982 fout3.n41 fout3.n40 4.5
R14983 fout3.n107 fout3.n105 4.314
R14984 fout3.n159 fout3.n156 3.944
R14985 fout3.n318 fout3.n317 3.937
R14986 fout3.n304 fout3.n303 3.567
R14987 fout3.n264 fout3.n257 3.033
R14988 fout3.n328 fout3.n327 3.033
R14989 fout3.n325 fout3.t1 2.9
R14990 fout3.n158 fout3.n157 2.258
R14991 fout3.n302 fout3.n301 2.258
R14992 fout3.n113 fout3.n112 1.882
R14993 fout3.n114 fout3.n113 1.882
R14994 fout3.n310 fout3.n309 1.882
R14995 fout3.n366 fout3.n30 1.64
R14996 fout3.n304 fout3.n302 1.505
R14997 fout3.n311 fout3.n310 1.505
R14998 fout3.n346 fout3.n345 1.5
R14999 fout3.n197 fout3.n196 1.5
R15000 fout3.n234 fout3.n233 1.5
R15001 fout3.n265 fout3.n264 1.5
R15002 fout3.n244 fout3.n243 1.5
R15003 fout3.n355 fout3.n354 1.5
R15004 fout3.n42 fout3.n41 1.5
R15005 fout3.n491 fout3.n490 1.435
R15006 fout3.n422 fout3.n421 1.435
R15007 fout3.n22 fout3.n8 1.388
R15008 fout3.n10 fout3.n9 1.354
R15009 fout3.n522 fout3.n520 1.354
R15010 fout3.n537 fout3.n536 1.354
R15011 fout3.n462 fout3.n460 1.354
R15012 fout3.n442 fout3.n440 1.354
R15013 fout3.n395 fout3.n393 1.354
R15014 fout3.n379 fout3.n378 1.354
R15015 fout3 fout3.n410 1.229
R15016 fout3.n396 fout3.n395 1.142
R15017 fout3.n523 fout3.n522 1.142
R15018 fout3.n423 fout3.n422 1.142
R15019 fout3.n463 fout3.n462 1.14
R15020 fout3.n397 fout3.n396 1.138
R15021 fout3.n435 fout3.n423 1.138
R15022 fout3.n524 fout3.n523 1.138
R15023 fout3.n380 fout3.n379 1.137
R15024 fout3.n406 fout3.n405 1.137
R15025 fout3.n371 fout3.n370 1.137
R15026 fout3.n401 fout3.n400 1.137
R15027 fout3.n386 fout3.n385 1.137
R15028 fout3.n477 fout3.n476 1.137
R15029 fout3.n468 fout3.n467 1.137
R15030 fout3.n473 fout3.n472 1.137
R15031 fout3.n483 fout3.n482 1.137
R15032 fout3.n492 fout3.n491 1.137
R15033 fout3.n538 fout3.n537 1.137
R15034 fout3.n507 fout3.n506 1.137
R15035 fout3.n529 fout3.n528 1.137
R15036 fout3.n503 fout3.n502 1.137
R15037 fout3.n513 fout3.n512 1.137
R15038 fout3.n432 fout3.n431 1.137
R15039 fout3.n448 fout3.n447 1.137
R15040 fout3.n427 fout3.n426 1.137
R15041 fout3.n414 fout3.n413 1.137
R15042 fout3.n443 fout3.n442 1.137
R15043 fout3.n408 fout3.n407 1.136
R15044 fout3.n509 fout3.n508 1.136
R15045 fout3.n434 fout3.n433 1.136
R15046 fout3.n382 fout3.n381 1.136
R15047 fout3.n540 fout3.n539 1.136
R15048 fout3.n494 fout3.n493 1.136
R15049 fout3.n451 fout3.n450 1.136
R15050 fout3.n83 fout3.n82 1.129
R15051 fout3.n159 fout3.n158 1.129
R15052 fout3.n151 fout3.n150 1.129
R15053 fout3.n161 fout3.n160 1.042
R15054 fout3.n54 fout3.n53 0.853
R15055 fout3.n178 fout3.n177 0.853
R15056 fout3.n267 fout3.n266 0.853
R15057 fout3.n361 fout3.n360 0.853
R15058 fout3.n410 fout3.n29 0.827
R15059 fout3.n40 fout3.n39 0.752
R15060 fout3.n232 fout3.n231 0.752
R15061 fout3.n242 fout3.n241 0.752
R15062 fout3.n318 fout3.n316 0.752
R15063 fout3.n338 fout3.n337 0.752
R15064 fout3.n351 fout3.n350 0.752
R15065 fout3.n44 fout3.n43 0.717
R15066 fout3.n366 fout3.n365 0.69
R15067 fout3.n367 fout3.n366 0.68
R15068 fout3.n223 fout3.n222 0.536
R15069 fout3.n123 fout3.n122 0.536
R15070 fout3.n145 fout3.n144 0.475
R15071 fout3.n262 fout3.n261 0.475
R15072 fout3.n410 fout3.n409 0.471
R15073 fout3.n23 fout3.n22 0.44
R15074 fout3.n327 fout3.n326 0.382
R15075 fout3.n94 fout3.n93 0.382
R15076 fout3.n95 fout3.n94 0.376
R15077 fout3.n107 fout3.n106 0.376
R15078 fout3.n139 fout3.n138 0.376
R15079 fout3.n120 fout3.n119 0.376
R15080 fout3.n195 fout3.n194 0.376
R15081 fout3.n219 fout3.n218 0.376
R15082 fout3.n82 fout3.n81 0.349
R15083 fout3.n337 fout3.n336 0.349
R15084 fout3.n499 fout3.n498 0.151
R15085 fout3.n496 fout3.n495 0.123
R15086 fout3.n453 fout3.n452 0.123
R15087 fout3.n454 fout3.n453 0.091
R15088 fout3.n393 fout3.n392 0.083
R15089 fout3.n378 fout3.n377 0.083
R15090 fout3.n460 fout3.n459 0.083
R15091 fout3.n440 fout3.n439 0.083
R15092 fout3.n8 fout3.n7 0.076
R15093 fout3.n520 fout3.n519 0.076
R15094 fout3.n536 fout3.n535 0.076
R15095 fout3.n498 fout3.n496 0.07
R15096 fout3.n487 fout3.n486 0.064
R15097 fout3.n4 fout3.n3 0.059
R15098 fout3 fout3.n541 0.055
R15099 fout3.n136 fout3.n135 0.047
R15100 fout3.n126 fout3.n125 0.047
R15101 fout3.n214 fout3.n213 0.047
R15102 fout3.n227 fout3.n226 0.047
R15103 fout3.n255 fout3.n254 0.047
R15104 fout3.n342 fout3.n341 0.047
R15105 fout3.n321 fout3.n320 0.043
R15106 fout3.n290 fout3.n289 0.043
R15107 fout3.n104 fout3.n103 0.041
R15108 fout3.n71 fout3.n70 0.041
R15109 fout3.n330 fout3.n329 0.035
R15110 fout3.n198 fout3.n197 0.035
R15111 fout3.n203 fout3.n202 0.035
R15112 fout3.n296 fout3.n295 0.035
R15113 fout3.n91 fout3.n90 0.034
R15114 fout3.n212 fout3.n211 0.034
R15115 fout3.n216 fout3.n215 0.034
R15116 fout3.n333 fout3.n331 0.034
R15117 fout3.n51 fout3.n50 0.034
R15118 fout3.n49 fout3.n48 0.034
R15119 fout3.n168 fout3.n167 0.034
R15120 fout3.n175 fout3.n174 0.034
R15121 fout3.n234 fout3.n210 0.034
R15122 fout3.n236 fout3.n235 0.034
R15123 fout3.n249 fout3.n248 0.034
R15124 fout3.n298 fout3.n297 0.034
R15125 fout3.n405 fout3.n403 0.032
R15126 fout3.n18 fout3.n17 0.032
R15127 fout3.n17 fout3.n16 0.032
R15128 fout3.n89 fout3.n88 0.032
R15129 fout3.n264 fout3.n263 0.032
R15130 fout3.n328 fout3.n324 0.032
R15131 fout3.n173 fout3.n172 0.032
R15132 fout3.n346 fout3.n298 0.032
R15133 fout3.n476 fout3.n475 0.032
R15134 fout3.n506 fout3.n504 0.032
R15135 fout3.n431 fout3.n429 0.032
R15136 fout3.n22 fout3.n21 0.032
R15137 fout3.n56 fout3.n55 0.031
R15138 fout3.n67 fout3.n66 0.031
R15139 fout3.n280 fout3.n279 0.031
R15140 fout3.n363 fout3.n362 0.031
R15141 fout3.n12 fout3.n11 0.03
R15142 fout3.n98 fout3.n96 0.03
R15143 fout3.n143 fout3.n141 0.03
R15144 fout3.n128 fout3.n127 0.03
R15145 fout3.n229 fout3.n228 0.03
R15146 fout3.n343 fout3.n342 0.03
R15147 fout3.n52 fout3.n51 0.03
R15148 fout3.n46 fout3.n45 0.03
R15149 fout3.n171 fout3.n170 0.03
R15150 fout3.n208 fout3.n207 0.03
R15151 fout3.n237 fout3.n236 0.03
R15152 fout3.n293 fout3.n292 0.03
R15153 fout3.n360 fout3.n359 0.03
R15154 fout3.n180 fout3.n179 0.03
R15155 fout3.n191 fout3.n190 0.03
R15156 fout3.n269 fout3.n268 0.03
R15157 fout3.n392 fout3.n391 0.028
R15158 fout3.n390 fout3.n389 0.028
R15159 fout3.n375 fout3.n374 0.028
R15160 fout3.n377 fout3.n376 0.028
R15161 fout3.n385 fout3.n384 0.028
R15162 fout3.n400 fout3.n399 0.028
R15163 fout3.n405 fout3.n404 0.028
R15164 fout3.n370 fout3.n368 0.028
R15165 fout3.n21 fout3.n20 0.028
R15166 fout3.n19 fout3.n18 0.028
R15167 fout3.n16 fout3.n15 0.028
R15168 fout3.n14 fout3.n13 0.028
R15169 fout3.n41 fout3.n38 0.028
R15170 fout3.n79 fout3.n78 0.028
R15171 fout3.n102 fout3.n101 0.028
R15172 fout3.n117 fout3.n116 0.028
R15173 fout3.n160 fout3.n118 0.028
R15174 fout3.n149 fout3.n148 0.028
R15175 fout3.n264 fout3.n256 0.028
R15176 fout3.n308 fout3.n307 0.028
R15177 fout3.n322 fout3.n321 0.028
R15178 fout3.n345 fout3.n335 0.028
R15179 fout3.n42 fout3.n34 0.028
R15180 fout3.n69 fout3.n68 0.028
R15181 fout3.n76 fout3.n75 0.028
R15182 fout3.n161 fout3.n77 0.028
R15183 fout3.n166 fout3.n165 0.028
R15184 fout3.n176 fout3.n175 0.028
R15185 fout3.n193 fout3.n192 0.028
R15186 fout3.n205 fout3.n204 0.028
R15187 fout3.n266 fout3.n265 0.028
R15188 fout3.n285 fout3.n284 0.028
R15189 fout3.n291 fout3.n290 0.028
R15190 fout3.n356 fout3.n355 0.028
R15191 fout3.n459 fout3.n458 0.028
R15192 fout3.n488 fout3.n487 0.028
R15193 fout3.n490 fout3.n489 0.028
R15194 fout3.n472 fout3.n471 0.028
R15195 fout3.n482 fout3.n480 0.028
R15196 fout3.n512 fout3.n511 0.028
R15197 fout3.n502 fout3.n501 0.028
R15198 fout3.n506 fout3.n505 0.028
R15199 fout3.n528 fout3.n526 0.028
R15200 fout3.n439 fout3.n438 0.028
R15201 fout3.n437 fout3.n436 0.028
R15202 fout3.n419 fout3.n418 0.028
R15203 fout3.n421 fout3.n420 0.028
R15204 fout3.n447 fout3.n446 0.028
R15205 fout3.n426 fout3.n425 0.028
R15206 fout3.n431 fout3.n430 0.028
R15207 fout3.n413 fout3.n411 0.028
R15208 fout3.n60 fout3.n59 0.027
R15209 fout3.n63 fout3.n62 0.027
R15210 fout3.n7 fout3.n6 0.026
R15211 fout3.n5 fout3.n4 0.026
R15212 fout3.n3 fout3.n2 0.026
R15213 fout3.n1 fout3.n0 0.026
R15214 fout3.n86 fout3.n84 0.026
R15215 fout3.n140 fout3.n137 0.026
R15216 fout3.n259 fout3.n258 0.026
R15217 fout3.n306 fout3.n305 0.026
R15218 fout3.n163 fout3.n162 0.026
R15219 fout3.n177 fout3.n169 0.026
R15220 fout3.n247 fout3.n246 0.026
R15221 fout3.n283 fout3.n282 0.026
R15222 fout3.n288 fout3.n287 0.026
R15223 fout3.n358 fout3.n357 0.026
R15224 fout3.n184 fout3.n183 0.026
R15225 fout3.n187 fout3.n186 0.026
R15226 fout3.n273 fout3.n272 0.026
R15227 fout3.n276 fout3.n275 0.026
R15228 fout3.n519 fout3.n518 0.026
R15229 fout3.n517 fout3.n516 0.026
R15230 fout3.n533 fout3.n532 0.026
R15231 fout3.n535 fout3.n534 0.026
R15232 fout3.n43 fout3.n42 0.024
R15233 fout3.n147 fout3.n146 0.024
R15234 fout3.n263 fout3.n260 0.024
R15235 fout3.n33 fout3.n32 0.024
R15236 fout3.n73 fout3.n72 0.024
R15237 fout3.n169 fout3.n168 0.024
R15238 fout3.n201 fout3.n200 0.024
R15239 fout3.n244 fout3.n238 0.024
R15240 fout3.n26 fout3.n25 0.023
R15241 fout3.n110 fout3.n109 0.022
R15242 fout3.n137 fout3.n136 0.022
R15243 fout3.n124 fout3.n121 0.022
R15244 fout3.n224 fout3.n221 0.022
R15245 fout3.n260 fout3.n259 0.022
R15246 fout3.n315 fout3.n314 0.022
R15247 fout3.n32 fout3.n31 0.022
R15248 fout3.n177 fout3.n176 0.022
R15249 fout3.n200 fout3.n199 0.022
R15250 fout3.n265 fout3.n249 0.022
R15251 fout3.n248 fout3.n247 0.022
R15252 fout3.n154 fout3.n153 0.02
R15253 fout3.n152 fout3.n149 0.02
R15254 fout3.n148 fout3.n147 0.02
R15255 fout3.n256 fout3.n255 0.02
R15256 fout3.n240 fout3.n239 0.02
R15257 fout3.n53 fout3.n52 0.02
R15258 fout3.n167 fout3.n166 0.02
R15259 fout3.n266 fout3.n237 0.02
R15260 fout3.n359 fout3.n358 0.02
R15261 fout3.n355 fout3.n349 0.02
R15262 fout3.n54 fout3.n44 0.019
R15263 fout3.n55 fout3.n54 0.019
R15264 fout3.n361 fout3.n280 0.019
R15265 fout3.n362 fout3.n361 0.019
R15266 fout3.n324 fout3.n322 0.018
R15267 fout3.n74 fout3.n73 0.018
R15268 fout3.n360 fout3.n346 0.018
R15269 fout3.n178 fout3.n67 0.018
R15270 fout3.n179 fout3.n178 0.018
R15271 fout3.n267 fout3.n191 0.018
R15272 fout3.n268 fout3.n267 0.018
R15273 fout3.n395 fout3.n394 0.017
R15274 fout3.n385 fout3.n383 0.017
R15275 fout3.n370 fout3.n369 0.017
R15276 fout3.n379 fout3.n373 0.017
R15277 fout3.n13 fout3.n12 0.017
R15278 fout3.n11 fout3.n10 0.017
R15279 fout3.n101 fout3.n100 0.017
R15280 fout3.n130 fout3.n129 0.017
R15281 fout3.n127 fout3.n126 0.017
R15282 fout3.n353 fout3.n352 0.017
R15283 fout3.n162 fout3.n161 0.017
R15284 fout3.n165 fout3.n164 0.017
R15285 fout3.n174 fout3.n173 0.017
R15286 fout3.n172 fout3.n171 0.017
R15287 fout3.n246 fout3.n245 0.017
R15288 fout3.n287 fout3.n286 0.017
R15289 fout3.n292 fout3.n291 0.017
R15290 fout3.n349 fout3.n348 0.017
R15291 fout3.n462 fout3.n461 0.017
R15292 fout3.n467 fout3.n466 0.017
R15293 fout3.n482 fout3.n481 0.017
R15294 fout3.n491 fout3.n485 0.017
R15295 fout3.n522 fout3.n521 0.017
R15296 fout3.n512 fout3.n510 0.017
R15297 fout3.n528 fout3.n527 0.017
R15298 fout3.n537 fout3.n531 0.017
R15299 fout3.n442 fout3.n441 0.017
R15300 fout3.n447 fout3.n445 0.017
R15301 fout3.n413 fout3.n412 0.017
R15302 fout3.n422 fout3.n417 0.017
R15303 fout3.n401 fout3.n398 0.016
R15304 fout3.n406 fout3.n402 0.016
R15305 fout3.n473 fout3.n469 0.016
R15306 fout3.n478 fout3.n477 0.016
R15307 fout3.n503 fout3.n500 0.016
R15308 fout3.n432 fout3.n428 0.016
R15309 fout3.n391 fout3.n390 0.015
R15310 fout3.n376 fout3.n375 0.015
R15311 fout3.n20 fout3.n19 0.015
R15312 fout3.n15 fout3.n14 0.015
R15313 fout3.n80 fout3.n79 0.015
R15314 fout3.n90 fout3.n89 0.015
R15315 fout3.n118 fout3.n117 0.015
R15316 fout3.n228 fout3.n227 0.015
R15317 fout3.n233 fout3.n230 0.015
R15318 fout3.n307 fout3.n306 0.015
R15319 fout3.n312 fout3.n308 0.015
R15320 fout3.n344 fout3.n343 0.015
R15321 fout3.n50 fout3.n49 0.015
R15322 fout3.n48 fout3.n47 0.015
R15323 fout3.n77 fout3.n76 0.015
R15324 fout3.n207 fout3.n206 0.015
R15325 fout3.n210 fout3.n209 0.015
R15326 fout3.n235 fout3.n234 0.015
R15327 fout3.n284 fout3.n283 0.015
R15328 fout3.n286 fout3.n285 0.015
R15329 fout3.n458 fout3.n457 0.015
R15330 fout3.n489 fout3.n488 0.015
R15331 fout3.n471 fout3.n470 0.015
R15332 fout3.n480 fout3.n479 0.015
R15333 fout3.n438 fout3.n437 0.015
R15334 fout3.n420 fout3.n419 0.015
R15335 fout3.n6 fout3.n5 0.013
R15336 fout3.n2 fout3.n1 0.013
R15337 fout3.n92 fout3.n91 0.013
R15338 fout3.n116 fout3.n115 0.013
R15339 fout3.n132 fout3.n130 0.013
R15340 fout3.n329 fout3.n328 0.013
R15341 fout3.n331 fout3.n330 0.013
R15342 fout3.n75 fout3.n74 0.013
R15343 fout3.n295 fout3.n294 0.013
R15344 fout3.n297 fout3.n296 0.013
R15345 fout3.n365 fout3.n364 0.013
R15346 fout3.n518 fout3.n517 0.013
R15347 fout3.n534 fout3.n533 0.013
R15348 fout3.n407 fout3.n401 0.012
R15349 fout3.n407 fout3.n406 0.012
R15350 fout3.n61 fout3.n60 0.012
R15351 fout3.n62 fout3.n61 0.012
R15352 fout3.n474 fout3.n473 0.012
R15353 fout3.n477 fout3.n474 0.012
R15354 fout3.n508 fout3.n503 0.012
R15355 fout3.n508 fout3.n507 0.012
R15356 fout3.n433 fout3.n427 0.012
R15357 fout3.n433 fout3.n432 0.012
R15358 fout3.n388 fout3.n387 0.011
R15359 fout3.n381 fout3.n372 0.011
R15360 fout3.n155 fout3.n154 0.011
R15361 fout3.n58 fout3.n57 0.011
R15362 fout3.n65 fout3.n64 0.011
R15363 fout3.n182 fout3.n181 0.011
R15364 fout3.n185 fout3.n184 0.011
R15365 fout3.n186 fout3.n185 0.011
R15366 fout3.n189 fout3.n188 0.011
R15367 fout3.n271 fout3.n270 0.011
R15368 fout3.n274 fout3.n273 0.011
R15369 fout3.n275 fout3.n274 0.011
R15370 fout3.n278 fout3.n277 0.011
R15371 fout3.n465 fout3.n464 0.011
R15372 fout3.n493 fout3.n484 0.011
R15373 fout3.n515 fout3.n514 0.011
R15374 fout3.n539 fout3.n530 0.011
R15375 fout3.n450 fout3.n449 0.011
R15376 fout3.n416 fout3.n415 0.011
R15377 fout3.n469 fout3.n468 0.01
R15378 fout3.n483 fout3.n478 0.01
R15379 fout3.n529 fout3.n525 0.01
R15380 fout3.n448 fout3.n444 0.01
R15381 fout3.n24 fout3.n23 0.01
R15382 fout3.n25 fout3.n24 0.01
R15383 fout3.n28 fout3.n27 0.009
R15384 fout3.n38 fout3.n37 0.009
R15385 fout3.n111 fout3.n110 0.009
R15386 fout3.n115 fout3.n111 0.009
R15387 fout3.n213 fout3.n212 0.009
R15388 fout3.n314 fout3.n313 0.009
R15389 fout3.n34 fout3.n33 0.009
R15390 fout3.n199 fout3.n198 0.009
R15391 fout3.n108 fout3.n104 0.007
R15392 fout3.n215 fout3.n214 0.007
R15393 fout3.n221 fout3.n220 0.007
R15394 fout3.n313 fout3.n312 0.007
R15395 fout3.n341 fout3.n340 0.007
R15396 fout3.n72 fout3.n71 0.007
R15397 fout3.n197 fout3.n193 0.007
R15398 fout3.n202 fout3.n201 0.007
R15399 fout3.n204 fout3.n203 0.007
R15400 fout3.n357 fout3.n356 0.007
R15401 fout3.n348 fout3.n347 0.007
R15402 fout3.n387 fout3.n386 0.006
R15403 fout3.n372 fout3.n371 0.006
R15404 fout3.n381 fout3.n380 0.006
R15405 fout3.n57 fout3.n56 0.006
R15406 fout3.n59 fout3.n58 0.006
R15407 fout3.n64 fout3.n63 0.006
R15408 fout3.n66 fout3.n65 0.006
R15409 fout3.n181 fout3.n180 0.006
R15410 fout3.n183 fout3.n182 0.006
R15411 fout3.n188 fout3.n187 0.006
R15412 fout3.n190 fout3.n189 0.006
R15413 fout3.n270 fout3.n269 0.006
R15414 fout3.n272 fout3.n271 0.006
R15415 fout3.n277 fout3.n276 0.006
R15416 fout3.n279 fout3.n278 0.006
R15417 fout3.n364 fout3.n363 0.006
R15418 fout3.n468 fout3.n465 0.006
R15419 fout3.n484 fout3.n483 0.006
R15420 fout3.n493 fout3.n492 0.006
R15421 fout3.n514 fout3.n513 0.006
R15422 fout3.n530 fout3.n529 0.006
R15423 fout3.n539 fout3.n538 0.006
R15424 fout3.n450 fout3.n443 0.006
R15425 fout3.n449 fout3.n448 0.006
R15426 fout3.n415 fout3.n414 0.006
R15427 fout3.n27 fout3.n26 0.005
R15428 fout3.n29 fout3.n28 0.005
R15429 fout3.n84 fout3.n80 0.005
R15430 fout3.n88 fout3.n86 0.005
R15431 fout3.n160 fout3.n155 0.005
R15432 fout3.n153 fout3.n152 0.005
R15433 fout3.n125 fout3.n124 0.005
R15434 fout3.n225 fout3.n224 0.005
R15435 fout3.n300 fout3.n299 0.005
R15436 fout3.n320 fout3.n319 0.005
R15437 fout3.n245 fout3.n244 0.005
R15438 fout3.n289 fout3.n288 0.005
R15439 fout3.n409 fout3.n408 0.004
R15440 fout3.n434 fout3.n424 0.004
R15441 fout3.n509 fout3.n499 0.004
R15442 fout3.n464 fout3.n463 0.003
R15443 fout3.n382 fout3.n367 0.003
R15444 fout3.n541 fout3.n540 0.003
R15445 fout3.n495 fout3.n494 0.003
R15446 fout3.n452 fout3.n451 0.003
R15447 fout3.n41 fout3.n35 0.003
R15448 fout3.n233 fout3.n229 0.003
R15449 fout3.n254 fout3.n251 0.003
R15450 fout3.n243 fout3.n240 0.003
R15451 fout3.n319 fout3.n315 0.003
R15452 fout3.n335 fout3.n333 0.003
R15453 fout3.n345 fout3.n344 0.003
R15454 fout3.n354 fout3.n353 0.003
R15455 fout3.n164 fout3.n163 0.003
R15456 fout3.n294 fout3.n293 0.003
R15457 fout3.n396 fout3.n388 0.003
R15458 fout3.n523 fout3.n515 0.003
R15459 fout3.n423 fout3.n416 0.003
R15460 fout3.n455 fout3.n454 0.002
R15461 fout3.n456 fout3.n455 0.002
R15462 fout3.n408 fout3.n397 0.002
R15463 fout3.n524 fout3.n509 0.002
R15464 fout3.n435 fout3.n434 0.002
R15465 fout3.n397 fout3.n382 0.002
R15466 fout3.n451 fout3.n435 0.002
R15467 fout3.n540 fout3.n524 0.002
R15468 fout3.n494 fout3.n456 0.002
R15469 fout3.n96 fout3.n92 0.001
R15470 fout3.n100 fout3.n98 0.001
R15471 fout3.n103 fout3.n102 0.001
R15472 fout3.n109 fout3.n108 0.001
R15473 fout3.n146 fout3.n143 0.001
R15474 fout3.n141 fout3.n140 0.001
R15475 fout3.n135 fout3.n132 0.001
R15476 fout3.n129 fout3.n128 0.001
R15477 fout3.n220 fout3.n216 0.001
R15478 fout3.n226 fout3.n225 0.001
R15479 fout3.n305 fout3.n300 0.001
R15480 fout3.n47 fout3.n46 0.001
R15481 fout3.n70 fout3.n69 0.001
R15482 fout3.n206 fout3.n205 0.001
R15483 fout3.n209 fout3.n208 0.001
R15484 fout3.n282 fout3.n281 0.001
R15485 fout3.n498 fout3.n497 0.001
R15486 fout.n388 fout.t4 1037.29
R15487 fout.n389 fout.t6 797.185
R15488 fout.n341 fout.t5 732.331
R15489 fout.n372 fout.t3 397.315
R15490 fout.n229 fout.n228 13.176
R15491 fout.n335 fout.t2 11.722
R15492 fout.n335 fout.t0 10.994
R15493 fout.n8 fout.n7 9.3
R15494 fout.n307 fout.n306 9.3
R15495 fout.n273 fout.n272 9.3
R15496 fout.n270 fout.n269 9.3
R15497 fout.n207 fout.n206 9.3
R15498 fout.n321 fout.n320 9.3
R15499 fout.n323 fout.n322 9.3
R15500 fout.n205 fout.n204 9.3
R15501 fout.n238 fout.n237 9.3
R15502 fout.n251 fout.n250 9.3
R15503 fout.n259 fout.n258 9.3
R15504 fout.n262 fout.n261 9.3
R15505 fout.n122 fout.n121 9.3
R15506 fout.n119 fout.n118 9.3
R15507 fout.n35 fout.n34 9.3
R15508 fout.n33 fout.n32 9.3
R15509 fout.n26 fout.n25 8.097
R15510 fout.n261 fout.n260 5.457
R15511 fout.n121 fout.n120 5.08
R15512 fout.n24 fout.n23 4.65
R15513 fout.n131 fout.n130 4.65
R15514 fout.n40 fout.n38 4.5
R15515 fout.n92 fout.n88 4.5
R15516 fout.n96 fout.n85 4.5
R15517 fout.n111 fout.n110 4.5
R15518 fout.n66 fout.n65 4.5
R15519 fout.n240 fout.n232 4.5
R15520 fout.n247 fout.n230 4.5
R15521 fout.n256 fout.n227 4.5
R15522 fout.n279 fout.n278 4.5
R15523 fout.n327 fout.n326 4.5
R15524 fout.n315 fout.n314 4.5
R15525 fout.n215 fout.n214 4.5
R15526 fout.n222 fout.n221 4.5
R15527 fout.n287 fout.n286 4.5
R15528 fout.n267 fout.n266 4.5
R15529 fout.n104 fout.n103 4.5
R15530 fout.n198 fout.n197 4.5
R15531 fout.n12 fout.n10 4.5
R15532 fout.n214 fout.n212 4.314
R15533 fout.n286 fout.n283 3.944
R15534 fout.n88 fout.n87 3.937
R15535 fout.n103 fout.n102 3.567
R15536 fout.n132 fout.n125 3.033
R15537 fout.n28 fout.n27 3.033
R15538 fout.n25 fout.t1 2.9
R15539 fout.n285 fout.n284 2.258
R15540 fout.n101 fout.n100 2.258
R15541 fout.n220 fout.n219 1.882
R15542 fout.n221 fout.n220 1.882
R15543 fout.n84 fout.n83 1.882
R15544 fout.n336 fout.n335 1.518
R15545 fout.n103 fout.n101 1.505
R15546 fout.n85 fout.n84 1.505
R15547 fout.n41 fout.n40 1.5
R15548 fout.n328 fout.n327 1.5
R15549 fout.n67 fout.n66 1.5
R15550 fout.n133 fout.n132 1.5
R15551 fout.n112 fout.n111 1.5
R15552 fout.n199 fout.n198 1.5
R15553 fout.n13 fout.n12 1.5
R15554 fout.n402 fout.n388 1.388
R15555 fout.n390 fout.n389 1.355
R15556 fout.n343 fout.n341 1.354
R15557 fout.n373 fout.n372 1.354
R15558 fout.n344 fout.n343 1.14
R15559 fout.n358 fout.n357 1.137
R15560 fout.n349 fout.n348 1.137
R15561 fout.n354 fout.n353 1.137
R15562 fout.n364 fout.n363 1.137
R15563 fout.n374 fout.n373 1.137
R15564 fout.n376 fout.n375 1.136
R15565 fout.n326 fout.n325 1.129
R15566 fout.n286 fout.n285 1.129
R15567 fout.n278 fout.n277 1.129
R15568 fout.n288 fout.n287 1.042
R15569 fout.n330 fout.n329 0.853
R15570 fout.n177 fout.n176 0.853
R15571 fout.n135 fout.n134 0.853
R15572 fout.n43 fout.n42 0.853
R15573 fout.n410 fout.n409 0.823
R15574 fout.n197 fout.n196 0.752
R15575 fout.n65 fout.n64 0.752
R15576 fout.n110 fout.n109 0.752
R15577 fout.n88 fout.n86 0.752
R15578 fout.n38 fout.n37 0.752
R15579 fout.n10 fout.n9 0.752
R15580 fout.n15 fout.n14 0.716
R15581 fout.n336 fout.n334 0.689
R15582 fout.n337 fout.n336 0.68
R15583 fout.n237 fout.n236 0.536
R15584 fout.n250 fout.n249 0.536
R15585 fout.n130 fout.n129 0.476
R15586 fout.n272 fout.n271 0.475
R15587 fout.n410 fout.n379 0.471
R15588 fout.n403 fout.n402 0.44
R15589 fout.n27 fout.n26 0.382
R15590 fout.n313 fout.n312 0.382
R15591 fout.n314 fout.n313 0.376
R15592 fout.n214 fout.n213 0.376
R15593 fout.n266 fout.n265 0.376
R15594 fout.n227 fout.n226 0.376
R15595 fout.n230 fout.n229 0.376
R15596 fout.n232 fout.n231 0.376
R15597 fout.n37 fout.n36 0.35
R15598 fout.n325 fout.n324 0.349
R15599 fout fout.n410 0.187
R15600 fout.n341 fout.n340 0.083
R15601 fout.n372 fout.n371 0.083
R15602 fout.n388 fout.n387 0.075
R15603 fout.n368 fout.n367 0.064
R15604 fout.n384 fout.n383 0.058
R15605 fout.n309 fout.n308 0.047
R15606 fout.n263 fout.n262 0.047
R15607 fout.n253 fout.n252 0.047
R15608 fout.n244 fout.n243 0.047
R15609 fout.n234 fout.n233 0.047
R15610 fout.n123 fout.n122 0.047
R15611 fout.n6 fout.n5 0.047
R15612 fout.n91 fout.n90 0.043
R15613 fout.n73 fout.n72 0.043
R15614 fout.n211 fout.n210 0.041
R15615 fout.n296 fout.n295 0.041
R15616 fout.n30 fout.n29 0.035
R15617 fout.n166 fout.n165 0.035
R15618 fout.n161 fout.n160 0.035
R15619 fout.n20 fout.n19 0.035
R15620 fout.n318 fout.n317 0.034
R15621 fout.n246 fout.n245 0.034
R15622 fout.n242 fout.n241 0.034
R15623 fout.n33 fout.n31 0.034
R15624 fout.n305 fout.n304 0.034
R15625 fout.n303 fout.n302 0.034
R15626 fout.n155 fout.n154 0.034
R15627 fout.n174 fout.n173 0.034
R15628 fout.n67 fout.n60 0.034
R15629 fout.n69 fout.n68 0.034
R15630 fout.n117 fout.n116 0.034
R15631 fout.n22 fout.n21 0.034
R15632 fout.n397 fout.n396 0.032
R15633 fout.n398 fout.n397 0.032
R15634 fout.n357 fout.n356 0.032
R15635 fout.n321 fout.n319 0.032
R15636 fout.n132 fout.n131 0.032
R15637 fout.n28 fout.n24 0.032
R15638 fout.n172 fout.n171 0.032
R15639 fout.n41 fout.n22 0.032
R15640 fout.n402 fout.n401 0.032
R15641 fout.n332 fout.n331 0.031
R15642 fout.n190 fout.n189 0.031
R15643 fout.n179 fout.n178 0.031
R15644 fout.n148 fout.n147 0.031
R15645 fout.n137 fout.n136 0.031
R15646 fout.n56 fout.n55 0.031
R15647 fout.n45 fout.n44 0.031
R15648 fout.n392 fout.n391 0.03
R15649 fout.n270 fout.n268 0.03
R15650 fout.n255 fout.n254 0.03
R15651 fout.n62 fout.n61 0.03
R15652 fout.n5 fout.n4 0.03
R15653 fout.n328 fout.n305 0.03
R15654 fout.n300 fout.n299 0.03
R15655 fout.n170 fout.n169 0.03
R15656 fout.n58 fout.n57 0.03
R15657 fout.n70 fout.n69 0.03
R15658 fout.n17 fout.n16 0.03
R15659 fout.n394 fout.n393 0.028
R15660 fout.n396 fout.n395 0.028
R15661 fout.n399 fout.n398 0.028
R15662 fout.n401 fout.n400 0.028
R15663 fout.n340 fout.n339 0.028
R15664 fout.n369 fout.n368 0.028
R15665 fout.n371 fout.n370 0.028
R15666 fout.n353 fout.n352 0.028
R15667 fout.n363 fout.n361 0.028
R15668 fout.n310 fout.n309 0.028
R15669 fout.n209 fout.n208 0.028
R15670 fout.n224 fout.n223 0.028
R15671 fout.n287 fout.n225 0.028
R15672 fout.n276 fout.n275 0.028
R15673 fout.n132 fout.n124 0.028
R15674 fout.n98 fout.n97 0.028
R15675 fout.n90 fout.n89 0.028
R15676 fout.n40 fout.n35 0.028
R15677 fout.n12 fout.n8 0.028
R15678 fout.n200 fout.n199 0.028
R15679 fout.n329 fout.n203 0.028
R15680 fout.n298 fout.n297 0.028
R15681 fout.n291 fout.n290 0.028
R15682 fout.n289 fout.n288 0.028
R15683 fout.n153 fout.n152 0.028
R15684 fout.n175 fout.n174 0.028
R15685 fout.n168 fout.n167 0.028
R15686 fout.n159 fout.n158 0.028
R15687 fout.n134 fout.n133 0.028
R15688 fout.n78 fout.n77 0.028
R15689 fout.n72 fout.n71 0.028
R15690 fout.n13 fout.n3 0.028
R15691 fout.n186 fout.n185 0.027
R15692 fout.n183 fout.n182 0.027
R15693 fout.n144 fout.n143 0.027
R15694 fout.n141 fout.n140 0.027
R15695 fout.n52 fout.n51 0.027
R15696 fout.n49 fout.n48 0.027
R15697 fout.n327 fout.n323 0.026
R15698 fout.n267 fout.n264 0.026
R15699 fout.n127 fout.n126 0.026
R15700 fout.n104 fout.n99 0.026
R15701 fout.n150 fout.n149 0.026
R15702 fout.n176 fout.n156 0.026
R15703 fout.n115 fout.n114 0.026
R15704 fout.n80 fout.n79 0.026
R15705 fout.n75 fout.n74 0.026
R15706 fout.n2 fout.n1 0.026
R15707 fout.n381 fout.n380 0.025
R15708 fout.n383 fout.n382 0.025
R15709 fout.n385 fout.n384 0.025
R15710 fout.n387 fout.n386 0.025
R15711 fout.n14 fout.n13 0.024
R15712 fout.n274 fout.n273 0.024
R15713 fout.n131 fout.n128 0.024
R15714 fout.n202 fout.n201 0.024
R15715 fout.n294 fout.n293 0.024
R15716 fout.n156 fout.n155 0.024
R15717 fout.n163 fout.n162 0.024
R15718 fout.n112 fout.n82 0.024
R15719 fout.n406 fout.n405 0.023
R15720 fout.n217 fout.n216 0.022
R15721 fout.n264 fout.n263 0.022
R15722 fout.n251 fout.n248 0.022
R15723 fout.n239 fout.n238 0.022
R15724 fout.n128 fout.n127 0.022
R15725 fout.n94 fout.n93 0.022
R15726 fout.n203 fout.n202 0.022
R15727 fout.n176 fout.n175 0.022
R15728 fout.n164 fout.n163 0.022
R15729 fout.n133 fout.n117 0.022
R15730 fout.n116 fout.n115 0.022
R15731 fout.n281 fout.n280 0.02
R15732 fout.n279 fout.n276 0.02
R15733 fout.n275 fout.n274 0.02
R15734 fout.n124 fout.n123 0.02
R15735 fout.n108 fout.n107 0.02
R15736 fout.n199 fout.n193 0.02
R15737 fout.n329 fout.n328 0.02
R15738 fout.n154 fout.n153 0.02
R15739 fout.n134 fout.n70 0.02
R15740 fout.n1 fout.n0 0.02
R15741 fout.n331 fout.n330 0.019
R15742 fout.n330 fout.n190 0.019
R15743 fout.n178 fout.n177 0.019
R15744 fout.n177 fout.n148 0.019
R15745 fout.n136 fout.n135 0.019
R15746 fout.n135 fout.n56 0.019
R15747 fout.n44 fout.n43 0.019
R15748 fout.n43 fout.n15 0.019
R15749 fout.n293 fout.n292 0.018
R15750 fout.n42 fout.n41 0.018
R15751 fout.n391 fout.n390 0.017
R15752 fout.n393 fout.n392 0.017
R15753 fout.n343 fout.n342 0.017
R15754 fout.n348 fout.n347 0.017
R15755 fout.n363 fout.n362 0.017
R15756 fout.n373 fout.n366 0.017
R15757 fout.n195 fout.n194 0.017
R15758 fout.n208 fout.n207 0.017
R15759 fout.n257 fout.n256 0.017
R15760 fout.n254 fout.n253 0.017
R15761 fout.n193 fout.n192 0.017
R15762 fout.n299 fout.n298 0.017
R15763 fout.n152 fout.n151 0.017
R15764 fout.n173 fout.n172 0.017
R15765 fout.n171 fout.n170 0.017
R15766 fout.n169 fout.n168 0.017
R15767 fout.n114 fout.n113 0.017
R15768 fout.n82 fout.n81 0.017
R15769 fout.n76 fout.n75 0.017
R15770 fout.n354 fout.n350 0.016
R15771 fout.n359 fout.n358 0.016
R15772 fout.n395 fout.n394 0.015
R15773 fout.n400 fout.n399 0.015
R15774 fout.n339 fout.n338 0.015
R15775 fout.n370 fout.n369 0.015
R15776 fout.n352 fout.n351 0.015
R15777 fout.n361 fout.n360 0.015
R15778 fout.n311 fout.n310 0.015
R15779 fout.n319 fout.n318 0.015
R15780 fout.n225 fout.n224 0.015
R15781 fout.n66 fout.n63 0.015
R15782 fout.n99 fout.n98 0.015
R15783 fout.n97 fout.n96 0.015
R15784 fout.n304 fout.n303 0.015
R15785 fout.n302 fout.n301 0.015
R15786 fout.n290 fout.n289 0.015
R15787 fout.n60 fout.n59 0.015
R15788 fout.n68 fout.n67 0.015
R15789 fout.n79 fout.n78 0.015
R15790 fout.n77 fout.n76 0.015
R15791 fout.n382 fout.n381 0.013
R15792 fout.n386 fout.n385 0.013
R15793 fout.n317 fout.n316 0.013
R15794 fout.n223 fout.n222 0.013
R15795 fout.n259 fout.n257 0.013
R15796 fout.n29 fout.n28 0.013
R15797 fout.n31 fout.n30 0.013
R15798 fout.n292 fout.n291 0.013
R15799 fout.n19 fout.n18 0.013
R15800 fout.n21 fout.n20 0.013
R15801 fout.n334 fout.n333 0.013
R15802 fout.n355 fout.n354 0.012
R15803 fout.n358 fout.n355 0.012
R15804 fout.n185 fout.n184 0.012
R15805 fout.n184 fout.n183 0.012
R15806 fout.n143 fout.n142 0.012
R15807 fout.n142 fout.n141 0.012
R15808 fout.n51 fout.n50 0.012
R15809 fout.n50 fout.n49 0.012
R15810 fout.n346 fout.n345 0.011
R15811 fout.n375 fout.n365 0.011
R15812 fout.n282 fout.n281 0.011
R15813 fout.n107 fout.n106 0.011
R15814 fout.n188 fout.n187 0.011
R15815 fout.n181 fout.n180 0.011
R15816 fout.n146 fout.n145 0.011
R15817 fout.n139 fout.n138 0.011
R15818 fout.n54 fout.n53 0.011
R15819 fout.n47 fout.n46 0.011
R15820 fout.n350 fout.n349 0.01
R15821 fout.n364 fout.n359 0.01
R15822 fout.n405 fout.n404 0.01
R15823 fout.n404 fout.n403 0.01
R15824 fout.n408 fout.n407 0.009
R15825 fout.n308 fout.n307 0.009
R15826 fout.n218 fout.n217 0.009
R15827 fout.n222 fout.n218 0.009
R15828 fout.n245 fout.n244 0.009
R15829 fout.n95 fout.n94 0.009
R15830 fout.n201 fout.n200 0.009
R15831 fout.n165 fout.n164 0.009
R15832 fout.n215 fout.n211 0.007
R15833 fout.n248 fout.n247 0.007
R15834 fout.n243 fout.n242 0.007
R15835 fout.n240 fout.n239 0.007
R15836 fout.n96 fout.n95 0.007
R15837 fout.n8 fout.n6 0.007
R15838 fout.n295 fout.n294 0.007
R15839 fout.n167 fout.n166 0.007
R15840 fout.n162 fout.n161 0.007
R15841 fout.n160 fout.n159 0.007
R15842 fout.n3 fout.n2 0.007
R15843 fout.n349 fout.n346 0.006
R15844 fout.n365 fout.n364 0.006
R15845 fout.n375 fout.n374 0.006
R15846 fout.n333 fout.n332 0.006
R15847 fout.n189 fout.n188 0.006
R15848 fout.n187 fout.n186 0.006
R15849 fout.n182 fout.n181 0.006
R15850 fout.n180 fout.n179 0.006
R15851 fout.n147 fout.n146 0.006
R15852 fout.n145 fout.n144 0.006
R15853 fout.n140 fout.n139 0.006
R15854 fout.n138 fout.n137 0.006
R15855 fout.n55 fout.n54 0.006
R15856 fout.n53 fout.n52 0.006
R15857 fout.n48 fout.n47 0.006
R15858 fout.n46 fout.n45 0.006
R15859 fout.n409 fout.n408 0.005
R15860 fout.n407 fout.n406 0.005
R15861 fout.n327 fout.n311 0.005
R15862 fout.n323 fout.n321 0.005
R15863 fout.n287 fout.n282 0.005
R15864 fout.n280 fout.n279 0.005
R15865 fout.n252 fout.n251 0.005
R15866 fout.n238 fout.n235 0.005
R15867 fout.n106 fout.n105 0.005
R15868 fout.n92 fout.n91 0.005
R15869 fout.n192 fout.n191 0.005
R15870 fout.n113 fout.n112 0.005
R15871 fout.n74 fout.n73 0.005
R15872 fout.n345 fout.n344 0.003
R15873 fout.n376 fout.n337 0.003
R15874 fout.n198 fout.n195 0.003
R15875 fout.n66 fout.n62 0.003
R15876 fout.n122 fout.n119 0.003
R15877 fout.n111 fout.n108 0.003
R15878 fout.n93 fout.n92 0.003
R15879 fout.n35 fout.n33 0.003
R15880 fout.n40 fout.n39 0.003
R15881 fout.n12 fout.n11 0.003
R15882 fout.n151 fout.n150 0.003
R15883 fout.n18 fout.n17 0.003
R15884 fout.n379 fout.n378 0.002
R15885 fout.n378 fout.n377 0.002
R15886 fout.n377 fout.n376 0.002
R15887 fout.n316 fout.n315 0.001
R15888 fout.n207 fout.n205 0.001
R15889 fout.n210 fout.n209 0.001
R15890 fout.n216 fout.n215 0.001
R15891 fout.n273 fout.n270 0.001
R15892 fout.n268 fout.n267 0.001
R15893 fout.n262 fout.n259 0.001
R15894 fout.n256 fout.n255 0.001
R15895 fout.n247 fout.n246 0.001
R15896 fout.n241 fout.n240 0.001
R15897 fout.n235 fout.n234 0.001
R15898 fout.n105 fout.n104 0.001
R15899 fout.n301 fout.n300 0.001
R15900 fout.n297 fout.n296 0.001
R15901 fout.n158 fout.n157 0.001
R15902 fout.n59 fout.n58 0.001
R15903 fout.n81 fout.n80 0.001
R15904 a_n8558_5866.n97 a_n8558_5866.t4 1040.33
R15905 a_n8558_5866.n97 a_n8558_5866.t5 794.533
R15906 a_n8558_5866.n41 a_n8558_5866.n40 13.176
R15907 a_n8558_5866.n95 a_n8558_5866.t0 11.614
R15908 a_n8558_5866.n95 a_n8558_5866.t2 11.298
R15909 a_n8558_5866.n96 a_n8558_5866.t3 10.061
R15910 a_n8558_5866.n151 a_n8558_5866.n34 9.3
R15911 a_n8558_5866.n151 a_n8558_5866.n142 9.3
R15912 a_n8558_5866.n151 a_n8558_5866.n136 9.3
R15913 a_n8558_5866.n151 a_n8558_5866.n49 9.3
R15914 a_n8558_5866.n151 a_n8558_5866.n54 9.3
R15915 a_n8558_5866.n151 a_n8558_5866.n124 9.3
R15916 a_n8558_5866.n151 a_n8558_5866.n150 8.469
R15917 a_n8558_5866.n151 a_n8558_5866.n114 8.469
R15918 a_n8558_5866.n151 a_n8558_5866.n119 8.125
R15919 a_n8558_5866.n151 a_n8558_5866.n29 8.124
R15920 a_n8558_5866.n151 a_n8558_5866.n111 8.097
R15921 a_n8558_5866.n151 a_n8558_5866.n147 8.096
R15922 a_n8558_5866.n151 a_n8558_5866.n127 8.016
R15923 a_n8558_5866.n151 a_n8558_5866.n39 8.016
R15924 a_n8558_5866.n151 a_n8558_5866.n131 7.964
R15925 a_n8558_5866.n151 a_n8558_5866.n44 7.964
R15926 a_n8558_5866.n126 a_n8558_5866.n125 6.4
R15927 a_n8558_5866.n110 a_n8558_5866.n55 6.4
R15928 a_n8558_5866.n145 a_n8558_5866.n144 6.023
R15929 a_n8558_5866.n37 a_n8558_5866.n36 6.023
R15930 a_n8558_5866.n136 a_n8558_5866.n135 6.023
R15931 a_n8558_5866.n43 a_n8558_5866.n42 6.023
R15932 a_n8558_5866.n130 a_n8558_5866.n129 6.023
R15933 a_n8558_5866.n149 a_n8558_5866.n148 5.647
R15934 a_n8558_5866.n49 a_n8558_5866.n46 5.647
R15935 a_n8558_5866.n117 a_n8558_5866.n116 5.647
R15936 a_n8558_5866.n113 a_n8558_5866.n112 5.647
R15937 a_n8558_5866.n133 a_n8558_5866.n132 5.457
R15938 a_n8558_5866.n27 a_n8558_5866.n26 5.27
R15939 a_n8558_5866.n48 a_n8558_5866.n47 5.08
R15940 a_n8558_5866.n34 a_n8558_5866.n33 4.517
R15941 a_n8558_5866.n124 a_n8558_5866.n121 4.517
R15942 a_n8558_5866.n63 a_n8558_5866.n62 4.5
R15943 a_n8558_5866.n2 a_n8558_5866.n1 4.5
R15944 a_n8558_5866.n31 a_n8558_5866.n30 4.314
R15945 a_n8558_5866.n141 a_n8558_5866.n140 4.141
R15946 a_n8558_5866.n51 a_n8558_5866.n50 4.141
R15947 a_n8558_5866.n138 a_n8558_5866.n137 3.944
R15948 a_n8558_5866.n123 a_n8558_5866.n122 3.937
R15949 a_n8558_5866.n53 a_n8558_5866.n52 3.567
R15950 a_n8558_5866.n98 a_n8558_5866.n97 3.396
R15951 a_n8558_5866.n110 a_n8558_5866.n109 3.033
R15952 a_n8558_5866.t1 a_n8558_5866.n151 2.9
R15953 a_n8558_5866.n142 a_n8558_5866.n141 2.258
R15954 a_n8558_5866.n54 a_n8558_5866.n51 2.258
R15955 a_n8558_5866.n99 a_n8558_5866.n98 2.166
R15956 a_n8558_5866.n33 a_n8558_5866.n32 1.882
R15957 a_n8558_5866.n121 a_n8558_5866.n120 1.882
R15958 a_n8558_5866.n54 a_n8558_5866.n53 1.505
R15959 a_n8558_5866.n82 a_n8558_5866.n103 1.5
R15960 a_n8558_5866.n64 a_n8558_5866.n66 1.5
R15961 a_n8558_5866.n63 a_n8558_5866.n61 1.5
R15962 a_n8558_5866.n21 a_n8558_5866.n24 1.5
R15963 a_n8558_5866.n12 a_n8558_5866.n11 1.5
R15964 a_n8558_5866.n109 a_n8558_5866.n80 1.5
R15965 a_n8558_5866.n28 a_n8558_5866.n27 1.129
R15966 a_n8558_5866.n26 a_n8558_5866.n25 1.129
R15967 a_n8558_5866.n142 a_n8558_5866.n138 1.129
R15968 a_n8558_5866.n140 a_n8558_5866.n139 1.129
R15969 a_n8558_5866.n98 a_n8558_5866.n96 1.033
R15970 a_n8558_5866.n102 a_n8558_5866.n101 0.853
R15971 a_n8558_5866.n150 a_n8558_5866.n149 0.752
R15972 a_n8558_5866.n46 a_n8558_5866.n45 0.752
R15973 a_n8558_5866.n49 a_n8558_5866.n48 0.752
R15974 a_n8558_5866.n124 a_n8558_5866.n123 0.752
R15975 a_n8558_5866.n116 a_n8558_5866.n115 0.752
R15976 a_n8558_5866.n118 a_n8558_5866.n117 0.752
R15977 a_n8558_5866.n114 a_n8558_5866.n113 0.752
R15978 a_n8558_5866.n89 a_n8558_5866.n88 0.716
R15979 a_n8558_5866.n131 a_n8558_5866.n130 0.536
R15980 a_n8558_5866.n44 a_n8558_5866.n43 0.536
R15981 a_n8558_5866.n127 a_n8558_5866.n126 0.476
R15982 a_n8558_5866.n39 a_n8558_5866.n38 0.475
R15983 a_n8558_5866.n111 a_n8558_5866.n110 0.382
R15984 a_n8558_5866.n147 a_n8558_5866.n146 0.382
R15985 a_n8558_5866.n146 a_n8558_5866.n145 0.376
R15986 a_n8558_5866.n144 a_n8558_5866.n143 0.376
R15987 a_n8558_5866.n34 a_n8558_5866.n31 0.376
R15988 a_n8558_5866.n38 a_n8558_5866.n37 0.376
R15989 a_n8558_5866.n36 a_n8558_5866.n35 0.376
R15990 a_n8558_5866.n136 a_n8558_5866.n133 0.376
R15991 a_n8558_5866.n135 a_n8558_5866.n134 0.376
R15992 a_n8558_5866.n42 a_n8558_5866.n41 0.376
R15993 a_n8558_5866.n129 a_n8558_5866.n128 0.376
R15994 a_n8558_5866.n119 a_n8558_5866.n118 0.35
R15995 a_n8558_5866.n29 a_n8558_5866.n28 0.349
R15996 a_n8558_5866.n96 a_n8558_5866.n95 0.308
R15997 a_n8558_5866.n2 a_n8558_5866.n0 0.066
R15998 a_n8558_5866.n87 a_n8558_5866.n86 0.047
R15999 a_n8558_5866.n72 a_n8558_5866.n71 0.043
R16000 a_n8558_5866.n68 a_n8558_5866.n67 0.043
R16001 a_n8558_5866.n64 a_n8558_5866.n63 0.041
R16002 a_n8558_5866.n79 a_n8558_5866.n78 0.035
R16003 a_n8558_5866.n108 a_n8558_5866.n107 0.035
R16004 a_n8558_5866.n19 a_n8558_5866.n18 0.034
R16005 a_n8558_5866.n23 a_n8558_5866.n22 0.034
R16006 a_n8558_5866.n8 a_n8558_5866.n7 0.034
R16007 a_n8558_5866.n77 a_n8558_5866.n76 0.034
R16008 a_n8558_5866.n106 a_n8558_5866.n105 0.034
R16009 a_n8558_5866.n12 a_n8558_5866.n6 0.032
R16010 a_n8558_5866.n109 a_n8558_5866.n70 0.032
R16011 a_n8558_5866.n100 a_n8558_5866.n99 0.031
R16012 a_n8558_5866.n9 a_n8558_5866.n8 0.03
R16013 a_n8558_5866.n75 a_n8558_5866.n74 0.03
R16014 a_n8558_5866.n102 a_n8558_5866.n94 0.03
R16015 a_n8558_5866.n81 a_n8558_5866.n87 0.03
R16016 a_n8558_5866.n11 a_n8558_5866.n10 0.028
R16017 a_n8558_5866.n60 a_n8558_5866.n58 0.028
R16018 a_n8558_5866.n73 a_n8558_5866.n72 0.028
R16019 a_n8558_5866.n91 a_n8558_5866.n90 0.028
R16020 a_n8558_5866.n13 a_n8558_5866.n12 0.028
R16021 a_n8558_5866.n57 a_n8558_5866.n56 0.028
R16022 a_n8558_5866.n69 a_n8558_5866.n68 0.028
R16023 a_n8558_5866.n104 a_n8558_5866.n82 0.028
R16024 a_n8558_5866.n85 a_n8558_5866.n83 0.028
R16025 a_n8558_5866.n17 a_n8558_5866.n15 0.026
R16026 a_n8558_5866.n66 a_n8558_5866.n65 0.026
R16027 a_n8558_5866.n93 a_n8558_5866.n92 0.026
R16028 a_n8558_5866.n4 a_n8558_5866.n3 0.026
R16029 a_n8558_5866.n90 a_n8558_5866.n89 0.024
R16030 a_n8558_5866.n18 a_n8558_5866.n17 0.024
R16031 a_n8558_5866.n6 a_n8558_5866.n5 0.024
R16032 a_n8558_5866.n15 a_n8558_5866.n16 0.022
R16033 a_n8558_5866.n5 a_n8558_5866.n4 0.022
R16034 a_n8558_5866.n3 a_n8558_5866.n2 0.022
R16035 a_n8558_5866.n20 a_n8558_5866.n19 0.02
R16036 a_n8558_5866.n10 a_n8558_5866.n9 0.02
R16037 a_n8558_5866.n94 a_n8558_5866.n93 0.02
R16038 a_n8558_5866.n14 a_n8558_5866.n13 0.02
R16039 a_n8558_5866.n101 a_n8558_5866.n100 0.019
R16040 a_n8558_5866.n82 a_n8558_5866.n81 0.018
R16041 a_n8558_5866.n103 a_n8558_5866.n102 0.018
R16042 a_n8558_5866.n70 a_n8558_5866.n69 0.018
R16043 a_n8558_5866.n24 a_n8558_5866.n23 0.017
R16044 a_n8558_5866.n74 a_n8558_5866.n73 0.017
R16045 a_n8558_5866.n58 a_n8558_5866.n59 0.015
R16046 a_n8558_5866.n61 a_n8558_5866.n60 0.015
R16047 a_n8558_5866.n56 a_n8558_5866.n0 0.015
R16048 a_n8558_5866.n63 a_n8558_5866.n57 0.015
R16049 a_n8558_5866.n80 a_n8558_5866.n79 0.013
R16050 a_n8558_5866.n78 a_n8558_5866.n77 0.013
R16051 a_n8558_5866.n109 a_n8558_5866.n108 0.013
R16052 a_n8558_5866.n107 a_n8558_5866.n106 0.013
R16053 a_n8558_5866.n92 a_n8558_5866.n91 0.007
R16054 a_n8558_5866.n86 a_n8558_5866.n85 0.007
R16055 a_n8558_5866.n21 a_n8558_5866.n20 1.424
R16056 a_n8558_5866.n67 a_n8558_5866.n64 0.005
R16057 a_n8558_5866.n80 a_n8558_5866.n75 0.003
R16058 a_n8558_5866.n105 a_n8558_5866.n104 0.003
R16059 a_n8558_5866.n83 a_n8558_5866.n84 0.003
R16060 a_n8558_5866.n14 a_n8558_5866.n21 0.47
R16061 a_n12888_11551.n97 a_n12888_11551.t5 1040.28
R16062 a_n12888_11551.n97 a_n12888_11551.t4 794.529
R16063 a_n12888_11551.n50 a_n12888_11551.n49 13.176
R16064 a_n12888_11551.n98 a_n12888_11551.t3 11.611
R16065 a_n12888_11551.n98 a_n12888_11551.t2 11.295
R16066 a_n12888_11551.n99 a_n12888_11551.t1 10.373
R16067 a_n12888_11551.n138 a_n12888_11551.n39 9.3
R16068 a_n12888_11551.n138 a_n12888_11551.n134 9.3
R16069 a_n12888_11551.n138 a_n12888_11551.n128 9.3
R16070 a_n12888_11551.n138 a_n12888_11551.n58 9.3
R16071 a_n12888_11551.n138 a_n12888_11551.n66 9.3
R16072 a_n12888_11551.n138 a_n12888_11551.n123 9.3
R16073 a_n12888_11551.n138 a_n12888_11551.n118 8.47
R16074 a_n12888_11551.n138 a_n12888_11551.n137 8.469
R16075 a_n12888_11551.n138 a_n12888_11551.n115 8.124
R16076 a_n12888_11551.n138 a_n12888_11551.n29 8.124
R16077 a_n12888_11551.n138 a_n12888_11551.n34 8.097
R16078 a_n12888_11551.n138 a_n12888_11551.n110 8.097
R16079 a_n12888_11551.n138 a_n12888_11551.n61 8.016
R16080 a_n12888_11551.n138 a_n12888_11551.n44 8.016
R16081 a_n12888_11551.n138 a_n12888_11551.n53 7.964
R16082 a_n12888_11551.n138 a_n12888_11551.n48 7.964
R16083 a_n12888_11551.n60 a_n12888_11551.n59 6.4
R16084 a_n12888_11551.n109 a_n12888_11551.n67 6.4
R16085 a_n12888_11551.n32 a_n12888_11551.n31 6.023
R16086 a_n12888_11551.n42 a_n12888_11551.n41 6.023
R16087 a_n12888_11551.n128 a_n12888_11551.n127 6.023
R16088 a_n12888_11551.n47 a_n12888_11551.n46 6.023
R16089 a_n12888_11551.n52 a_n12888_11551.n51 6.023
R16090 a_n12888_11551.n136 a_n12888_11551.n135 5.647
R16091 a_n12888_11551.n58 a_n12888_11551.n55 5.647
R16092 a_n12888_11551.n113 a_n12888_11551.n112 5.647
R16093 a_n12888_11551.n117 a_n12888_11551.n116 5.647
R16094 a_n12888_11551.n125 a_n12888_11551.n124 5.457
R16095 a_n12888_11551.n27 a_n12888_11551.n26 5.27
R16096 a_n12888_11551.n57 a_n12888_11551.n56 5.08
R16097 a_n12888_11551.n39 a_n12888_11551.n38 4.517
R16098 a_n12888_11551.n123 a_n12888_11551.n120 4.517
R16099 a_n12888_11551.n75 a_n12888_11551.n74 4.5
R16100 a_n12888_11551.n2 a_n12888_11551.n1 4.5
R16101 a_n12888_11551.n36 a_n12888_11551.n35 4.314
R16102 a_n12888_11551.n133 a_n12888_11551.n132 4.141
R16103 a_n12888_11551.n63 a_n12888_11551.n62 4.141
R16104 a_n12888_11551.n130 a_n12888_11551.n129 3.944
R16105 a_n12888_11551.n122 a_n12888_11551.n121 3.937
R16106 a_n12888_11551.n65 a_n12888_11551.n64 3.567
R16107 a_n12888_11551.n100 a_n12888_11551.n97 3.395
R16108 a_n12888_11551.n109 a_n12888_11551.n108 3.033
R16109 a_n12888_11551.t0 a_n12888_11551.n138 2.9
R16110 a_n12888_11551.n101 a_n12888_11551.n100 2.399
R16111 a_n12888_11551.n134 a_n12888_11551.n133 2.258
R16112 a_n12888_11551.n66 a_n12888_11551.n63 2.258
R16113 a_n12888_11551.n38 a_n12888_11551.n37 1.882
R16114 a_n12888_11551.n120 a_n12888_11551.n119 1.882
R16115 a_n12888_11551.n66 a_n12888_11551.n65 1.505
R16116 a_n12888_11551.n94 a_n12888_11551.n102 1.5
R16117 a_n12888_11551.n76 a_n12888_11551.n78 1.5
R16118 a_n12888_11551.n75 a_n12888_11551.n73 1.5
R16119 a_n12888_11551.n21 a_n12888_11551.n24 1.5
R16120 a_n12888_11551.n12 a_n12888_11551.n11 1.5
R16121 a_n12888_11551.n108 a_n12888_11551.n92 1.5
R16122 a_n12888_11551.n28 a_n12888_11551.n27 1.129
R16123 a_n12888_11551.n26 a_n12888_11551.n25 1.129
R16124 a_n12888_11551.n134 a_n12888_11551.n130 1.129
R16125 a_n12888_11551.n132 a_n12888_11551.n131 1.129
R16126 a_n12888_11551.n100 a_n12888_11551.n99 1.022
R16127 a_n12888_11551.n137 a_n12888_11551.n136 0.752
R16128 a_n12888_11551.n55 a_n12888_11551.n54 0.752
R16129 a_n12888_11551.n58 a_n12888_11551.n57 0.752
R16130 a_n12888_11551.n123 a_n12888_11551.n122 0.752
R16131 a_n12888_11551.n112 a_n12888_11551.n111 0.752
R16132 a_n12888_11551.n114 a_n12888_11551.n113 0.752
R16133 a_n12888_11551.n118 a_n12888_11551.n117 0.752
R16134 a_n12888_11551.n53 a_n12888_11551.n52 0.536
R16135 a_n12888_11551.n48 a_n12888_11551.n47 0.536
R16136 a_n12888_11551.n61 a_n12888_11551.n60 0.475
R16137 a_n12888_11551.n44 a_n12888_11551.n43 0.475
R16138 a_n12888_11551.n34 a_n12888_11551.n33 0.382
R16139 a_n12888_11551.n110 a_n12888_11551.n109 0.382
R16140 a_n12888_11551.n33 a_n12888_11551.n32 0.376
R16141 a_n12888_11551.n31 a_n12888_11551.n30 0.376
R16142 a_n12888_11551.n39 a_n12888_11551.n36 0.376
R16143 a_n12888_11551.n43 a_n12888_11551.n42 0.376
R16144 a_n12888_11551.n41 a_n12888_11551.n40 0.376
R16145 a_n12888_11551.n128 a_n12888_11551.n125 0.376
R16146 a_n12888_11551.n127 a_n12888_11551.n126 0.376
R16147 a_n12888_11551.n46 a_n12888_11551.n45 0.376
R16148 a_n12888_11551.n51 a_n12888_11551.n50 0.376
R16149 a_n12888_11551.n29 a_n12888_11551.n28 0.349
R16150 a_n12888_11551.n115 a_n12888_11551.n114 0.349
R16151 a_n12888_11551.n99 a_n12888_11551.n98 0.316
R16152 a_n12888_11551.n94 a_n12888_11551.n93 0.15
R16153 a_n12888_11551.n101 a_n12888_11551.n95 0.148
R16154 a_n12888_11551.n2 a_n12888_11551.n0 0.066
R16155 a_n12888_11551.n84 a_n12888_11551.n83 0.043
R16156 a_n12888_11551.n80 a_n12888_11551.n79 0.043
R16157 a_n12888_11551.n76 a_n12888_11551.n75 0.041
R16158 a_n12888_11551.n91 a_n12888_11551.n90 0.035
R16159 a_n12888_11551.n107 a_n12888_11551.n106 0.035
R16160 a_n12888_11551.n19 a_n12888_11551.n18 0.034
R16161 a_n12888_11551.n23 a_n12888_11551.n22 0.034
R16162 a_n12888_11551.n8 a_n12888_11551.n7 0.034
R16163 a_n12888_11551.n89 a_n12888_11551.n88 0.034
R16164 a_n12888_11551.n105 a_n12888_11551.n104 0.034
R16165 a_n12888_11551.n12 a_n12888_11551.n6 0.032
R16166 a_n12888_11551.n108 a_n12888_11551.n82 0.032
R16167 a_n12888_11551.n9 a_n12888_11551.n8 0.03
R16168 a_n12888_11551.n87 a_n12888_11551.n86 0.03
R16169 a_n12888_11551.n11 a_n12888_11551.n10 0.028
R16170 a_n12888_11551.n72 a_n12888_11551.n70 0.028
R16171 a_n12888_11551.n85 a_n12888_11551.n84 0.028
R16172 a_n12888_11551.n13 a_n12888_11551.n12 0.028
R16173 a_n12888_11551.n69 a_n12888_11551.n68 0.028
R16174 a_n12888_11551.n81 a_n12888_11551.n80 0.028
R16175 a_n12888_11551.n103 a_n12888_11551.n94 0.028
R16176 a_n12888_11551.n17 a_n12888_11551.n15 0.026
R16177 a_n12888_11551.n78 a_n12888_11551.n77 0.026
R16178 a_n12888_11551.n4 a_n12888_11551.n3 0.026
R16179 a_n12888_11551.n18 a_n12888_11551.n17 0.024
R16180 a_n12888_11551.n6 a_n12888_11551.n5 0.024
R16181 a_n12888_11551.n15 a_n12888_11551.n16 0.022
R16182 a_n12888_11551.n5 a_n12888_11551.n4 0.022
R16183 a_n12888_11551.n3 a_n12888_11551.n2 0.022
R16184 a_n12888_11551.n20 a_n12888_11551.n19 0.02
R16185 a_n12888_11551.n10 a_n12888_11551.n9 0.02
R16186 a_n12888_11551.n14 a_n12888_11551.n13 0.02
R16187 a_n12888_11551.n102 a_n12888_11551.n101 0.018
R16188 a_n12888_11551.n82 a_n12888_11551.n81 0.018
R16189 a_n12888_11551.n24 a_n12888_11551.n23 0.017
R16190 a_n12888_11551.n86 a_n12888_11551.n85 0.017
R16191 a_n12888_11551.n70 a_n12888_11551.n71 0.015
R16192 a_n12888_11551.n73 a_n12888_11551.n72 0.015
R16193 a_n12888_11551.n68 a_n12888_11551.n0 0.015
R16194 a_n12888_11551.n75 a_n12888_11551.n69 0.015
R16195 a_n12888_11551.n92 a_n12888_11551.n91 0.013
R16196 a_n12888_11551.n90 a_n12888_11551.n89 0.013
R16197 a_n12888_11551.n108 a_n12888_11551.n107 0.013
R16198 a_n12888_11551.n106 a_n12888_11551.n105 0.013
R16199 a_n12888_11551.n95 a_n12888_11551.n96 0.007
R16200 a_n12888_11551.n21 a_n12888_11551.n20 1.424
R16201 a_n12888_11551.n79 a_n12888_11551.n76 0.005
R16202 a_n12888_11551.n92 a_n12888_11551.n87 0.003
R16203 a_n12888_11551.n104 a_n12888_11551.n103 0.003
R16204 a_n12888_11551.n14 a_n12888_11551.n21 0.47
R16205 a_n7083_11551.n97 a_n7083_11551.t4 1040.28
R16206 a_n7083_11551.n97 a_n7083_11551.t5 794.529
R16207 a_n7083_11551.n46 a_n7083_11551.n45 13.176
R16208 a_n7083_11551.n98 a_n7083_11551.t2 11.611
R16209 a_n7083_11551.n98 a_n7083_11551.t0 11.295
R16210 a_n7083_11551.n142 a_n7083_11551.n39 9.3
R16211 a_n7083_11551.n142 a_n7083_11551.n138 9.3
R16212 a_n7083_11551.n142 a_n7083_11551.n132 9.3
R16213 a_n7083_11551.n142 a_n7083_11551.n58 9.3
R16214 a_n7083_11551.n142 a_n7083_11551.n66 9.3
R16215 a_n7083_11551.n142 a_n7083_11551.n127 9.3
R16216 a_n7083_11551.n101 a_n7083_11551.t1 9.017
R16217 a_n7083_11551.n142 a_n7083_11551.n122 8.47
R16218 a_n7083_11551.n142 a_n7083_11551.n141 8.469
R16219 a_n7083_11551.n142 a_n7083_11551.n119 8.124
R16220 a_n7083_11551.n142 a_n7083_11551.n29 8.124
R16221 a_n7083_11551.n142 a_n7083_11551.n34 8.097
R16222 a_n7083_11551.n142 a_n7083_11551.n114 8.097
R16223 a_n7083_11551.n142 a_n7083_11551.n61 8.016
R16224 a_n7083_11551.n142 a_n7083_11551.n44 8.016
R16225 a_n7083_11551.n142 a_n7083_11551.n53 7.964
R16226 a_n7083_11551.n142 a_n7083_11551.n49 7.964
R16227 a_n7083_11551.n60 a_n7083_11551.n59 6.4
R16228 a_n7083_11551.n113 a_n7083_11551.n67 6.4
R16229 a_n7083_11551.n32 a_n7083_11551.n31 6.023
R16230 a_n7083_11551.n42 a_n7083_11551.n41 6.023
R16231 a_n7083_11551.n132 a_n7083_11551.n131 6.023
R16232 a_n7083_11551.n48 a_n7083_11551.n47 6.023
R16233 a_n7083_11551.n52 a_n7083_11551.n51 6.023
R16234 a_n7083_11551.n140 a_n7083_11551.n139 5.647
R16235 a_n7083_11551.n58 a_n7083_11551.n55 5.647
R16236 a_n7083_11551.n117 a_n7083_11551.n116 5.647
R16237 a_n7083_11551.n121 a_n7083_11551.n120 5.647
R16238 a_n7083_11551.n129 a_n7083_11551.n128 5.457
R16239 a_n7083_11551.n27 a_n7083_11551.n26 5.27
R16240 a_n7083_11551.n57 a_n7083_11551.n56 5.08
R16241 a_n7083_11551.n39 a_n7083_11551.n38 4.517
R16242 a_n7083_11551.n127 a_n7083_11551.n124 4.517
R16243 a_n7083_11551.n75 a_n7083_11551.n74 4.5
R16244 a_n7083_11551.n2 a_n7083_11551.n1 4.5
R16245 a_n7083_11551.n36 a_n7083_11551.n35 4.314
R16246 a_n7083_11551.n137 a_n7083_11551.n136 4.141
R16247 a_n7083_11551.n63 a_n7083_11551.n62 4.141
R16248 a_n7083_11551.n134 a_n7083_11551.n133 3.944
R16249 a_n7083_11551.n126 a_n7083_11551.n125 3.937
R16250 a_n7083_11551.n65 a_n7083_11551.n64 3.567
R16251 a_n7083_11551.n104 a_n7083_11551.n97 3.395
R16252 a_n7083_11551.n113 a_n7083_11551.n112 3.033
R16253 a_n7083_11551.t3 a_n7083_11551.n142 2.9
R16254 a_n7083_11551.n105 a_n7083_11551.n104 2.376
R16255 a_n7083_11551.n138 a_n7083_11551.n137 2.258
R16256 a_n7083_11551.n66 a_n7083_11551.n63 2.258
R16257 a_n7083_11551.n102 a_n7083_11551.n101 2.237
R16258 a_n7083_11551.n38 a_n7083_11551.n37 1.882
R16259 a_n7083_11551.n124 a_n7083_11551.n123 1.882
R16260 a_n7083_11551.n66 a_n7083_11551.n65 1.505
R16261 a_n7083_11551.n94 a_n7083_11551.n106 1.5
R16262 a_n7083_11551.n76 a_n7083_11551.n78 1.5
R16263 a_n7083_11551.n75 a_n7083_11551.n73 1.5
R16264 a_n7083_11551.n21 a_n7083_11551.n24 1.5
R16265 a_n7083_11551.n12 a_n7083_11551.n11 1.5
R16266 a_n7083_11551.n112 a_n7083_11551.n92 1.5
R16267 a_n7083_11551.n28 a_n7083_11551.n27 1.129
R16268 a_n7083_11551.n26 a_n7083_11551.n25 1.129
R16269 a_n7083_11551.n138 a_n7083_11551.n134 1.129
R16270 a_n7083_11551.n136 a_n7083_11551.n135 1.129
R16271 a_n7083_11551.n104 a_n7083_11551.n103 1.02
R16272 a_n7083_11551.n141 a_n7083_11551.n140 0.752
R16273 a_n7083_11551.n55 a_n7083_11551.n54 0.752
R16274 a_n7083_11551.n58 a_n7083_11551.n57 0.752
R16275 a_n7083_11551.n127 a_n7083_11551.n126 0.752
R16276 a_n7083_11551.n116 a_n7083_11551.n115 0.752
R16277 a_n7083_11551.n118 a_n7083_11551.n117 0.752
R16278 a_n7083_11551.n122 a_n7083_11551.n121 0.752
R16279 a_n7083_11551.n53 a_n7083_11551.n52 0.536
R16280 a_n7083_11551.n49 a_n7083_11551.n48 0.536
R16281 a_n7083_11551.n61 a_n7083_11551.n60 0.475
R16282 a_n7083_11551.n44 a_n7083_11551.n43 0.475
R16283 a_n7083_11551.n34 a_n7083_11551.n33 0.382
R16284 a_n7083_11551.n114 a_n7083_11551.n113 0.382
R16285 a_n7083_11551.n33 a_n7083_11551.n32 0.376
R16286 a_n7083_11551.n31 a_n7083_11551.n30 0.376
R16287 a_n7083_11551.n39 a_n7083_11551.n36 0.376
R16288 a_n7083_11551.n43 a_n7083_11551.n42 0.376
R16289 a_n7083_11551.n41 a_n7083_11551.n40 0.376
R16290 a_n7083_11551.n132 a_n7083_11551.n129 0.376
R16291 a_n7083_11551.n131 a_n7083_11551.n130 0.376
R16292 a_n7083_11551.n47 a_n7083_11551.n46 0.376
R16293 a_n7083_11551.n51 a_n7083_11551.n50 0.376
R16294 a_n7083_11551.n29 a_n7083_11551.n28 0.349
R16295 a_n7083_11551.n119 a_n7083_11551.n118 0.349
R16296 a_n7083_11551.n99 a_n7083_11551.n98 0.276
R16297 a_n7083_11551.n94 a_n7083_11551.n93 0.15
R16298 a_n7083_11551.n105 a_n7083_11551.n95 0.148
R16299 a_n7083_11551.n2 a_n7083_11551.n0 0.066
R16300 a_n7083_11551.n84 a_n7083_11551.n83 0.043
R16301 a_n7083_11551.n80 a_n7083_11551.n79 0.043
R16302 a_n7083_11551.n76 a_n7083_11551.n75 0.041
R16303 a_n7083_11551.n102 a_n7083_11551.n99 0.039
R16304 a_n7083_11551.n91 a_n7083_11551.n90 0.035
R16305 a_n7083_11551.n111 a_n7083_11551.n110 0.035
R16306 a_n7083_11551.n19 a_n7083_11551.n18 0.034
R16307 a_n7083_11551.n23 a_n7083_11551.n22 0.034
R16308 a_n7083_11551.n8 a_n7083_11551.n7 0.034
R16309 a_n7083_11551.n89 a_n7083_11551.n88 0.034
R16310 a_n7083_11551.n109 a_n7083_11551.n108 0.034
R16311 a_n7083_11551.n12 a_n7083_11551.n6 0.032
R16312 a_n7083_11551.n112 a_n7083_11551.n82 0.032
R16313 a_n7083_11551.n101 a_n7083_11551.n100 0.032
R16314 a_n7083_11551.n9 a_n7083_11551.n8 0.03
R16315 a_n7083_11551.n87 a_n7083_11551.n86 0.03
R16316 a_n7083_11551.n11 a_n7083_11551.n10 0.028
R16317 a_n7083_11551.n72 a_n7083_11551.n70 0.028
R16318 a_n7083_11551.n85 a_n7083_11551.n84 0.028
R16319 a_n7083_11551.n13 a_n7083_11551.n12 0.028
R16320 a_n7083_11551.n69 a_n7083_11551.n68 0.028
R16321 a_n7083_11551.n81 a_n7083_11551.n80 0.028
R16322 a_n7083_11551.n107 a_n7083_11551.n94 0.028
R16323 a_n7083_11551.n17 a_n7083_11551.n15 0.026
R16324 a_n7083_11551.n78 a_n7083_11551.n77 0.026
R16325 a_n7083_11551.n4 a_n7083_11551.n3 0.026
R16326 a_n7083_11551.n18 a_n7083_11551.n17 0.024
R16327 a_n7083_11551.n6 a_n7083_11551.n5 0.024
R16328 a_n7083_11551.n15 a_n7083_11551.n16 0.022
R16329 a_n7083_11551.n5 a_n7083_11551.n4 0.022
R16330 a_n7083_11551.n3 a_n7083_11551.n2 0.022
R16331 a_n7083_11551.n20 a_n7083_11551.n19 0.02
R16332 a_n7083_11551.n10 a_n7083_11551.n9 0.02
R16333 a_n7083_11551.n14 a_n7083_11551.n13 0.02
R16334 a_n7083_11551.n106 a_n7083_11551.n105 0.018
R16335 a_n7083_11551.n82 a_n7083_11551.n81 0.018
R16336 a_n7083_11551.n24 a_n7083_11551.n23 0.017
R16337 a_n7083_11551.n86 a_n7083_11551.n85 0.017
R16338 a_n7083_11551.n70 a_n7083_11551.n71 0.015
R16339 a_n7083_11551.n73 a_n7083_11551.n72 0.015
R16340 a_n7083_11551.n68 a_n7083_11551.n0 0.015
R16341 a_n7083_11551.n75 a_n7083_11551.n69 0.015
R16342 a_n7083_11551.n92 a_n7083_11551.n91 0.013
R16343 a_n7083_11551.n90 a_n7083_11551.n89 0.013
R16344 a_n7083_11551.n112 a_n7083_11551.n111 0.013
R16345 a_n7083_11551.n110 a_n7083_11551.n109 0.013
R16346 a_n7083_11551.n95 a_n7083_11551.n96 0.007
R16347 a_n7083_11551.n21 a_n7083_11551.n20 1.424
R16348 a_n7083_11551.n79 a_n7083_11551.n76 0.005
R16349 a_n7083_11551.n92 a_n7083_11551.n87 0.003
R16350 a_n7083_11551.n108 a_n7083_11551.n107 0.003
R16351 a_n7083_11551.n103 a_n7083_11551.n102 0.001
R16352 a_n7083_11551.n14 a_n7083_11551.n21 0.47
R16353 a_n12880_6001.n13 a_n12880_6001.t2 732.456
R16354 a_n12880_6001.n13 a_n12880_6001.t3 397.58
R16355 a_n12880_6001.n51 a_n12880_6001.n50 92.5
R16356 a_n12880_6001.n9 a_n12880_6001.n8 92.5
R16357 a_n12880_6001.n50 a_n12880_6001.t1 70.344
R16358 a_n12880_6001.n45 a_n12880_6001.n44 31.034
R16359 a_n12880_6001.n24 a_n12880_6001.n23 31.034
R16360 a_n12880_6001.n27 a_n12880_6001.n28 9.3
R16361 a_n12880_6001.n38 a_n12880_6001.n39 9.3
R16362 a_n12880_6001.n46 a_n12880_6001.n45 9.3
R16363 a_n12880_6001.n25 a_n12880_6001.n24 9.3
R16364 a_n12880_6001.n105 a_n12880_6001.n98 9.154
R16365 a_n12880_6001.n105 a_n12880_6001.n4 9.143
R16366 a_n12880_6001.n105 a_n12880_6001.n3 9.143
R16367 a_n12880_6001.n105 a_n12880_6001.n78 9.132
R16368 a_n12880_6001.n105 a_n12880_6001.n62 9.132
R16369 a_n12880_6001.n105 a_n12880_6001.n102 8.885
R16370 a_n12880_6001.n105 a_n12880_6001.n82 8.885
R16371 a_n12880_6001.n105 a_n12880_6001.n86 8.875
R16372 a_n12880_6001.n105 a_n12880_6001.n56 8.875
R16373 a_n12880_6001.n105 a_n12880_6001.n104 8.864
R16374 a_n12880_6001.n105 a_n12880_6001.n88 8.864
R16375 a_n12880_6001.n52 a_n12880_6001.n51 8.282
R16376 a_n12880_6001.n10 a_n12880_6001.n9 8.282
R16377 a_n12880_6001.t0 a_n12880_6001.n105 7.141
R16378 a_n12880_6001.n46 a_n12880_6001.n42 5.647
R16379 a_n12880_6001.n25 a_n12880_6001.n21 5.647
R16380 a_n12880_6001.n1 a_n12880_6001.n11 4.65
R16381 a_n12880_6001.n16 a_n12880_6001.n15 4.566
R16382 a_n12880_6001.n98 a_n12880_6001.n90 4.517
R16383 a_n12880_6001.n0 a_n12880_6001.n10 4.5
R16384 a_n12880_6001.n1 a_n12880_6001.n7 4.5
R16385 a_n12880_6001.n6 a_n12880_6001.n52 4.5
R16386 a_n12880_6001.n40 a_n12880_6001.n48 4.5
R16387 a_n12880_6001.n12 a_n12880_6001.n37 4.5
R16388 a_n12880_6001.n17 a_n12880_6001.n32 4.5
R16389 a_n12880_6001.n15 a_n12880_6001.n14 4.481
R16390 a_n12880_6001.n100 a_n12880_6001.n99 4.141
R16391 a_n12880_6001.n98 a_n12880_6001.n89 4.141
R16392 a_n12880_6001.n80 a_n12880_6001.n79 4.141
R16393 a_n12880_6001.n44 a_n12880_6001.n43 4.137
R16394 a_n12880_6001.n23 a_n12880_6001.n22 4.137
R16395 a_n12880_6001.n37 a_n12880_6001.n35 3.764
R16396 a_n12880_6001.n26 a_n12880_6001.n19 3.764
R16397 a_n12880_6001.n58 a_n12880_6001.n57 3.764
R16398 a_n12880_6001.n3 a_n12880_6001.n69 3.764
R16399 a_n12880_6001.n62 a_n12880_6001.n61 3.736
R16400 a_n12880_6001.n48 a_n12880_6001.n47 3.388
R16401 a_n12880_6001.n32 a_n12880_6001.n31 3.388
R16402 a_n12880_6001.n54 a_n12880_6001.n53 3.388
R16403 a_n12880_6001.n4 a_n12880_6001.n67 3.388
R16404 a_n12880_6001.n76 a_n12880_6001.n75 3.388
R16405 a_n12880_6001.n84 a_n12880_6001.n83 3.388
R16406 a_n12880_6001.n78 a_n12880_6001.n74 3.36
R16407 a_n12880_6001.n48 a_n12880_6001.n46 3.011
R16408 a_n12880_6001.n52 a_n12880_6001.n49 3.011
R16409 a_n12880_6001.n32 a_n12880_6001.n30 3.011
R16410 a_n12880_6001.n55 a_n12880_6001.n54 3.011
R16411 a_n12880_6001.n67 a_n12880_6001.n66 3.011
R16412 a_n12880_6001.n65 a_n12880_6001.n64 3.011
R16413 a_n12880_6001.n74 a_n12880_6001.n73 3.011
R16414 a_n12880_6001.n77 a_n12880_6001.n76 3.011
R16415 a_n12880_6001.n85 a_n12880_6001.n84 3.011
R16416 a_n12880_6001.n91 a_n12880_6001.n14 2.921
R16417 a_n12880_6001.n37 a_n12880_6001.n36 2.635
R16418 a_n12880_6001.n26 a_n12880_6001.n25 2.635
R16419 a_n12880_6001.n59 a_n12880_6001.n58 2.635
R16420 a_n12880_6001.n61 a_n12880_6001.n60 2.635
R16421 a_n12880_6001.n72 a_n12880_6001.n71 2.635
R16422 a_n12880_6001.n69 a_n12880_6001.n68 2.635
R16423 a_n12880_6001.n15 a_n12880_6001.n13 2.354
R16424 a_n12880_6001.n101 a_n12880_6001.n100 2.258
R16425 a_n12880_6001.n81 a_n12880_6001.n80 2.258
R16426 a_n12880_6001.n5 a_n12880_6001.n96 1.633
R16427 a_n12880_6001.n2 a_n12880_6001.n95 1.619
R16428 a_n12880_6001.n92 a_n12880_6001.n93 1.588
R16429 a_n12880_6001.n5 a_n12880_6001.n106 1.587
R16430 a_n12880_6001.n71 a_n12880_6001.n70 1.505
R16431 a_n12880_6001.n12 a_n12880_6001.n34 1.5
R16432 a_n12880_6001.n64 a_n12880_6001.n63 1.129
R16433 a_n12880_6001.n42 a_n12880_6001.n41 0.752
R16434 a_n12880_6001.n21 a_n12880_6001.n20 0.752
R16435 a_n12880_6001.n104 a_n12880_6001.n103 0.155
R16436 a_n12880_6001.n88 a_n12880_6001.n87 0.155
R16437 a_n12880_6001.n56 a_n12880_6001.n55 0.144
R16438 a_n12880_6001.n86 a_n12880_6001.n85 0.144
R16439 a_n12880_6001.n102 a_n12880_6001.n101 0.132
R16440 a_n12880_6001.n82 a_n12880_6001.n81 0.132
R16441 a_n12880_6001.n91 a_n12880_6001.n92 0.125
R16442 a_n12880_6001.n106 a_n12880_6001.n107 0.037
R16443 a_n12880_6001.n96 a_n12880_6001.n97 0.034
R16444 a_n12880_6001.n40 a_n12880_6001.n38 0.094
R16445 a_n12880_6001.n34 a_n12880_6001.n33 0.293
R16446 a_n12880_6001.n34 a_n12880_6001.n18 0.877
R16447 a_n12880_6001.n93 a_n12880_6001.n94 0.024
R16448 a_n12880_6001.n62 a_n12880_6001.n59 0.024
R16449 a_n12880_6001.n78 a_n12880_6001.n77 0.024
R16450 a_n12880_6001.n98 a_n12880_6001.n91 4.672
R16451 a_n12880_6001.n18 a_n12880_6001.n16 0.019
R16452 a_n12880_6001.n18 a_n12880_6001.n17 2.433
R16453 a_n12880_6001.n6 a_n12880_6001.n40 0.044
R16454 a_n12880_6001.n17 a_n12880_6001.n27 0.032
R16455 a_n12880_6001.n38 a_n12880_6001.n12 0.031
R16456 a_n12880_6001.n17 a_n12880_6001.n29 0.017
R16457 a_n12880_6001.n27 a_n12880_6001.n26 4.595
R16458 a_n12880_6001.n4 a_n12880_6001.n65 2.257
R16459 a_n12880_6001.n3 a_n12880_6001.n72 2.257
R16460 a_n12880_6001.n2 a_n12880_6001.n5 0.256
R16461 a_n12880_6001.n92 a_n12880_6001.n2 0.124
R16462 a_n12880_6001.n6 a_n12880_6001.n1 0.07
R16463 a_n12880_6001.n1 a_n12880_6001.n0 0.053
R16464 P7 P7.t1 1038.31
R16465 P7 P7.t0 796.504
R16466 a_n20175_5871.n97 a_n20175_5871.t5 1040.33
R16467 a_n20175_5871.n97 a_n20175_5871.t4 794.533
R16468 a_n20175_5871.n41 a_n20175_5871.n40 13.176
R16469 a_n20175_5871.n95 a_n20175_5871.t3 11.611
R16470 a_n20175_5871.n95 a_n20175_5871.t2 11.295
R16471 a_n20175_5871.n96 a_n20175_5871.t1 10.376
R16472 a_n20175_5871.n151 a_n20175_5871.n34 9.3
R16473 a_n20175_5871.n151 a_n20175_5871.n142 9.3
R16474 a_n20175_5871.n151 a_n20175_5871.n136 9.3
R16475 a_n20175_5871.n151 a_n20175_5871.n49 9.3
R16476 a_n20175_5871.n151 a_n20175_5871.n54 9.3
R16477 a_n20175_5871.n151 a_n20175_5871.n124 9.3
R16478 a_n20175_5871.n151 a_n20175_5871.n150 8.469
R16479 a_n20175_5871.n151 a_n20175_5871.n114 8.469
R16480 a_n20175_5871.n151 a_n20175_5871.n119 8.125
R16481 a_n20175_5871.n151 a_n20175_5871.n29 8.124
R16482 a_n20175_5871.n151 a_n20175_5871.n111 8.097
R16483 a_n20175_5871.n151 a_n20175_5871.n147 8.096
R16484 a_n20175_5871.n151 a_n20175_5871.n127 8.016
R16485 a_n20175_5871.n151 a_n20175_5871.n39 8.016
R16486 a_n20175_5871.n151 a_n20175_5871.n131 7.964
R16487 a_n20175_5871.n151 a_n20175_5871.n44 7.964
R16488 a_n20175_5871.n126 a_n20175_5871.n125 6.4
R16489 a_n20175_5871.n110 a_n20175_5871.n55 6.4
R16490 a_n20175_5871.n145 a_n20175_5871.n144 6.023
R16491 a_n20175_5871.n37 a_n20175_5871.n36 6.023
R16492 a_n20175_5871.n136 a_n20175_5871.n135 6.023
R16493 a_n20175_5871.n43 a_n20175_5871.n42 6.023
R16494 a_n20175_5871.n130 a_n20175_5871.n129 6.023
R16495 a_n20175_5871.n149 a_n20175_5871.n148 5.647
R16496 a_n20175_5871.n49 a_n20175_5871.n46 5.647
R16497 a_n20175_5871.n117 a_n20175_5871.n116 5.647
R16498 a_n20175_5871.n113 a_n20175_5871.n112 5.647
R16499 a_n20175_5871.n133 a_n20175_5871.n132 5.457
R16500 a_n20175_5871.n27 a_n20175_5871.n26 5.27
R16501 a_n20175_5871.n48 a_n20175_5871.n47 5.08
R16502 a_n20175_5871.n34 a_n20175_5871.n33 4.517
R16503 a_n20175_5871.n124 a_n20175_5871.n121 4.517
R16504 a_n20175_5871.n63 a_n20175_5871.n62 4.5
R16505 a_n20175_5871.n2 a_n20175_5871.n1 4.5
R16506 a_n20175_5871.n31 a_n20175_5871.n30 4.314
R16507 a_n20175_5871.n141 a_n20175_5871.n140 4.141
R16508 a_n20175_5871.n51 a_n20175_5871.n50 4.141
R16509 a_n20175_5871.n138 a_n20175_5871.n137 3.944
R16510 a_n20175_5871.n123 a_n20175_5871.n122 3.937
R16511 a_n20175_5871.n53 a_n20175_5871.n52 3.567
R16512 a_n20175_5871.n98 a_n20175_5871.n97 3.395
R16513 a_n20175_5871.n110 a_n20175_5871.n109 3.033
R16514 a_n20175_5871.t0 a_n20175_5871.n151 2.9
R16515 a_n20175_5871.n142 a_n20175_5871.n141 2.258
R16516 a_n20175_5871.n54 a_n20175_5871.n51 2.258
R16517 a_n20175_5871.n99 a_n20175_5871.n98 2.168
R16518 a_n20175_5871.n33 a_n20175_5871.n32 1.882
R16519 a_n20175_5871.n121 a_n20175_5871.n120 1.882
R16520 a_n20175_5871.n54 a_n20175_5871.n53 1.505
R16521 a_n20175_5871.n82 a_n20175_5871.n103 1.5
R16522 a_n20175_5871.n64 a_n20175_5871.n66 1.5
R16523 a_n20175_5871.n63 a_n20175_5871.n61 1.5
R16524 a_n20175_5871.n21 a_n20175_5871.n24 1.5
R16525 a_n20175_5871.n12 a_n20175_5871.n11 1.5
R16526 a_n20175_5871.n109 a_n20175_5871.n80 1.5
R16527 a_n20175_5871.n28 a_n20175_5871.n27 1.129
R16528 a_n20175_5871.n26 a_n20175_5871.n25 1.129
R16529 a_n20175_5871.n142 a_n20175_5871.n138 1.129
R16530 a_n20175_5871.n140 a_n20175_5871.n139 1.129
R16531 a_n20175_5871.n98 a_n20175_5871.n96 1.021
R16532 a_n20175_5871.n102 a_n20175_5871.n101 0.853
R16533 a_n20175_5871.n150 a_n20175_5871.n149 0.752
R16534 a_n20175_5871.n46 a_n20175_5871.n45 0.752
R16535 a_n20175_5871.n49 a_n20175_5871.n48 0.752
R16536 a_n20175_5871.n124 a_n20175_5871.n123 0.752
R16537 a_n20175_5871.n116 a_n20175_5871.n115 0.752
R16538 a_n20175_5871.n118 a_n20175_5871.n117 0.752
R16539 a_n20175_5871.n114 a_n20175_5871.n113 0.752
R16540 a_n20175_5871.n89 a_n20175_5871.n88 0.716
R16541 a_n20175_5871.n131 a_n20175_5871.n130 0.536
R16542 a_n20175_5871.n44 a_n20175_5871.n43 0.536
R16543 a_n20175_5871.n127 a_n20175_5871.n126 0.476
R16544 a_n20175_5871.n39 a_n20175_5871.n38 0.475
R16545 a_n20175_5871.n111 a_n20175_5871.n110 0.382
R16546 a_n20175_5871.n147 a_n20175_5871.n146 0.382
R16547 a_n20175_5871.n146 a_n20175_5871.n145 0.376
R16548 a_n20175_5871.n144 a_n20175_5871.n143 0.376
R16549 a_n20175_5871.n34 a_n20175_5871.n31 0.376
R16550 a_n20175_5871.n38 a_n20175_5871.n37 0.376
R16551 a_n20175_5871.n36 a_n20175_5871.n35 0.376
R16552 a_n20175_5871.n136 a_n20175_5871.n133 0.376
R16553 a_n20175_5871.n135 a_n20175_5871.n134 0.376
R16554 a_n20175_5871.n42 a_n20175_5871.n41 0.376
R16555 a_n20175_5871.n129 a_n20175_5871.n128 0.376
R16556 a_n20175_5871.n119 a_n20175_5871.n118 0.35
R16557 a_n20175_5871.n29 a_n20175_5871.n28 0.349
R16558 a_n20175_5871.n96 a_n20175_5871.n95 0.316
R16559 a_n20175_5871.n2 a_n20175_5871.n0 0.066
R16560 a_n20175_5871.n87 a_n20175_5871.n86 0.047
R16561 a_n20175_5871.n72 a_n20175_5871.n71 0.043
R16562 a_n20175_5871.n68 a_n20175_5871.n67 0.043
R16563 a_n20175_5871.n64 a_n20175_5871.n63 0.041
R16564 a_n20175_5871.n79 a_n20175_5871.n78 0.035
R16565 a_n20175_5871.n108 a_n20175_5871.n107 0.035
R16566 a_n20175_5871.n19 a_n20175_5871.n18 0.034
R16567 a_n20175_5871.n23 a_n20175_5871.n22 0.034
R16568 a_n20175_5871.n8 a_n20175_5871.n7 0.034
R16569 a_n20175_5871.n77 a_n20175_5871.n76 0.034
R16570 a_n20175_5871.n106 a_n20175_5871.n105 0.034
R16571 a_n20175_5871.n12 a_n20175_5871.n6 0.032
R16572 a_n20175_5871.n109 a_n20175_5871.n70 0.032
R16573 a_n20175_5871.n100 a_n20175_5871.n99 0.031
R16574 a_n20175_5871.n9 a_n20175_5871.n8 0.03
R16575 a_n20175_5871.n75 a_n20175_5871.n74 0.03
R16576 a_n20175_5871.n102 a_n20175_5871.n94 0.03
R16577 a_n20175_5871.n81 a_n20175_5871.n87 0.03
R16578 a_n20175_5871.n11 a_n20175_5871.n10 0.028
R16579 a_n20175_5871.n60 a_n20175_5871.n58 0.028
R16580 a_n20175_5871.n73 a_n20175_5871.n72 0.028
R16581 a_n20175_5871.n91 a_n20175_5871.n90 0.028
R16582 a_n20175_5871.n13 a_n20175_5871.n12 0.028
R16583 a_n20175_5871.n57 a_n20175_5871.n56 0.028
R16584 a_n20175_5871.n69 a_n20175_5871.n68 0.028
R16585 a_n20175_5871.n104 a_n20175_5871.n82 0.028
R16586 a_n20175_5871.n85 a_n20175_5871.n83 0.028
R16587 a_n20175_5871.n17 a_n20175_5871.n15 0.026
R16588 a_n20175_5871.n66 a_n20175_5871.n65 0.026
R16589 a_n20175_5871.n93 a_n20175_5871.n92 0.026
R16590 a_n20175_5871.n4 a_n20175_5871.n3 0.026
R16591 a_n20175_5871.n90 a_n20175_5871.n89 0.024
R16592 a_n20175_5871.n18 a_n20175_5871.n17 0.024
R16593 a_n20175_5871.n6 a_n20175_5871.n5 0.024
R16594 a_n20175_5871.n15 a_n20175_5871.n16 0.022
R16595 a_n20175_5871.n5 a_n20175_5871.n4 0.022
R16596 a_n20175_5871.n3 a_n20175_5871.n2 0.022
R16597 a_n20175_5871.n20 a_n20175_5871.n19 0.02
R16598 a_n20175_5871.n10 a_n20175_5871.n9 0.02
R16599 a_n20175_5871.n94 a_n20175_5871.n93 0.02
R16600 a_n20175_5871.n14 a_n20175_5871.n13 0.02
R16601 a_n20175_5871.n101 a_n20175_5871.n100 0.019
R16602 a_n20175_5871.n82 a_n20175_5871.n81 0.018
R16603 a_n20175_5871.n103 a_n20175_5871.n102 0.018
R16604 a_n20175_5871.n70 a_n20175_5871.n69 0.018
R16605 a_n20175_5871.n24 a_n20175_5871.n23 0.017
R16606 a_n20175_5871.n74 a_n20175_5871.n73 0.017
R16607 a_n20175_5871.n58 a_n20175_5871.n59 0.015
R16608 a_n20175_5871.n61 a_n20175_5871.n60 0.015
R16609 a_n20175_5871.n56 a_n20175_5871.n0 0.015
R16610 a_n20175_5871.n63 a_n20175_5871.n57 0.015
R16611 a_n20175_5871.n80 a_n20175_5871.n79 0.013
R16612 a_n20175_5871.n78 a_n20175_5871.n77 0.013
R16613 a_n20175_5871.n109 a_n20175_5871.n108 0.013
R16614 a_n20175_5871.n107 a_n20175_5871.n106 0.013
R16615 a_n20175_5871.n92 a_n20175_5871.n91 0.007
R16616 a_n20175_5871.n86 a_n20175_5871.n85 0.007
R16617 a_n20175_5871.n21 a_n20175_5871.n20 1.424
R16618 a_n20175_5871.n67 a_n20175_5871.n64 0.005
R16619 a_n20175_5871.n80 a_n20175_5871.n75 0.003
R16620 a_n20175_5871.n105 a_n20175_5871.n104 0.003
R16621 a_n20175_5871.n83 a_n20175_5871.n84 0.003
R16622 a_n20175_5871.n14 a_n20175_5871.n21 0.47
R16623 a_n17722_2897.n33 a_n17722_2897.t5 733.434
R16624 a_n17722_2897.n53 a_n17722_2897.t4 733.434
R16625 a_n17722_2897.n24 a_n17722_2897.t3 399.25
R16626 a_n17722_2897.n44 a_n17722_2897.t2 399.25
R16627 a_n17722_2897.n95 a_n17722_2897.n94 92.5
R16628 a_n17722_2897.n12 a_n17722_2897.n11 92.5
R16629 a_n17722_2897.n94 a_n17722_2897.t1 70.344
R16630 a_n17722_2897.n89 a_n17722_2897.n88 31.034
R16631 a_n17722_2897.n68 a_n17722_2897.n67 31.034
R16632 a_n17722_2897.n71 a_n17722_2897.n72 9.3
R16633 a_n17722_2897.n82 a_n17722_2897.n83 9.3
R16634 a_n17722_2897.n90 a_n17722_2897.n89 9.3
R16635 a_n17722_2897.n69 a_n17722_2897.n68 9.3
R16636 a_n17722_2897.n162 a_n17722_2897.n155 9.154
R16637 a_n17722_2897.n162 a_n17722_2897.n113 9.143
R16638 a_n17722_2897.n162 a_n17722_2897.n120 9.143
R16639 a_n17722_2897.n162 a_n17722_2897.n126 9.132
R16640 a_n17722_2897.n162 a_n17722_2897.n106 9.132
R16641 a_n17722_2897.n162 a_n17722_2897.n159 8.885
R16642 a_n17722_2897.n162 a_n17722_2897.n130 8.885
R16643 a_n17722_2897.n162 a_n17722_2897.n134 8.875
R16644 a_n17722_2897.n162 a_n17722_2897.n100 8.875
R16645 a_n17722_2897.n162 a_n17722_2897.n161 8.864
R16646 a_n17722_2897.n162 a_n17722_2897.n136 8.864
R16647 a_n17722_2897.n96 a_n17722_2897.n95 8.282
R16648 a_n17722_2897.n13 a_n17722_2897.n12 8.282
R16649 a_n17722_2897.t0 a_n17722_2897.n162 7.141
R16650 a_n17722_2897.n59 a_n17722_2897.n58 6.392
R16651 a_n17722_2897.n90 a_n17722_2897.n86 5.647
R16652 a_n17722_2897.n69 a_n17722_2897.n65 5.647
R16653 a_n17722_2897.n16 a_n17722_2897.n15 4.65
R16654 a_n17722_2897.n155 a_n17722_2897.n5 4.65
R16655 a_n17722_2897.n155 a_n17722_2897.n138 4.517
R16656 a_n17722_2897.n14 a_n17722_2897.n13 4.5
R16657 a_n17722_2897.n17 a_n17722_2897.n10 4.5
R16658 a_n17722_2897.n9 a_n17722_2897.n96 4.5
R16659 a_n17722_2897.n84 a_n17722_2897.n92 4.5
R16660 a_n17722_2897.n18 a_n17722_2897.n81 4.5
R16661 a_n17722_2897.n61 a_n17722_2897.n76 4.5
R16662 a_n17722_2897.n157 a_n17722_2897.n156 4.141
R16663 a_n17722_2897.n155 a_n17722_2897.n137 4.141
R16664 a_n17722_2897.n128 a_n17722_2897.n127 4.141
R16665 a_n17722_2897.n88 a_n17722_2897.n87 4.137
R16666 a_n17722_2897.n67 a_n17722_2897.n66 4.137
R16667 a_n17722_2897.n81 a_n17722_2897.n79 3.764
R16668 a_n17722_2897.n70 a_n17722_2897.n63 3.764
R16669 a_n17722_2897.n102 a_n17722_2897.n101 3.764
R16670 a_n17722_2897.n116 a_n17722_2897.n115 3.764
R16671 a_n17722_2897.n106 a_n17722_2897.n105 3.736
R16672 a_n17722_2897.n92 a_n17722_2897.n91 3.388
R16673 a_n17722_2897.n76 a_n17722_2897.n75 3.388
R16674 a_n17722_2897.n98 a_n17722_2897.n97 3.388
R16675 a_n17722_2897.n112 a_n17722_2897.n111 3.388
R16676 a_n17722_2897.n124 a_n17722_2897.n123 3.388
R16677 a_n17722_2897.n132 a_n17722_2897.n131 3.388
R16678 a_n17722_2897.n126 a_n17722_2897.n122 3.36
R16679 a_n17722_2897.n92 a_n17722_2897.n90 3.011
R16680 a_n17722_2897.n96 a_n17722_2897.n93 3.011
R16681 a_n17722_2897.n76 a_n17722_2897.n74 3.011
R16682 a_n17722_2897.n99 a_n17722_2897.n98 3.011
R16683 a_n17722_2897.n111 a_n17722_2897.n110 3.011
R16684 a_n17722_2897.n109 a_n17722_2897.n108 3.011
R16685 a_n17722_2897.n122 a_n17722_2897.n121 3.011
R16686 a_n17722_2897.n125 a_n17722_2897.n124 3.011
R16687 a_n17722_2897.n133 a_n17722_2897.n132 3.011
R16688 a_n17722_2897.n139 a_n17722_2897.n58 2.921
R16689 a_n17722_2897.n81 a_n17722_2897.n80 2.635
R16690 a_n17722_2897.n70 a_n17722_2897.n69 2.635
R16691 a_n17722_2897.n103 a_n17722_2897.n102 2.635
R16692 a_n17722_2897.n105 a_n17722_2897.n104 2.635
R16693 a_n17722_2897.n119 a_n17722_2897.n118 2.635
R16694 a_n17722_2897.n115 a_n17722_2897.n114 2.635
R16695 a_n17722_2897.n60 a_n17722_2897.n59 2.631
R16696 a_n17722_2897.n158 a_n17722_2897.n157 2.258
R16697 a_n17722_2897.n129 a_n17722_2897.n128 2.258
R16698 a_n17722_2897.n113 a_n17722_2897.n109 2.245
R16699 a_n17722_2897.n120 a_n17722_2897.n119 2.245
R16700 a_n17722_2897.n151 a_n17722_2897.n150 1.633
R16701 a_n17722_2897.n147 a_n17722_2897.n146 1.619
R16702 a_n17722_2897.n149 a_n17722_2897.n164 1.594
R16703 a_n17722_2897.n140 a_n17722_2897.n143 1.588
R16704 a_n17722_2897.n151 a_n17722_2897.n163 1.587
R16705 a_n17722_2897.n118 a_n17722_2897.n117 1.505
R16706 a_n17722_2897.n18 a_n17722_2897.n78 1.5
R16707 a_n17722_2897.n4 a_n17722_2897.n6 1.5
R16708 a_n17722_2897.n141 a_n17722_2897.n153 1.5
R16709 a_n17722_2897.n34 a_n17722_2897.n33 2.49
R16710 a_n17722_2897.n54 a_n17722_2897.n53 2.49
R16711 a_n17722_2897.n22 a_n17722_2897.n28 1.137
R16712 a_n17722_2897.n25 a_n17722_2897.n26 1.137
R16713 a_n17722_2897.n41 a_n17722_2897.n48 1.137
R16714 a_n17722_2897.n45 a_n17722_2897.n46 1.137
R16715 a_n17722_2897.n3 a_n17722_2897.n36 1.136
R16716 a_n17722_2897.n0 a_n17722_2897.n42 1.136
R16717 a_n17722_2897.n1 a_n17722_2897.n56 1.136
R16718 a_n17722_2897.n108 a_n17722_2897.n107 1.129
R16719 a_n17722_2897.n86 a_n17722_2897.n85 0.752
R16720 a_n17722_2897.n65 a_n17722_2897.n64 0.752
R16721 a_n17722_2897.n161 a_n17722_2897.n160 0.155
R16722 a_n17722_2897.n136 a_n17722_2897.n135 0.155
R16723 a_n17722_2897.n100 a_n17722_2897.n99 0.144
R16724 a_n17722_2897.n134 a_n17722_2897.n133 0.144
R16725 a_n17722_2897.n159 a_n17722_2897.n158 0.132
R16726 a_n17722_2897.n130 a_n17722_2897.n129 0.132
R16727 a_n17722_2897.n149 a_n17722_2897.n148 0.127
R16728 a_n17722_2897.n147 a_n17722_2897.n145 0.119
R16729 a_n17722_2897.n140 a_n17722_2897.n142 0.111
R16730 a_n17722_2897.n4 a_n17722_2897.n5 0.103
R16731 a_n17722_2897.n33 a_n17722_2897.n32 0.126
R16732 a_n17722_2897.n53 a_n17722_2897.n52 0.126
R16733 a_n17722_2897.n20 a_n17722_2897.n19 0.064
R16734 a_n17722_2897.n31 a_n17722_2897.n30 0.064
R16735 a_n17722_2897.n39 a_n17722_2897.n38 0.064
R16736 a_n17722_2897.n51 a_n17722_2897.n50 0.064
R16737 a_n17722_2897.n139 a_n17722_2897.n141 0.083
R16738 a_n17722_2897.n141 a_n17722_2897.n140 0.042
R16739 a_n17722_2897.n163 a_n17722_2897.n168 0.037
R16740 a_n17722_2897.n150 a_n17722_2897.n152 0.034
R16741 a_n17722_2897.n28 a_n17722_2897.n29 0.032
R16742 a_n17722_2897.n35 a_n17722_2897.n37 0.032
R16743 a_n17722_2897.n48 a_n17722_2897.n49 0.032
R16744 a_n17722_2897.n55 a_n17722_2897.n57 0.032
R16745 a_n17722_2897.n84 a_n17722_2897.n82 0.094
R16746 a_n17722_2897.n21 a_n17722_2897.n20 0.028
R16747 a_n17722_2897.n32 a_n17722_2897.n31 0.028
R16748 a_n17722_2897.n40 a_n17722_2897.n39 0.028
R16749 a_n17722_2897.n52 a_n17722_2897.n51 0.028
R16750 a_n17722_2897.n78 a_n17722_2897.n77 0.293
R16751 a_n17722_2897.n78 a_n17722_2897.n62 0.877
R16752 a_n17722_2897.n143 a_n17722_2897.n144 0.024
R16753 a_n17722_2897.n164 a_n17722_2897.n169 0.024
R16754 a_n17722_2897.n106 a_n17722_2897.n103 0.024
R16755 a_n17722_2897.n126 a_n17722_2897.n125 0.024
R16756 a_n17722_2897.n5 a_n17722_2897.n139 0.022
R16757 a_n17722_2897.n16 a_n17722_2897.n14 0.022
R16758 a_n17722_2897.n17 a_n17722_2897.n16 0.02
R16759 a_n17722_2897.n62 a_n17722_2897.n60 0.019
R16760 a_n17722_2897.n62 a_n17722_2897.n61 2.433
R16761 a_n17722_2897.n9 a_n17722_2897.n84 0.044
R16762 a_n17722_2897.n61 a_n17722_2897.n71 0.032
R16763 a_n17722_2897.n82 a_n17722_2897.n18 0.031
R16764 a_n17722_2897.n61 a_n17722_2897.n73 0.017
R16765 a_n17722_2897.n26 a_n17722_2897.n27 0.017
R16766 a_n17722_2897.n46 a_n17722_2897.n47 0.017
R16767 a_n17722_2897.n166 a_n17722_2897.n165 0.016
R16768 a_n17722_2897.n71 a_n17722_2897.n70 4.595
R16769 a_n17722_2897.n56 a_n17722_2897.n55 1.181
R16770 a_n17722_2897.n42 a_n17722_2897.n41 0.044
R16771 a_n17722_2897.n41 a_n17722_2897.n43 0.04
R16772 a_n17722_2897.n45 a_n17722_2897.n44 0.02
R16773 a_n17722_2897.n6 a_n17722_2897.n7 0.013
R16774 a_n17722_2897.n142 a_n17722_2897.n147 0.013
R16775 a_n17722_2897.n120 a_n17722_2897.n116 0.012
R16776 a_n17722_2897.n113 a_n17722_2897.n112 0.012
R16777 a_n17722_2897.n8 a_n17722_2897.n17 0.011
R16778 a_n17722_2897.n153 a_n17722_2897.n154 0.011
R16779 a_n17722_2897.n23 a_n17722_2897.n25 0.01
R16780 a_n17722_2897.n43 a_n17722_2897.n45 0.01
R16781 a_n17722_2897.n169 a_n17722_2897.n167 0.009
R16782 a_n17722_2897.n2 a_n17722_2897.n21 2.621
R16783 a_n17722_2897.n36 a_n17722_2897.n34 0.006
R16784 a_n17722_2897.n42 a_n17722_2897.n40 2.621
R16785 a_n17722_2897.n36 a_n17722_2897.n35 1.181
R16786 a_n17722_2897.n2 a_n17722_2897.n22 0.044
R16787 a_n17722_2897.n22 a_n17722_2897.n23 0.04
R16788 a_n17722_2897.n25 a_n17722_2897.n24 0.02
R16789 a_n17722_2897.n56 a_n17722_2897.n54 0.006
R16790 a_n17722_2897.n145 a_n17722_2897.n149 0.005
R16791 a_n17722_2897.n148 a_n17722_2897.n151 0.005
R16792 a_n17722_2897.n3 a_n17722_2897.n2 1.245
R16793 a_n17722_2897.n4 a_n17722_2897.n166 2.057
R16794 a_n17722_2897.n0 a_n17722_2897.n3 0.11
R16795 a_n17722_2897.n1 a_n17722_2897.n0 0.109
R16796 a_n17722_2897.n59 a_n17722_2897.n1 0.071
R16797 a_n17722_2897.n9 a_n17722_2897.n8 0.07
R16798 modi6.n1 modi6.t4 1037.94
R16799 modi6.n41 modi6.t5 1037.29
R16800 modi6.n1 modi6.t3 798.529
R16801 modi6.n41 modi6.t2 797.574
R16802 modi6.n276 modi6.n275 92.5
R16803 modi6.n261 modi6.n260 92.5
R16804 modi6.n275 modi6.t0 70.344
R16805 modi6.n290 modi6.n289 31.034
R16806 modi6.n230 modi6.n229 31.034
R16807 modi6.n216 modi6.n215 9.3
R16808 modi6.n291 modi6.n290 9.3
R16809 modi6.n231 modi6.n230 9.3
R16810 modi6.n238 modi6.n237 9.3
R16811 modi6.n87 modi6.n86 9.3
R16812 modi6.n176 modi6.n175 9.3
R16813 modi6.n125 modi6.n124 9.154
R16814 modi6.n277 modi6.n276 8.282
R16815 modi6.n262 modi6.n261 8.282
R16816 modi6.n124 modi6.t1 7.141
R16817 modi6.n157 modi6.n153 7.033
R16818 modi6.n46 modi6.n45 7.033
R16819 modi6.n299 modi6.n298 6.416
R16820 modi6.n291 modi6.n287 5.647
R16821 modi6.n231 modi6.n227 5.647
R16822 modi6.n269 modi6.n268 4.65
R16823 modi6.n126 modi6.n125 4.65
R16824 modi6.n244 modi6.n242 4.5
R16825 modi6.n236 modi6.n232 4.5
R16826 modi6.n254 modi6.n251 4.5
R16827 modi6.n294 modi6.n293 4.5
R16828 modi6.n280 modi6.n277 4.5
R16829 modi6.n270 modi6.n267 4.5
R16830 modi6.n263 modi6.n262 4.5
R16831 modi6.n221 modi6.n220 4.5
R16832 modi6.n204 modi6.n203 4.5
R16833 modi6.n192 modi6.n191 4.5
R16834 modi6.n182 modi6.n181 4.5
R16835 modi6.n170 modi6.n169 4.5
R16836 modi6.n163 modi6.n162 4.5
R16837 modi6.n128 modi6.n127 4.5
R16838 modi6.n122 modi6.n121 4.5
R16839 modi6.n113 modi6.n112 4.5
R16840 modi6.n106 modi6.n105 4.5
R16841 modi6.n93 modi6.n92 4.5
R16842 modi6.n63 modi6.n62 4.5
R16843 modi6.n73 modi6.n72 4.5
R16844 modi6.n62 modi6.n59 4.141
R16845 modi6.n191 modi6.n190 4.141
R16846 modi6.n289 modi6.n288 4.137
R16847 modi6.n229 modi6.n228 4.137
R16848 modi6.n300 modi6.n299 3.846
R16849 modi6.n220 modi6.n218 3.764
R16850 modi6.n232 modi6.n225 3.764
R16851 modi6.n92 modi6.n89 3.764
R16852 modi6.n169 modi6.n167 3.764
R16853 modi6.n8 modi6.n1 3.461
R16854 modi6.n293 modi6.n292 3.388
R16855 modi6.n242 modi6.n241 3.388
R16856 modi6.n72 modi6.n69 3.388
R16857 modi6.n105 modi6.n104 3.388
R16858 modi6.n181 modi6.n180 3.388
R16859 modi6.n203 modi6.n202 3.388
R16860 modi6.n293 modi6.n291 3.011
R16861 modi6.n277 modi6.n274 3.011
R16862 modi6.n242 modi6.n240 3.011
R16863 modi6.n72 modi6.n71 3.011
R16864 modi6.n105 modi6.n102 3.011
R16865 modi6.n112 modi6.n110 3.011
R16866 modi6.n175 modi6.n174 3.011
R16867 modi6.n181 modi6.n179 3.011
R16868 modi6.n203 modi6.n201 3.011
R16869 modi6.n220 modi6.n219 2.635
R16870 modi6.n251 modi6.n250 2.635
R16871 modi6.n232 modi6.n231 2.635
R16872 modi6.n92 modi6.n91 2.635
R16873 modi6.n86 modi6.n85 2.635
R16874 modi6.n162 modi6.n161 2.635
R16875 modi6.n169 modi6.n168 2.635
R16876 modi6.n62 modi6.n61 2.258
R16877 modi6.n191 modi6.n189 2.258
R16878 modi6.n299 modi6.n41 2.25
R16879 modi6.n76 modi6.n47 1.754
R16880 modi6.n249 modi6.n224 1.754
R16881 modi6.n76 modi6.n75 1.705
R16882 modi6.n151 modi6.n150 1.705
R16883 modi6.n145 modi6.n144 1.705
R16884 modi6.n139 modi6.n138 1.705
R16885 modi6.n133 modi6.n132 1.705
R16886 modi6.n116 modi6.n115 1.705
R16887 modi6.n96 modi6.n95 1.705
R16888 modi6.n82 modi6.n81 1.705
R16889 modi6.n297 modi6.n223 1.705
R16890 modi6.n296 modi6.n295 1.705
R16891 modi6.n266 modi6.n265 1.705
R16892 modi6.n249 modi6.n248 1.705
R16893 modi6.n210 modi6.n209 1.705
R16894 modi6.n301 modi6.n300 1.705
R16895 modi6.n304 modi6.n0 1.705
R16896 modi6.n162 modi6.n160 1.505
R16897 modi6.n245 modi6.n244 1.5
R16898 modi6.n248 modi6.n236 1.5
R16899 modi6.n295 modi6.n294 1.5
R16900 modi6.n281 modi6.n280 1.5
R16901 modi6.n255 modi6.n254 1.5
R16902 modi6.n271 modi6.n270 1.5
R16903 modi6.n264 modi6.n263 1.5
R16904 modi6.n222 modi6.n221 1.5
R16905 modi6.n129 modi6.n128 1.5
R16906 modi6.n123 modi6.n122 1.5
R16907 modi6.n114 modi6.n113 1.5
R16908 modi6.n107 modi6.n106 1.5
R16909 modi6.n94 modi6.n93 1.5
R16910 modi6.n14 modi6.n13 1.402
R16911 modi6.n10 modi6.n8 1.355
R16912 modi6.n298 modi6.n210 1.267
R16913 modi6.n40 modi6.n10 1.14
R16914 modi6.n15 modi6.n14 1.137
R16915 modi6.n26 modi6.n25 1.137
R16916 modi6.n20 modi6.n19 1.137
R16917 modi6.n30 modi6.n29 1.137
R16918 modi6.n37 modi6.n36 1.137
R16919 modi6.n112 modi6.n111 1.129
R16920 modi6.n209 modi6.n157 1.127
R16921 modi6.n47 modi6.n46 1.127
R16922 modi6.n205 modi6.n204 1.125
R16923 modi6.n74 modi6.n73 1.125
R16924 modi6.n287 modi6.n286 0.752
R16925 modi6.n227 modi6.n226 0.752
R16926 modi6.n298 modi6.n297 0.71
R16927 modi6.n301 modi6.n40 0.682
R16928 modi6.n45 modi6.n44 0.155
R16929 modi6.n153 modi6.n152 0.155
R16930 modi6.n71 modi6.n70 0.144
R16931 modi6.n201 modi6.n200 0.144
R16932 modi6.n61 modi6.n60 0.133
R16933 modi6.n189 modi6.n188 0.132
R16934 modi6.n216 modi6.n214 0.053
R16935 modi6.n52 modi6.n51 0.053
R16936 modi6.n67 modi6.n66 0.053
R16937 modi6.n57 modi6.n56 0.053
R16938 modi6.n176 modi6.n173 0.053
R16939 modi6.n186 modi6.n185 0.053
R16940 modi6.n196 modi6.n195 0.053
R16941 modi6.n82 modi6.n76 0.049
R16942 modi6.n96 modi6.n82 0.049
R16943 modi6.n116 modi6.n96 0.049
R16944 modi6.n133 modi6.n116 0.049
R16945 modi6.n139 modi6.n133 0.049
R16946 modi6.n145 modi6.n139 0.049
R16947 modi6.n151 modi6.n145 0.049
R16948 modi6.n210 modi6.n151 0.049
R16949 modi6.n297 modi6.n296 0.049
R16950 modi6.n296 modi6.n266 0.049
R16951 modi6.n266 modi6.n249 0.049
R16952 modi6.n8 modi6.n7 0.048
R16953 modi6.n122 modi6.n120 0.045
R16954 modi6.n163 modi6.n159 0.045
R16955 modi6.n280 modi6.n279 0.043
R16956 modi6.n263 modi6.n259 0.043
R16957 modi6.n4 modi6.n3 0.037
R16958 modi6.n195 modi6.n194 0.032
R16959 modi6.n155 modi6.n154 0.032
R16960 modi6.n222 modi6.n212 0.03
R16961 modi6.n246 modi6.n245 0.03
R16962 modi6.n68 modi6.n67 0.03
R16963 modi6.n66 modi6.n65 0.03
R16964 modi6.n185 modi6.n184 0.03
R16965 modi6.n56 modi6.n55 0.028
R16966 modi6.n197 modi6.n196 0.028
R16967 modi6.n199 modi6.n198 0.028
R16968 modi6.n53 modi6.n52 0.025
R16969 modi6.n58 modi6.n57 0.025
R16970 modi6.n128 modi6.n126 0.025
R16971 modi6.n91 modi6.n90 0.024
R16972 modi6.n179 modi6.n178 0.024
R16973 modi6.n270 modi6.n269 0.023
R16974 modi6.n187 modi6.n186 0.023
R16975 modi6.n29 modi6.n28 0.021
R16976 modi6.n221 modi6.n213 0.021
R16977 modi6.n217 modi6.n216 0.021
R16978 modi6.n234 modi6.n233 0.021
R16979 modi6.n88 modi6.n87 0.021
R16980 modi6.n170 modi6.n165 0.021
R16981 modi6.n173 modi6.n172 0.021
R16982 modi6.n283 modi6.n282 0.019
R16983 modi6.n294 modi6.n285 0.019
R16984 modi6.n235 modi6.n234 0.019
R16985 modi6.n239 modi6.n238 0.019
R16986 modi6.n244 modi6.n243 0.019
R16987 modi6.n73 modi6.n53 0.019
R16988 modi6.n100 modi6.n99 0.019
R16989 modi6.n101 modi6.n100 0.019
R16990 modi6.n172 modi6.n171 0.019
R16991 modi6.n177 modi6.n176 0.019
R16992 modi6.n183 modi6.n182 0.019
R16993 modi6.n204 modi6.n199 0.019
R16994 modi6.n46 modi6.n43 0.019
R16995 modi6.n157 modi6.n156 0.019
R16996 modi6.n36 modi6.n35 0.018
R16997 modi6.n25 modi6.n24 0.018
R16998 modi6.n95 modi6.n94 0.018
R16999 modi6.n294 modi6.n283 0.017
R17000 modi6.n244 modi6.n239 0.017
R17001 modi6.n73 modi6.n68 0.017
R17002 modi6.n64 modi6.n63 0.017
R17003 modi6.n106 modi6.n101 0.017
R17004 modi6.n113 modi6.n109 0.017
R17005 modi6.n182 modi6.n177 0.017
R17006 modi6.n193 modi6.n192 0.017
R17007 modi6.n204 modi6.n197 0.017
R17008 modi6.n7 modi6.n6 0.016
R17009 modi6.n5 modi6.n4 0.016
R17010 modi6.n3 modi6.n2 0.016
R17011 modi6.n13 modi6.n12 0.016
R17012 modi6.n295 modi6.n281 0.016
R17013 modi6.n50 modi6.n49 0.016
R17014 modi6.n78 modi6.n77 0.016
R17015 modi6.n143 modi6.n142 0.016
R17016 modi6.n149 modi6.n148 0.016
R17017 modi6.n207 modi6.n206 0.016
R17018 modi6.n221 modi6.n217 0.015
R17019 modi6.n254 modi6.n253 0.015
R17020 modi6.n236 modi6.n235 0.015
R17021 modi6.n272 modi6.n271 0.015
R17022 modi6.n256 modi6.n255 0.015
R17023 modi6.n93 modi6.n88 0.015
R17024 modi6.n164 modi6.n163 0.015
R17025 modi6.n171 modi6.n170 0.015
R17026 modi6.n114 modi6.n107 0.015
R17027 modi6.n129 modi6.n123 0.015
R17028 modi6.n135 modi6.n134 0.015
R17029 modi6.n281 modi6.n273 0.014
R17030 modi6.n264 modi6.n257 0.014
R17031 modi6.n206 modi6.n205 0.014
R17032 modi6.n74 modi6.n50 0.013
R17033 modi6.n123 modi6.n118 0.013
R17034 modi6.n130 modi6.n129 0.013
R17035 modi6.n104 modi6.n103 0.012
R17036 modi6.n167 modi6.n166 0.012
R17037 modi6.n285 modi6.n284 0.012
R17038 modi6.n253 modi6.n252 0.012
R17039 modi6.n63 modi6.n58 0.012
R17040 modi6.n109 modi6.n108 0.012
R17041 modi6.n165 modi6.n164 0.012
R17042 modi6.n192 modi6.n187 0.012
R17043 modi6.n10 modi6.n9 0.011
R17044 modi6.n36 modi6.n33 0.011
R17045 modi6.n19 modi6.n18 0.011
R17046 modi6.n14 modi6.n11 0.011
R17047 modi6.n49 modi6.n48 0.011
R17048 modi6.n79 modi6.n78 0.011
R17049 modi6.n81 modi6.n80 0.011
R17050 modi6.n107 modi6.n98 0.011
R17051 modi6.n115 modi6.n114 0.011
R17052 modi6.n148 modi6.n147 0.011
R17053 modi6.n208 modi6.n207 0.011
R17054 modi6.n35 modi6.n34 0.01
R17055 modi6.n24 modi6.n23 0.01
R17056 modi6.n248 modi6.n247 0.01
R17057 modi6.n136 modi6.n135 0.01
R17058 modi6.n32 modi6.n31 0.009
R17059 modi6.n22 modi6.n21 0.009
R17060 modi6.n138 modi6.n137 0.009
R17061 modi6.n142 modi6.n141 0.009
R17062 modi6.n150 modi6.n149 0.009
R17063 modi6.n6 modi6.n5 0.008
R17064 modi6.n279 modi6.n278 0.008
R17065 modi6.n259 modi6.n258 0.008
R17066 modi6.n223 modi6.n222 0.008
R17067 modi6.n120 modi6.n119 0.008
R17068 modi6.n159 modi6.n158 0.008
R17069 modi6.n84 modi6.n83 0.008
R17070 modi6.n94 modi6.n84 0.008
R17071 modi6.n39 modi6.n38 0.007
R17072 modi6.n30 modi6.n27 0.007
R17073 modi6.n27 modi6.n26 0.007
R17074 modi6.n17 modi6.n16 0.007
R17075 modi6.n265 modi6.n264 0.007
R17076 modi6.n247 modi6.n246 0.007
R17077 modi6.n141 modi6.n140 0.007
R17078 modi6.n31 modi6.n30 0.006
R17079 modi6.n26 modi6.n22 0.006
R17080 modi6.n212 modi6.n211 0.006
R17081 modi6.n65 modi6.n64 0.006
R17082 modi6.n55 modi6.n54 0.006
R17083 modi6.n184 modi6.n183 0.006
R17084 modi6.n194 modi6.n193 0.006
R17085 modi6.n137 modi6.n136 0.006
R17086 modi6.n75 modi6.n74 0.005
R17087 modi6.n80 modi6.n79 0.005
R17088 modi6.n98 modi6.n97 0.005
R17089 modi6.n147 modi6.n146 0.005
R17090 modi6.n209 modi6.n208 0.005
R17091 modi6.n38 modi6.n37 0.004
R17092 modi6.n20 modi6.n17 0.004
R17093 modi6.n16 modi6.n15 0.004
R17094 modi6.n43 modi6.n42 0.004
R17095 modi6.n156 modi6.n155 0.004
R17096 modi6.n302 modi6.n301 0.004
R17097 modi6.n304 modi6.n303 0.004
R17098 modi6.n305 modi6.n304 0.004
R17099 modi6.n307 modi6.n306 0.004
R17100 modi6.n308 modi6.n307 0.004
R17101 modi6 modi6.n308 0.004
R17102 modi6.n132 modi6.n131 0.003
R17103 modi6.n303 modi6.n302 0.003
R17104 modi6.n306 modi6.n305 0.003
R17105 modi6.n37 modi6.n32 0.002
R17106 modi6.n21 modi6.n20 0.002
R17107 modi6.n273 modi6.n272 0.002
R17108 modi6.n257 modi6.n256 0.002
R17109 modi6.n118 modi6.n117 0.002
R17110 modi6.n131 modi6.n130 0.002
R17111 modi6.n40 modi6.n39 0.001
R17112 modi6.n144 modi6.n143 0.001
R17113 P1 P1.t0 1038.7
R17114 P1 P1.t1 796.11
R17115 a_n5892_12356.n60 a_n5892_12356.t4 735.929
R17116 a_n5892_12356.n54 a_n5892_12356.t2 396.755
R17117 a_n5892_12356.n66 a_n5892_12356.t3 396.755
R17118 a_n5892_12356.n80 a_n5892_12356.n79 92.5
R17119 a_n5892_12356.n98 a_n5892_12356.n97 92.5
R17120 a_n5892_12356.n79 a_n5892_12356.t1 70.344
R17121 a_n5892_12356.n87 a_n5892_12356.n86 31.034
R17122 a_n5892_12356.n110 a_n5892_12356.n109 31.034
R17123 a_n5892_12356.n1 a_n5892_12356.n91 9.3
R17124 a_n5892_12356.n0 a_n5892_12356.n113 9.3
R17125 a_n5892_12356.n111 a_n5892_12356.n110 9.3
R17126 a_n5892_12356.n88 a_n5892_12356.n87 9.3
R17127 a_n5892_12356.n137 a_n5892_12356.n124 9.154
R17128 a_n5892_12356.n137 a_n5892_12356.n7 9.143
R17129 a_n5892_12356.n137 a_n5892_12356.n6 9.143
R17130 a_n5892_12356.n137 a_n5892_12356.n30 9.132
R17131 a_n5892_12356.n137 a_n5892_12356.n130 9.132
R17132 a_n5892_12356.n137 a_n5892_12356.n134 8.886
R17133 a_n5892_12356.n137 a_n5892_12356.n34 8.885
R17134 a_n5892_12356.n137 a_n5892_12356.n19 8.875
R17135 a_n5892_12356.n137 a_n5892_12356.n40 8.875
R17136 a_n5892_12356.n137 a_n5892_12356.n136 8.864
R17137 a_n5892_12356.n137 a_n5892_12356.n36 8.864
R17138 a_n5892_12356.n81 a_n5892_12356.n80 8.282
R17139 a_n5892_12356.n99 a_n5892_12356.n98 8.282
R17140 a_n5892_12356.t0 a_n5892_12356.n137 7.141
R17141 a_n5892_12356.n118 a_n5892_12356.n117 6.632
R17142 a_n5892_12356.n88 a_n5892_12356.n84 5.647
R17143 a_n5892_12356.n111 a_n5892_12356.n107 5.647
R17144 a_n5892_12356.n2 a_n5892_12356.n96 4.65
R17145 a_n5892_12356.n124 a_n5892_12356.n119 4.65
R17146 a_n5892_12356.n124 a_n5892_12356.n47 4.517
R17147 a_n5892_12356.n100 a_n5892_12356.n99 4.5
R17148 a_n5892_12356.n101 a_n5892_12356.n103 4.5
R17149 a_n5892_12356.n77 a_n5892_12356.n81 4.5
R17150 a_n5892_12356.n104 a_n5892_12356.n112 4.5
R17151 a_n5892_12356.n2 a_n5892_12356.n95 4.5
R17152 a_n5892_12356.n4 a_n5892_12356.n90 4.5
R17153 a_n5892_12356.n0 a_n5892_12356.n116 4.5
R17154 a_n5892_12356.n1 a_n5892_12356.n94 4.5
R17155 a_n5892_12356.n132 a_n5892_12356.n131 4.141
R17156 a_n5892_12356.n124 a_n5892_12356.n46 4.141
R17157 a_n5892_12356.n32 a_n5892_12356.n31 4.141
R17158 a_n5892_12356.n86 a_n5892_12356.n85 4.137
R17159 a_n5892_12356.n109 a_n5892_12356.n108 4.137
R17160 a_n5892_12356.n94 a_n5892_12356.n92 3.764
R17161 a_n5892_12356.n112 a_n5892_12356.n105 3.764
R17162 a_n5892_12356.n126 a_n5892_12356.n125 3.764
R17163 a_n5892_12356.n7 a_n5892_12356.n42 3.764
R17164 a_n5892_12356.n13 a_n5892_12356.n55 3.758
R17165 a_n5892_12356.n130 a_n5892_12356.n129 3.736
R17166 a_n5892_12356.n12 a_n5892_12356.n66 3.633
R17167 a_n5892_12356.n90 a_n5892_12356.n89 3.388
R17168 a_n5892_12356.n116 a_n5892_12356.n115 3.388
R17169 a_n5892_12356.n17 a_n5892_12356.n16 3.388
R17170 a_n5892_12356.n6 a_n5892_12356.n21 3.388
R17171 a_n5892_12356.n26 a_n5892_12356.n25 3.388
R17172 a_n5892_12356.n38 a_n5892_12356.n37 3.388
R17173 a_n5892_12356.n30 a_n5892_12356.n29 3.36
R17174 a_n5892_12356.n90 a_n5892_12356.n88 3.011
R17175 a_n5892_12356.n81 a_n5892_12356.n78 3.011
R17176 a_n5892_12356.n116 a_n5892_12356.n114 3.011
R17177 a_n5892_12356.n18 a_n5892_12356.n17 3.011
R17178 a_n5892_12356.n21 a_n5892_12356.n20 3.011
R17179 a_n5892_12356.n24 a_n5892_12356.n23 3.011
R17180 a_n5892_12356.n29 a_n5892_12356.n28 3.011
R17181 a_n5892_12356.n27 a_n5892_12356.n26 3.011
R17182 a_n5892_12356.n39 a_n5892_12356.n38 3.011
R17183 a_n5892_12356.n94 a_n5892_12356.n93 2.635
R17184 a_n5892_12356.n103 a_n5892_12356.n102 2.635
R17185 a_n5892_12356.n112 a_n5892_12356.n111 2.635
R17186 a_n5892_12356.n127 a_n5892_12356.n126 2.635
R17187 a_n5892_12356.n129 a_n5892_12356.n128 2.635
R17188 a_n5892_12356.n45 a_n5892_12356.n44 2.635
R17189 a_n5892_12356.n42 a_n5892_12356.n41 2.635
R17190 a_n5892_12356.n117 a_n5892_12356.n3 2.631
R17191 a_n5892_12356.n74 a_n5892_12356.n71 2.621
R17192 a_n5892_12356.n15 a_n5892_12356.n54 3.627
R17193 a_n5892_12356.n133 a_n5892_12356.n132 2.258
R17194 a_n5892_12356.n33 a_n5892_12356.n32 2.258
R17195 a_n5892_12356.n5 a_n5892_12356.n123 1.619
R17196 a_n5892_12356.n120 a_n5892_12356.n121 1.588
R17197 a_n5892_12356.n5 a_n5892_12356.n138 1.88
R17198 a_n5892_12356.n3 a_n5892_12356.n0 2.375
R17199 a_n5892_12356.n44 a_n5892_12356.n43 1.505
R17200 a_n5892_12356.n76 a_n5892_12356.n1 1.5
R17201 a_n5892_12356.n7 a_n5892_12356.n45 2.257
R17202 a_n5892_12356.n6 a_n5892_12356.n24 2.257
R17203 a_n5892_12356.n9 a_n5892_12356.n8 1.149
R17204 a_n5892_12356.n59 a_n5892_12356.n57 1.149
R17205 a_n5892_12356.n11 a_n5892_12356.n10 1.149
R17206 a_n5892_12356.n12 a_n5892_12356.n63 1.148
R17207 a_n5892_12356.n15 a_n5892_12356.n9 1.138
R17208 a_n5892_12356.n14 a_n5892_12356.t5 737.068
R17209 a_n5892_12356.n63 a_n5892_12356.n61 1.137
R17210 a_n5892_12356.n11 a_n5892_12356.n67 1.137
R17211 a_n5892_12356.n14 a_n5892_12356.n74 1.136
R17212 a_n5892_12356.n13 a_n5892_12356.n59 1.136
R17213 a_n5892_12356.n23 a_n5892_12356.n22 1.129
R17214 a_n5892_12356.n84 a_n5892_12356.n83 0.752
R17215 a_n5892_12356.n107 a_n5892_12356.n106 0.752
R17216 a_n5892_12356.n9 a_n5892_12356.n48 1.149
R17217 a_n5892_12356.n14 a_n5892_12356.n11 1.148
R17218 a_n5892_12356.n76 a_n5892_12356.n75 0.24
R17219 a_n5892_12356.n136 a_n5892_12356.n135 0.155
R17220 a_n5892_12356.n36 a_n5892_12356.n35 0.155
R17221 a_n5892_12356.n19 a_n5892_12356.n18 0.144
R17222 a_n5892_12356.n40 a_n5892_12356.n39 0.144
R17223 a_n5892_12356.n134 a_n5892_12356.n133 0.133
R17224 a_n5892_12356.n34 a_n5892_12356.n33 0.132
R17225 a_n5892_12356.n54 a_n5892_12356.n52 0.126
R17226 a_n5892_12356.n66 a_n5892_12356.n64 0.126
R17227 a_n5892_12356.n13 a_n5892_12356.n15 0.114
R17228 a_n5892_12356.n14 a_n5892_12356.n12 0.11
R17229 a_n5892_12356.n12 a_n5892_12356.n13 0.107
R17230 a_n5892_12356.n101 a_n5892_12356.n100 0.082
R17231 a_n5892_12356.n77 a_n5892_12356.n82 0.071
R17232 a_n5892_12356.n104 a_n5892_12356.n101 0.042
R17233 a_n5892_12356.n59 a_n5892_12356.n60 0.059
R17234 a_n5892_12356.n8 a_n5892_12356.n50 0.032
R17235 a_n5892_12356.n10 a_n5892_12356.n69 0.032
R17236 a_n5892_12356.n52 a_n5892_12356.n53 0.028
R17237 a_n5892_12356.n48 a_n5892_12356.n49 0.028
R17238 a_n5892_12356.n8 a_n5892_12356.n51 0.028
R17239 a_n5892_12356.n55 a_n5892_12356.n56 0.028
R17240 a_n5892_12356.n57 a_n5892_12356.n58 0.028
R17241 a_n5892_12356.n64 a_n5892_12356.n65 0.028
R17242 a_n5892_12356.n61 a_n5892_12356.n62 0.028
R17243 a_n5892_12356.n71 a_n5892_12356.n72 0.028
R17244 a_n5892_12356.n67 a_n5892_12356.n68 0.028
R17245 a_n5892_12356.n10 a_n5892_12356.n70 0.028
R17246 a_n5892_12356.n74 a_n5892_12356.n73 0.027
R17247 a_n5892_12356.n121 a_n5892_12356.n122 0.024
R17248 a_n5892_12356.n30 a_n5892_12356.n27 0.024
R17249 a_n5892_12356.n130 a_n5892_12356.n127 0.024
R17250 a_n5892_12356.n119 a_n5892_12356.n120 0.147
R17251 a_n5892_12356.n120 a_n5892_12356.n5 0.124
R17252 a_n5892_12356.n117 a_n5892_12356.n14 0.072
R17253 a_n5892_12356.n119 a_n5892_12356.n118 2.702
R17254 a_n5892_12356.n3 a_n5892_12356.n76 0.955
R17255 a_n5892_12356.n0 a_n5892_12356.n104 0.127
R17256 a_n5892_12356.n1 a_n5892_12356.n4 0.11
R17257 a_n5892_12356.n4 a_n5892_12356.n77 0.058
R17258 a_n5892_12356.n100 a_n5892_12356.n2 0.042
R17259 a_n11858_2898.n33 a_n11858_2898.t2 733.434
R17260 a_n11858_2898.n53 a_n11858_2898.t5 733.434
R17261 a_n11858_2898.n24 a_n11858_2898.t3 399.25
R17262 a_n11858_2898.n44 a_n11858_2898.t4 399.25
R17263 a_n11858_2898.n95 a_n11858_2898.n94 92.5
R17264 a_n11858_2898.n12 a_n11858_2898.n11 92.5
R17265 a_n11858_2898.n94 a_n11858_2898.t1 70.344
R17266 a_n11858_2898.n89 a_n11858_2898.n88 31.034
R17267 a_n11858_2898.n68 a_n11858_2898.n67 31.034
R17268 a_n11858_2898.n71 a_n11858_2898.n72 9.3
R17269 a_n11858_2898.n82 a_n11858_2898.n83 9.3
R17270 a_n11858_2898.n90 a_n11858_2898.n89 9.3
R17271 a_n11858_2898.n69 a_n11858_2898.n68 9.3
R17272 a_n11858_2898.n162 a_n11858_2898.n155 9.154
R17273 a_n11858_2898.n162 a_n11858_2898.n113 9.143
R17274 a_n11858_2898.n162 a_n11858_2898.n120 9.143
R17275 a_n11858_2898.n162 a_n11858_2898.n126 9.132
R17276 a_n11858_2898.n162 a_n11858_2898.n106 9.132
R17277 a_n11858_2898.n162 a_n11858_2898.n159 8.885
R17278 a_n11858_2898.n162 a_n11858_2898.n130 8.885
R17279 a_n11858_2898.n162 a_n11858_2898.n134 8.875
R17280 a_n11858_2898.n162 a_n11858_2898.n100 8.875
R17281 a_n11858_2898.n162 a_n11858_2898.n161 8.864
R17282 a_n11858_2898.n162 a_n11858_2898.n136 8.864
R17283 a_n11858_2898.n96 a_n11858_2898.n95 8.282
R17284 a_n11858_2898.n13 a_n11858_2898.n12 8.282
R17285 a_n11858_2898.t0 a_n11858_2898.n162 7.141
R17286 a_n11858_2898.n59 a_n11858_2898.n58 6.381
R17287 a_n11858_2898.n90 a_n11858_2898.n86 5.647
R17288 a_n11858_2898.n69 a_n11858_2898.n65 5.647
R17289 a_n11858_2898.n16 a_n11858_2898.n15 4.65
R17290 a_n11858_2898.n155 a_n11858_2898.n5 4.65
R17291 a_n11858_2898.n155 a_n11858_2898.n138 4.517
R17292 a_n11858_2898.n14 a_n11858_2898.n13 4.5
R17293 a_n11858_2898.n17 a_n11858_2898.n10 4.5
R17294 a_n11858_2898.n9 a_n11858_2898.n96 4.5
R17295 a_n11858_2898.n84 a_n11858_2898.n92 4.5
R17296 a_n11858_2898.n18 a_n11858_2898.n81 4.5
R17297 a_n11858_2898.n61 a_n11858_2898.n76 4.5
R17298 a_n11858_2898.n157 a_n11858_2898.n156 4.141
R17299 a_n11858_2898.n155 a_n11858_2898.n137 4.141
R17300 a_n11858_2898.n128 a_n11858_2898.n127 4.141
R17301 a_n11858_2898.n88 a_n11858_2898.n87 4.137
R17302 a_n11858_2898.n67 a_n11858_2898.n66 4.137
R17303 a_n11858_2898.n81 a_n11858_2898.n79 3.764
R17304 a_n11858_2898.n70 a_n11858_2898.n63 3.764
R17305 a_n11858_2898.n102 a_n11858_2898.n101 3.764
R17306 a_n11858_2898.n116 a_n11858_2898.n115 3.764
R17307 a_n11858_2898.n106 a_n11858_2898.n105 3.736
R17308 a_n11858_2898.n92 a_n11858_2898.n91 3.388
R17309 a_n11858_2898.n76 a_n11858_2898.n75 3.388
R17310 a_n11858_2898.n98 a_n11858_2898.n97 3.388
R17311 a_n11858_2898.n112 a_n11858_2898.n111 3.388
R17312 a_n11858_2898.n124 a_n11858_2898.n123 3.388
R17313 a_n11858_2898.n132 a_n11858_2898.n131 3.388
R17314 a_n11858_2898.n126 a_n11858_2898.n122 3.36
R17315 a_n11858_2898.n92 a_n11858_2898.n90 3.011
R17316 a_n11858_2898.n96 a_n11858_2898.n93 3.011
R17317 a_n11858_2898.n76 a_n11858_2898.n74 3.011
R17318 a_n11858_2898.n99 a_n11858_2898.n98 3.011
R17319 a_n11858_2898.n111 a_n11858_2898.n110 3.011
R17320 a_n11858_2898.n109 a_n11858_2898.n108 3.011
R17321 a_n11858_2898.n122 a_n11858_2898.n121 3.011
R17322 a_n11858_2898.n125 a_n11858_2898.n124 3.011
R17323 a_n11858_2898.n133 a_n11858_2898.n132 3.011
R17324 a_n11858_2898.n139 a_n11858_2898.n58 2.921
R17325 a_n11858_2898.n81 a_n11858_2898.n80 2.635
R17326 a_n11858_2898.n70 a_n11858_2898.n69 2.635
R17327 a_n11858_2898.n103 a_n11858_2898.n102 2.635
R17328 a_n11858_2898.n105 a_n11858_2898.n104 2.635
R17329 a_n11858_2898.n119 a_n11858_2898.n118 2.635
R17330 a_n11858_2898.n115 a_n11858_2898.n114 2.635
R17331 a_n11858_2898.n60 a_n11858_2898.n59 2.632
R17332 a_n11858_2898.n158 a_n11858_2898.n157 2.258
R17333 a_n11858_2898.n129 a_n11858_2898.n128 2.258
R17334 a_n11858_2898.n113 a_n11858_2898.n109 2.245
R17335 a_n11858_2898.n120 a_n11858_2898.n119 2.245
R17336 a_n11858_2898.n151 a_n11858_2898.n150 1.633
R17337 a_n11858_2898.n147 a_n11858_2898.n146 1.619
R17338 a_n11858_2898.n149 a_n11858_2898.n164 1.594
R17339 a_n11858_2898.n140 a_n11858_2898.n143 1.588
R17340 a_n11858_2898.n151 a_n11858_2898.n163 1.587
R17341 a_n11858_2898.n118 a_n11858_2898.n117 1.505
R17342 a_n11858_2898.n18 a_n11858_2898.n78 1.5
R17343 a_n11858_2898.n4 a_n11858_2898.n6 1.5
R17344 a_n11858_2898.n141 a_n11858_2898.n153 1.5
R17345 a_n11858_2898.n34 a_n11858_2898.n33 2.49
R17346 a_n11858_2898.n54 a_n11858_2898.n53 2.49
R17347 a_n11858_2898.n22 a_n11858_2898.n28 1.137
R17348 a_n11858_2898.n25 a_n11858_2898.n26 1.137
R17349 a_n11858_2898.n41 a_n11858_2898.n48 1.137
R17350 a_n11858_2898.n45 a_n11858_2898.n46 1.137
R17351 a_n11858_2898.n3 a_n11858_2898.n36 1.136
R17352 a_n11858_2898.n0 a_n11858_2898.n42 1.136
R17353 a_n11858_2898.n1 a_n11858_2898.n56 1.136
R17354 a_n11858_2898.n108 a_n11858_2898.n107 1.129
R17355 a_n11858_2898.n86 a_n11858_2898.n85 0.752
R17356 a_n11858_2898.n65 a_n11858_2898.n64 0.752
R17357 a_n11858_2898.n161 a_n11858_2898.n160 0.155
R17358 a_n11858_2898.n136 a_n11858_2898.n135 0.155
R17359 a_n11858_2898.n100 a_n11858_2898.n99 0.144
R17360 a_n11858_2898.n134 a_n11858_2898.n133 0.144
R17361 a_n11858_2898.n159 a_n11858_2898.n158 0.132
R17362 a_n11858_2898.n130 a_n11858_2898.n129 0.132
R17363 a_n11858_2898.n149 a_n11858_2898.n148 0.127
R17364 a_n11858_2898.n147 a_n11858_2898.n145 0.119
R17365 a_n11858_2898.n140 a_n11858_2898.n142 0.111
R17366 a_n11858_2898.n4 a_n11858_2898.n5 0.103
R17367 a_n11858_2898.n33 a_n11858_2898.n32 0.126
R17368 a_n11858_2898.n53 a_n11858_2898.n52 0.126
R17369 a_n11858_2898.n20 a_n11858_2898.n19 0.064
R17370 a_n11858_2898.n31 a_n11858_2898.n30 0.064
R17371 a_n11858_2898.n39 a_n11858_2898.n38 0.064
R17372 a_n11858_2898.n51 a_n11858_2898.n50 0.064
R17373 a_n11858_2898.n139 a_n11858_2898.n141 0.083
R17374 a_n11858_2898.n141 a_n11858_2898.n140 0.042
R17375 a_n11858_2898.n163 a_n11858_2898.n168 0.037
R17376 a_n11858_2898.n150 a_n11858_2898.n152 0.034
R17377 a_n11858_2898.n28 a_n11858_2898.n29 0.032
R17378 a_n11858_2898.n35 a_n11858_2898.n37 0.032
R17379 a_n11858_2898.n48 a_n11858_2898.n49 0.032
R17380 a_n11858_2898.n55 a_n11858_2898.n57 0.032
R17381 a_n11858_2898.n84 a_n11858_2898.n82 0.094
R17382 a_n11858_2898.n21 a_n11858_2898.n20 0.028
R17383 a_n11858_2898.n32 a_n11858_2898.n31 0.028
R17384 a_n11858_2898.n40 a_n11858_2898.n39 0.028
R17385 a_n11858_2898.n52 a_n11858_2898.n51 0.028
R17386 a_n11858_2898.n78 a_n11858_2898.n77 0.293
R17387 a_n11858_2898.n78 a_n11858_2898.n62 0.877
R17388 a_n11858_2898.n143 a_n11858_2898.n144 0.024
R17389 a_n11858_2898.n164 a_n11858_2898.n169 0.024
R17390 a_n11858_2898.n106 a_n11858_2898.n103 0.024
R17391 a_n11858_2898.n126 a_n11858_2898.n125 0.024
R17392 a_n11858_2898.n5 a_n11858_2898.n139 0.022
R17393 a_n11858_2898.n16 a_n11858_2898.n14 0.022
R17394 a_n11858_2898.n17 a_n11858_2898.n16 0.02
R17395 a_n11858_2898.n62 a_n11858_2898.n60 0.019
R17396 a_n11858_2898.n62 a_n11858_2898.n61 2.433
R17397 a_n11858_2898.n9 a_n11858_2898.n84 0.044
R17398 a_n11858_2898.n61 a_n11858_2898.n71 0.032
R17399 a_n11858_2898.n82 a_n11858_2898.n18 0.031
R17400 a_n11858_2898.n61 a_n11858_2898.n73 0.017
R17401 a_n11858_2898.n26 a_n11858_2898.n27 0.017
R17402 a_n11858_2898.n46 a_n11858_2898.n47 0.017
R17403 a_n11858_2898.n166 a_n11858_2898.n165 0.016
R17404 a_n11858_2898.n71 a_n11858_2898.n70 4.595
R17405 a_n11858_2898.n56 a_n11858_2898.n55 1.181
R17406 a_n11858_2898.n42 a_n11858_2898.n41 0.044
R17407 a_n11858_2898.n41 a_n11858_2898.n43 0.04
R17408 a_n11858_2898.n45 a_n11858_2898.n44 0.02
R17409 a_n11858_2898.n6 a_n11858_2898.n7 0.013
R17410 a_n11858_2898.n142 a_n11858_2898.n147 0.013
R17411 a_n11858_2898.n120 a_n11858_2898.n116 0.012
R17412 a_n11858_2898.n113 a_n11858_2898.n112 0.012
R17413 a_n11858_2898.n8 a_n11858_2898.n17 0.011
R17414 a_n11858_2898.n153 a_n11858_2898.n154 0.011
R17415 a_n11858_2898.n23 a_n11858_2898.n25 0.01
R17416 a_n11858_2898.n43 a_n11858_2898.n45 0.01
R17417 a_n11858_2898.n169 a_n11858_2898.n167 0.009
R17418 a_n11858_2898.n2 a_n11858_2898.n21 2.621
R17419 a_n11858_2898.n36 a_n11858_2898.n34 0.006
R17420 a_n11858_2898.n42 a_n11858_2898.n40 2.621
R17421 a_n11858_2898.n36 a_n11858_2898.n35 1.181
R17422 a_n11858_2898.n2 a_n11858_2898.n22 0.044
R17423 a_n11858_2898.n22 a_n11858_2898.n23 0.04
R17424 a_n11858_2898.n25 a_n11858_2898.n24 0.02
R17425 a_n11858_2898.n56 a_n11858_2898.n54 0.006
R17426 a_n11858_2898.n145 a_n11858_2898.n149 0.005
R17427 a_n11858_2898.n148 a_n11858_2898.n151 0.005
R17428 a_n11858_2898.n3 a_n11858_2898.n2 1.245
R17429 a_n11858_2898.n4 a_n11858_2898.n166 2.057
R17430 a_n11858_2898.n0 a_n11858_2898.n3 0.11
R17431 a_n11858_2898.n1 a_n11858_2898.n0 0.109
R17432 a_n11858_2898.n59 a_n11858_2898.n1 0.071
R17433 a_n11858_2898.n9 a_n11858_2898.n8 0.07
R17434 a_n23475_2903.n33 a_n23475_2903.t5 733.436
R17435 a_n23475_2903.n53 a_n23475_2903.t3 733.436
R17436 a_n23475_2903.n24 a_n23475_2903.t4 399.248
R17437 a_n23475_2903.n44 a_n23475_2903.t2 399.248
R17438 a_n23475_2903.n95 a_n23475_2903.n94 92.5
R17439 a_n23475_2903.n12 a_n23475_2903.n11 92.5
R17440 a_n23475_2903.n94 a_n23475_2903.t1 70.344
R17441 a_n23475_2903.n89 a_n23475_2903.n88 31.034
R17442 a_n23475_2903.n68 a_n23475_2903.n67 31.034
R17443 a_n23475_2903.n71 a_n23475_2903.n72 9.3
R17444 a_n23475_2903.n82 a_n23475_2903.n83 9.3
R17445 a_n23475_2903.n90 a_n23475_2903.n89 9.3
R17446 a_n23475_2903.n69 a_n23475_2903.n68 9.3
R17447 a_n23475_2903.n162 a_n23475_2903.n155 9.154
R17448 a_n23475_2903.n162 a_n23475_2903.n113 9.143
R17449 a_n23475_2903.n162 a_n23475_2903.n120 9.143
R17450 a_n23475_2903.n162 a_n23475_2903.n126 9.132
R17451 a_n23475_2903.n162 a_n23475_2903.n106 9.132
R17452 a_n23475_2903.n162 a_n23475_2903.n159 8.885
R17453 a_n23475_2903.n162 a_n23475_2903.n130 8.885
R17454 a_n23475_2903.n162 a_n23475_2903.n134 8.875
R17455 a_n23475_2903.n162 a_n23475_2903.n100 8.875
R17456 a_n23475_2903.n162 a_n23475_2903.n161 8.864
R17457 a_n23475_2903.n162 a_n23475_2903.n136 8.864
R17458 a_n23475_2903.n96 a_n23475_2903.n95 8.282
R17459 a_n23475_2903.n13 a_n23475_2903.n12 8.282
R17460 a_n23475_2903.t0 a_n23475_2903.n162 7.141
R17461 a_n23475_2903.n59 a_n23475_2903.n58 6.381
R17462 a_n23475_2903.n90 a_n23475_2903.n86 5.647
R17463 a_n23475_2903.n69 a_n23475_2903.n65 5.647
R17464 a_n23475_2903.n16 a_n23475_2903.n15 4.65
R17465 a_n23475_2903.n155 a_n23475_2903.n5 4.65
R17466 a_n23475_2903.n155 a_n23475_2903.n138 4.517
R17467 a_n23475_2903.n14 a_n23475_2903.n13 4.5
R17468 a_n23475_2903.n17 a_n23475_2903.n10 4.5
R17469 a_n23475_2903.n9 a_n23475_2903.n96 4.5
R17470 a_n23475_2903.n84 a_n23475_2903.n92 4.5
R17471 a_n23475_2903.n18 a_n23475_2903.n81 4.5
R17472 a_n23475_2903.n61 a_n23475_2903.n76 4.5
R17473 a_n23475_2903.n157 a_n23475_2903.n156 4.141
R17474 a_n23475_2903.n155 a_n23475_2903.n137 4.141
R17475 a_n23475_2903.n128 a_n23475_2903.n127 4.141
R17476 a_n23475_2903.n88 a_n23475_2903.n87 4.137
R17477 a_n23475_2903.n67 a_n23475_2903.n66 4.137
R17478 a_n23475_2903.n81 a_n23475_2903.n79 3.764
R17479 a_n23475_2903.n70 a_n23475_2903.n63 3.764
R17480 a_n23475_2903.n102 a_n23475_2903.n101 3.764
R17481 a_n23475_2903.n116 a_n23475_2903.n115 3.764
R17482 a_n23475_2903.n106 a_n23475_2903.n105 3.736
R17483 a_n23475_2903.n92 a_n23475_2903.n91 3.388
R17484 a_n23475_2903.n76 a_n23475_2903.n75 3.388
R17485 a_n23475_2903.n98 a_n23475_2903.n97 3.388
R17486 a_n23475_2903.n112 a_n23475_2903.n111 3.388
R17487 a_n23475_2903.n124 a_n23475_2903.n123 3.388
R17488 a_n23475_2903.n132 a_n23475_2903.n131 3.388
R17489 a_n23475_2903.n126 a_n23475_2903.n122 3.36
R17490 a_n23475_2903.n92 a_n23475_2903.n90 3.011
R17491 a_n23475_2903.n96 a_n23475_2903.n93 3.011
R17492 a_n23475_2903.n76 a_n23475_2903.n74 3.011
R17493 a_n23475_2903.n99 a_n23475_2903.n98 3.011
R17494 a_n23475_2903.n111 a_n23475_2903.n110 3.011
R17495 a_n23475_2903.n109 a_n23475_2903.n108 3.011
R17496 a_n23475_2903.n122 a_n23475_2903.n121 3.011
R17497 a_n23475_2903.n125 a_n23475_2903.n124 3.011
R17498 a_n23475_2903.n133 a_n23475_2903.n132 3.011
R17499 a_n23475_2903.n139 a_n23475_2903.n58 2.921
R17500 a_n23475_2903.n81 a_n23475_2903.n80 2.635
R17501 a_n23475_2903.n70 a_n23475_2903.n69 2.635
R17502 a_n23475_2903.n103 a_n23475_2903.n102 2.635
R17503 a_n23475_2903.n105 a_n23475_2903.n104 2.635
R17504 a_n23475_2903.n119 a_n23475_2903.n118 2.635
R17505 a_n23475_2903.n115 a_n23475_2903.n114 2.635
R17506 a_n23475_2903.n60 a_n23475_2903.n59 2.63
R17507 a_n23475_2903.n158 a_n23475_2903.n157 2.258
R17508 a_n23475_2903.n129 a_n23475_2903.n128 2.258
R17509 a_n23475_2903.n113 a_n23475_2903.n109 2.245
R17510 a_n23475_2903.n120 a_n23475_2903.n119 2.245
R17511 a_n23475_2903.n151 a_n23475_2903.n150 1.633
R17512 a_n23475_2903.n147 a_n23475_2903.n146 1.619
R17513 a_n23475_2903.n149 a_n23475_2903.n164 1.594
R17514 a_n23475_2903.n140 a_n23475_2903.n143 1.588
R17515 a_n23475_2903.n151 a_n23475_2903.n163 1.587
R17516 a_n23475_2903.n118 a_n23475_2903.n117 1.505
R17517 a_n23475_2903.n18 a_n23475_2903.n78 1.5
R17518 a_n23475_2903.n4 a_n23475_2903.n6 1.5
R17519 a_n23475_2903.n141 a_n23475_2903.n153 1.5
R17520 a_n23475_2903.n34 a_n23475_2903.n33 2.49
R17521 a_n23475_2903.n54 a_n23475_2903.n53 2.49
R17522 a_n23475_2903.n22 a_n23475_2903.n28 1.137
R17523 a_n23475_2903.n25 a_n23475_2903.n26 1.137
R17524 a_n23475_2903.n41 a_n23475_2903.n48 1.137
R17525 a_n23475_2903.n45 a_n23475_2903.n46 1.137
R17526 a_n23475_2903.n3 a_n23475_2903.n36 1.136
R17527 a_n23475_2903.n0 a_n23475_2903.n42 1.136
R17528 a_n23475_2903.n1 a_n23475_2903.n56 1.136
R17529 a_n23475_2903.n108 a_n23475_2903.n107 1.129
R17530 a_n23475_2903.n86 a_n23475_2903.n85 0.752
R17531 a_n23475_2903.n65 a_n23475_2903.n64 0.752
R17532 a_n23475_2903.n161 a_n23475_2903.n160 0.155
R17533 a_n23475_2903.n136 a_n23475_2903.n135 0.155
R17534 a_n23475_2903.n100 a_n23475_2903.n99 0.144
R17535 a_n23475_2903.n134 a_n23475_2903.n133 0.144
R17536 a_n23475_2903.n159 a_n23475_2903.n158 0.132
R17537 a_n23475_2903.n130 a_n23475_2903.n129 0.132
R17538 a_n23475_2903.n149 a_n23475_2903.n148 0.127
R17539 a_n23475_2903.n147 a_n23475_2903.n145 0.119
R17540 a_n23475_2903.n140 a_n23475_2903.n142 0.111
R17541 a_n23475_2903.n4 a_n23475_2903.n5 0.103
R17542 a_n23475_2903.n33 a_n23475_2903.n32 0.126
R17543 a_n23475_2903.n53 a_n23475_2903.n52 0.126
R17544 a_n23475_2903.n20 a_n23475_2903.n19 0.064
R17545 a_n23475_2903.n31 a_n23475_2903.n30 0.064
R17546 a_n23475_2903.n39 a_n23475_2903.n38 0.064
R17547 a_n23475_2903.n51 a_n23475_2903.n50 0.064
R17548 a_n23475_2903.n139 a_n23475_2903.n141 0.083
R17549 a_n23475_2903.n141 a_n23475_2903.n140 0.042
R17550 a_n23475_2903.n163 a_n23475_2903.n168 0.037
R17551 a_n23475_2903.n150 a_n23475_2903.n152 0.034
R17552 a_n23475_2903.n28 a_n23475_2903.n29 0.032
R17553 a_n23475_2903.n35 a_n23475_2903.n37 0.032
R17554 a_n23475_2903.n48 a_n23475_2903.n49 0.032
R17555 a_n23475_2903.n55 a_n23475_2903.n57 0.032
R17556 a_n23475_2903.n84 a_n23475_2903.n82 0.094
R17557 a_n23475_2903.n21 a_n23475_2903.n20 0.028
R17558 a_n23475_2903.n32 a_n23475_2903.n31 0.028
R17559 a_n23475_2903.n40 a_n23475_2903.n39 0.028
R17560 a_n23475_2903.n52 a_n23475_2903.n51 0.028
R17561 a_n23475_2903.n78 a_n23475_2903.n77 0.293
R17562 a_n23475_2903.n78 a_n23475_2903.n62 0.877
R17563 a_n23475_2903.n143 a_n23475_2903.n144 0.024
R17564 a_n23475_2903.n164 a_n23475_2903.n169 0.024
R17565 a_n23475_2903.n106 a_n23475_2903.n103 0.024
R17566 a_n23475_2903.n126 a_n23475_2903.n125 0.024
R17567 a_n23475_2903.n5 a_n23475_2903.n139 0.022
R17568 a_n23475_2903.n16 a_n23475_2903.n14 0.022
R17569 a_n23475_2903.n17 a_n23475_2903.n16 0.02
R17570 a_n23475_2903.n62 a_n23475_2903.n60 0.019
R17571 a_n23475_2903.n62 a_n23475_2903.n61 2.433
R17572 a_n23475_2903.n9 a_n23475_2903.n84 0.044
R17573 a_n23475_2903.n61 a_n23475_2903.n71 0.032
R17574 a_n23475_2903.n82 a_n23475_2903.n18 0.031
R17575 a_n23475_2903.n61 a_n23475_2903.n73 0.017
R17576 a_n23475_2903.n26 a_n23475_2903.n27 0.017
R17577 a_n23475_2903.n46 a_n23475_2903.n47 0.017
R17578 a_n23475_2903.n166 a_n23475_2903.n165 0.016
R17579 a_n23475_2903.n71 a_n23475_2903.n70 4.595
R17580 a_n23475_2903.n56 a_n23475_2903.n55 1.181
R17581 a_n23475_2903.n42 a_n23475_2903.n41 0.044
R17582 a_n23475_2903.n41 a_n23475_2903.n43 0.04
R17583 a_n23475_2903.n45 a_n23475_2903.n44 0.02
R17584 a_n23475_2903.n6 a_n23475_2903.n7 0.013
R17585 a_n23475_2903.n142 a_n23475_2903.n147 0.013
R17586 a_n23475_2903.n120 a_n23475_2903.n116 0.012
R17587 a_n23475_2903.n113 a_n23475_2903.n112 0.012
R17588 a_n23475_2903.n8 a_n23475_2903.n17 0.011
R17589 a_n23475_2903.n153 a_n23475_2903.n154 0.011
R17590 a_n23475_2903.n23 a_n23475_2903.n25 0.01
R17591 a_n23475_2903.n43 a_n23475_2903.n45 0.01
R17592 a_n23475_2903.n169 a_n23475_2903.n167 0.009
R17593 a_n23475_2903.n2 a_n23475_2903.n21 2.621
R17594 a_n23475_2903.n36 a_n23475_2903.n34 0.006
R17595 a_n23475_2903.n42 a_n23475_2903.n40 2.621
R17596 a_n23475_2903.n36 a_n23475_2903.n35 1.181
R17597 a_n23475_2903.n2 a_n23475_2903.n22 0.044
R17598 a_n23475_2903.n22 a_n23475_2903.n23 0.04
R17599 a_n23475_2903.n25 a_n23475_2903.n24 0.02
R17600 a_n23475_2903.n56 a_n23475_2903.n54 0.006
R17601 a_n23475_2903.n145 a_n23475_2903.n149 0.005
R17602 a_n23475_2903.n148 a_n23475_2903.n151 0.005
R17603 a_n23475_2903.n3 a_n23475_2903.n2 1.245
R17604 a_n23475_2903.n4 a_n23475_2903.n166 2.057
R17605 a_n23475_2903.n0 a_n23475_2903.n3 0.11
R17606 a_n23475_2903.n1 a_n23475_2903.n0 0.109
R17607 a_n23475_2903.n59 a_n23475_2903.n1 0.072
R17608 a_n23475_2903.n9 a_n23475_2903.n8 0.07
R17609 a_n2702_5867.n97 a_n2702_5867.t5 1040.33
R17610 a_n2702_5867.n97 a_n2702_5867.t4 794.533
R17611 a_n2702_5867.n41 a_n2702_5867.n40 13.176
R17612 a_n2702_5867.n95 a_n2702_5867.t3 11.614
R17613 a_n2702_5867.n95 a_n2702_5867.t0 11.298
R17614 a_n2702_5867.n96 a_n2702_5867.t2 10.376
R17615 a_n2702_5867.n151 a_n2702_5867.n34 9.3
R17616 a_n2702_5867.n151 a_n2702_5867.n142 9.3
R17617 a_n2702_5867.n151 a_n2702_5867.n136 9.3
R17618 a_n2702_5867.n151 a_n2702_5867.n49 9.3
R17619 a_n2702_5867.n151 a_n2702_5867.n54 9.3
R17620 a_n2702_5867.n151 a_n2702_5867.n124 9.3
R17621 a_n2702_5867.n151 a_n2702_5867.n150 8.469
R17622 a_n2702_5867.n151 a_n2702_5867.n114 8.469
R17623 a_n2702_5867.n151 a_n2702_5867.n119 8.125
R17624 a_n2702_5867.n151 a_n2702_5867.n29 8.124
R17625 a_n2702_5867.n151 a_n2702_5867.n111 8.097
R17626 a_n2702_5867.n151 a_n2702_5867.n147 8.096
R17627 a_n2702_5867.n151 a_n2702_5867.n127 8.016
R17628 a_n2702_5867.n151 a_n2702_5867.n39 8.016
R17629 a_n2702_5867.n151 a_n2702_5867.n131 7.964
R17630 a_n2702_5867.n151 a_n2702_5867.n44 7.964
R17631 a_n2702_5867.n126 a_n2702_5867.n125 6.4
R17632 a_n2702_5867.n110 a_n2702_5867.n55 6.4
R17633 a_n2702_5867.n145 a_n2702_5867.n144 6.023
R17634 a_n2702_5867.n37 a_n2702_5867.n36 6.023
R17635 a_n2702_5867.n136 a_n2702_5867.n135 6.023
R17636 a_n2702_5867.n43 a_n2702_5867.n42 6.023
R17637 a_n2702_5867.n130 a_n2702_5867.n129 6.023
R17638 a_n2702_5867.n149 a_n2702_5867.n148 5.647
R17639 a_n2702_5867.n49 a_n2702_5867.n46 5.647
R17640 a_n2702_5867.n117 a_n2702_5867.n116 5.647
R17641 a_n2702_5867.n113 a_n2702_5867.n112 5.647
R17642 a_n2702_5867.n133 a_n2702_5867.n132 5.457
R17643 a_n2702_5867.n27 a_n2702_5867.n26 5.27
R17644 a_n2702_5867.n48 a_n2702_5867.n47 5.08
R17645 a_n2702_5867.n34 a_n2702_5867.n33 4.517
R17646 a_n2702_5867.n124 a_n2702_5867.n121 4.517
R17647 a_n2702_5867.n63 a_n2702_5867.n62 4.5
R17648 a_n2702_5867.n2 a_n2702_5867.n1 4.5
R17649 a_n2702_5867.n31 a_n2702_5867.n30 4.314
R17650 a_n2702_5867.n141 a_n2702_5867.n140 4.141
R17651 a_n2702_5867.n51 a_n2702_5867.n50 4.141
R17652 a_n2702_5867.n138 a_n2702_5867.n137 3.944
R17653 a_n2702_5867.n123 a_n2702_5867.n122 3.937
R17654 a_n2702_5867.n53 a_n2702_5867.n52 3.567
R17655 a_n2702_5867.n98 a_n2702_5867.n97 3.395
R17656 a_n2702_5867.n110 a_n2702_5867.n109 3.033
R17657 a_n2702_5867.t1 a_n2702_5867.n151 2.9
R17658 a_n2702_5867.n142 a_n2702_5867.n141 2.258
R17659 a_n2702_5867.n54 a_n2702_5867.n51 2.258
R17660 a_n2702_5867.n99 a_n2702_5867.n98 2.168
R17661 a_n2702_5867.n33 a_n2702_5867.n32 1.882
R17662 a_n2702_5867.n121 a_n2702_5867.n120 1.882
R17663 a_n2702_5867.n54 a_n2702_5867.n53 1.505
R17664 a_n2702_5867.n82 a_n2702_5867.n103 1.5
R17665 a_n2702_5867.n64 a_n2702_5867.n66 1.5
R17666 a_n2702_5867.n63 a_n2702_5867.n61 1.5
R17667 a_n2702_5867.n21 a_n2702_5867.n24 1.5
R17668 a_n2702_5867.n12 a_n2702_5867.n11 1.5
R17669 a_n2702_5867.n109 a_n2702_5867.n80 1.5
R17670 a_n2702_5867.n28 a_n2702_5867.n27 1.129
R17671 a_n2702_5867.n26 a_n2702_5867.n25 1.129
R17672 a_n2702_5867.n142 a_n2702_5867.n138 1.129
R17673 a_n2702_5867.n140 a_n2702_5867.n139 1.129
R17674 a_n2702_5867.n98 a_n2702_5867.n96 1.022
R17675 a_n2702_5867.n102 a_n2702_5867.n101 0.853
R17676 a_n2702_5867.n150 a_n2702_5867.n149 0.752
R17677 a_n2702_5867.n46 a_n2702_5867.n45 0.752
R17678 a_n2702_5867.n49 a_n2702_5867.n48 0.752
R17679 a_n2702_5867.n124 a_n2702_5867.n123 0.752
R17680 a_n2702_5867.n116 a_n2702_5867.n115 0.752
R17681 a_n2702_5867.n118 a_n2702_5867.n117 0.752
R17682 a_n2702_5867.n114 a_n2702_5867.n113 0.752
R17683 a_n2702_5867.n89 a_n2702_5867.n88 0.716
R17684 a_n2702_5867.n131 a_n2702_5867.n130 0.536
R17685 a_n2702_5867.n44 a_n2702_5867.n43 0.536
R17686 a_n2702_5867.n127 a_n2702_5867.n126 0.476
R17687 a_n2702_5867.n39 a_n2702_5867.n38 0.475
R17688 a_n2702_5867.n111 a_n2702_5867.n110 0.382
R17689 a_n2702_5867.n147 a_n2702_5867.n146 0.382
R17690 a_n2702_5867.n146 a_n2702_5867.n145 0.376
R17691 a_n2702_5867.n144 a_n2702_5867.n143 0.376
R17692 a_n2702_5867.n34 a_n2702_5867.n31 0.376
R17693 a_n2702_5867.n38 a_n2702_5867.n37 0.376
R17694 a_n2702_5867.n36 a_n2702_5867.n35 0.376
R17695 a_n2702_5867.n136 a_n2702_5867.n133 0.376
R17696 a_n2702_5867.n135 a_n2702_5867.n134 0.376
R17697 a_n2702_5867.n42 a_n2702_5867.n41 0.376
R17698 a_n2702_5867.n129 a_n2702_5867.n128 0.376
R17699 a_n2702_5867.n119 a_n2702_5867.n118 0.35
R17700 a_n2702_5867.n29 a_n2702_5867.n28 0.349
R17701 a_n2702_5867.n96 a_n2702_5867.n95 0.316
R17702 a_n2702_5867.n2 a_n2702_5867.n0 0.066
R17703 a_n2702_5867.n87 a_n2702_5867.n86 0.047
R17704 a_n2702_5867.n72 a_n2702_5867.n71 0.043
R17705 a_n2702_5867.n68 a_n2702_5867.n67 0.043
R17706 a_n2702_5867.n64 a_n2702_5867.n63 0.041
R17707 a_n2702_5867.n79 a_n2702_5867.n78 0.035
R17708 a_n2702_5867.n108 a_n2702_5867.n107 0.035
R17709 a_n2702_5867.n19 a_n2702_5867.n18 0.034
R17710 a_n2702_5867.n23 a_n2702_5867.n22 0.034
R17711 a_n2702_5867.n8 a_n2702_5867.n7 0.034
R17712 a_n2702_5867.n77 a_n2702_5867.n76 0.034
R17713 a_n2702_5867.n106 a_n2702_5867.n105 0.034
R17714 a_n2702_5867.n12 a_n2702_5867.n6 0.032
R17715 a_n2702_5867.n109 a_n2702_5867.n70 0.032
R17716 a_n2702_5867.n100 a_n2702_5867.n99 0.031
R17717 a_n2702_5867.n9 a_n2702_5867.n8 0.03
R17718 a_n2702_5867.n75 a_n2702_5867.n74 0.03
R17719 a_n2702_5867.n102 a_n2702_5867.n94 0.03
R17720 a_n2702_5867.n81 a_n2702_5867.n87 0.03
R17721 a_n2702_5867.n11 a_n2702_5867.n10 0.028
R17722 a_n2702_5867.n60 a_n2702_5867.n58 0.028
R17723 a_n2702_5867.n73 a_n2702_5867.n72 0.028
R17724 a_n2702_5867.n91 a_n2702_5867.n90 0.028
R17725 a_n2702_5867.n13 a_n2702_5867.n12 0.028
R17726 a_n2702_5867.n57 a_n2702_5867.n56 0.028
R17727 a_n2702_5867.n69 a_n2702_5867.n68 0.028
R17728 a_n2702_5867.n104 a_n2702_5867.n82 0.028
R17729 a_n2702_5867.n85 a_n2702_5867.n83 0.028
R17730 a_n2702_5867.n17 a_n2702_5867.n15 0.026
R17731 a_n2702_5867.n66 a_n2702_5867.n65 0.026
R17732 a_n2702_5867.n93 a_n2702_5867.n92 0.026
R17733 a_n2702_5867.n4 a_n2702_5867.n3 0.026
R17734 a_n2702_5867.n90 a_n2702_5867.n89 0.024
R17735 a_n2702_5867.n18 a_n2702_5867.n17 0.024
R17736 a_n2702_5867.n6 a_n2702_5867.n5 0.024
R17737 a_n2702_5867.n15 a_n2702_5867.n16 0.022
R17738 a_n2702_5867.n5 a_n2702_5867.n4 0.022
R17739 a_n2702_5867.n3 a_n2702_5867.n2 0.022
R17740 a_n2702_5867.n20 a_n2702_5867.n19 0.02
R17741 a_n2702_5867.n10 a_n2702_5867.n9 0.02
R17742 a_n2702_5867.n94 a_n2702_5867.n93 0.02
R17743 a_n2702_5867.n14 a_n2702_5867.n13 0.02
R17744 a_n2702_5867.n101 a_n2702_5867.n100 0.019
R17745 a_n2702_5867.n82 a_n2702_5867.n81 0.018
R17746 a_n2702_5867.n103 a_n2702_5867.n102 0.018
R17747 a_n2702_5867.n70 a_n2702_5867.n69 0.018
R17748 a_n2702_5867.n24 a_n2702_5867.n23 0.017
R17749 a_n2702_5867.n74 a_n2702_5867.n73 0.017
R17750 a_n2702_5867.n58 a_n2702_5867.n59 0.015
R17751 a_n2702_5867.n61 a_n2702_5867.n60 0.015
R17752 a_n2702_5867.n56 a_n2702_5867.n0 0.015
R17753 a_n2702_5867.n63 a_n2702_5867.n57 0.015
R17754 a_n2702_5867.n80 a_n2702_5867.n79 0.013
R17755 a_n2702_5867.n78 a_n2702_5867.n77 0.013
R17756 a_n2702_5867.n109 a_n2702_5867.n108 0.013
R17757 a_n2702_5867.n107 a_n2702_5867.n106 0.013
R17758 a_n2702_5867.n92 a_n2702_5867.n91 0.007
R17759 a_n2702_5867.n86 a_n2702_5867.n85 0.007
R17760 a_n2702_5867.n21 a_n2702_5867.n20 1.424
R17761 a_n2702_5867.n67 a_n2702_5867.n64 0.005
R17762 a_n2702_5867.n80 a_n2702_5867.n75 0.003
R17763 a_n2702_5867.n105 a_n2702_5867.n104 0.003
R17764 a_n2702_5867.n83 a_n2702_5867.n84 0.003
R17765 a_n2702_5867.n14 a_n2702_5867.n21 0.47
R17766 modi3.n5 modi3.t2 1037.94
R17767 modi3.n43 modi3.t3 1037.29
R17768 modi3.n43 modi3.t4 799.181
R17769 modi3.n5 modi3.t5 796.922
R17770 modi3.n151 modi3.n48 585
R17771 modi3.n127 modi3.n48 585
R17772 modi3.n69 modi3.n48 585
R17773 modi3.n61 modi3.n48 585
R17774 modi3.n250 modi3.n248 185
R17775 modi3.n232 modi3.n219 185
R17776 modi3.n231 modi3.n230 185
R17777 modi3.n270 modi3.n269 185
R17778 modi3.n231 modi3.n221 118.319
R17779 modi3.n271 modi3.n270 118.319
R17780 modi3.n292 modi3.n291 109.655
R17781 modi3.n281 modi3.n280 109.655
R17782 modi3.n291 modi3.n290 92.5
R17783 modi3.n282 modi3.n281 92.5
R17784 modi3.n291 modi3.t1 70.344
R17785 modi3.n281 modi3.t1 70.344
R17786 modi3.n292 modi3.n232 31.034
R17787 modi3.n280 modi3.n248 31.034
R17788 modi3.n120 modi3.n119 19.744
R17789 modi3.n182 modi3.n181 19.744
R17790 modi3.n195 modi3.n194 19.727
R17791 modi3.n110 modi3.n109 19.727
R17792 modi3.n97 modi3.n96 19.708
R17793 modi3.n206 modi3.n205 19.708
R17794 modi3.n149 modi3.n69 15.811
R17795 modi3.n152 modi3.n151 15.435
R17796 modi3.n136 modi3.n127 13.552
R17797 modi3.n164 modi3.n61 13.552
R17798 modi3.n269 modi3.n268 10.164
R17799 modi3.n230 modi3.n229 9.788
R17800 modi3.n227 modi3.n222 9.3
R17801 modi3.n229 modi3.n228 9.3
R17802 modi3.n240 modi3.n239 9.3
R17803 modi3.n294 modi3.n293 9.3
R17804 modi3.n293 modi3.n292 9.3
R17805 modi3.n238 modi3.n237 9.3
R17806 modi3.n279 modi3.n278 9.3
R17807 modi3.n280 modi3.n279 9.3
R17808 modi3.n256 modi3.n255 9.3
R17809 modi3.n258 modi3.n257 9.3
R17810 modi3.n223 modi3.n221 9.3
R17811 modi3.n272 modi3.n271 9.3
R17812 modi3.n266 modi3.n264 9.3
R17813 modi3.n268 modi3.n267 9.3
R17814 modi3.n126 modi3.n75 9.3
R17815 modi3.n132 modi3.n131 9.3
R17816 modi3.n161 modi3.n160 9.3
R17817 modi3.n172 modi3.n171 9.3
R17818 modi3.n164 modi3.n62 9.3
R17819 modi3.n99 modi3.n98 9.3
R17820 modi3.n108 modi3.n107 9.3
R17821 modi3.n111 modi3.n110 9.3
R17822 modi3.n118 modi3.n117 9.3
R17823 modi3.n121 modi3.n120 9.3
R17824 modi3.n124 modi3.n123 9.3
R17825 modi3.n137 modi3.n136 9.3
R17826 modi3.n134 modi3.n133 9.3
R17827 modi3.n96 modi3.n95 9.3
R17828 modi3.n174 modi3.n59 9.3
R17829 modi3.n182 modi3.n60 9.3
R17830 modi3.n180 modi3.n179 9.3
R17831 modi3.n194 modi3.n193 9.3
R17832 modi3.n197 modi3.n196 9.3
R17833 modi3.n205 modi3.n204 9.3
R17834 modi3.n208 modi3.n207 9.3
R17835 modi3.n163 modi3.n64 9.3
R17836 modi3.n150 modi3.n48 9.154
R17837 modi3.n162 modi3.n48 9.143
R17838 modi3.n128 modi3.n48 9.143
R17839 modi3.n125 modi3.n48 9.132
R17840 modi3.n173 modi3.n48 9.132
R17841 modi3.n181 modi3.n48 8.886
R17842 modi3.n119 modi3.n48 8.886
R17843 modi3.n109 modi3.n48 8.875
R17844 modi3.n195 modi3.n48 8.875
R17845 modi3.n97 modi3.n48 8.864
R17846 modi3.n206 modi3.n48 8.864
R17847 modi3.n290 modi3.n289 8.658
R17848 modi3.n282 modi3.n247 8.658
R17849 modi3.n290 modi3.n233 8.282
R17850 modi3.n283 modi3.n282 8.282
R17851 modi3.n48 modi3.t0 7.141
R17852 modi3.n207 modi3.n45 7.033
R17853 modi3.n98 modi3.n90 7.033
R17854 modi3.n301 modi3.n300 6.416
R17855 modi3.n302 modi3.n42 5.734
R17856 modi3.n293 modi3.n219 5.647
R17857 modi3.n279 modi3.n250 5.647
R17858 modi3.n236 modi3.n234 4.65
R17859 modi3.n150 modi3.n68 4.65
R17860 modi3.n283 modi3.n234 4.517
R17861 modi3.n152 modi3.n150 4.517
R17862 modi3.n273 modi3.n265 4.5
R17863 modi3.n296 modi3.n295 4.5
R17864 modi3.n244 modi3.n235 4.5
R17865 modi3.n246 modi3.n245 4.5
R17866 modi3.n251 modi3.n249 4.5
R17867 modi3.n259 modi3.n247 4.5
R17868 modi3.n254 modi3.n253 4.5
R17869 modi3.n243 modi3.n242 4.5
R17870 modi3.n218 modi3.n217 4.5
R17871 modi3.n220 modi3.n215 4.5
R17872 modi3.n241 modi3.n233 4.5
R17873 modi3.n289 modi3.n288 4.5
R17874 modi3.n284 modi3.n283 4.5
R17875 modi3.n275 modi3.n252 4.5
R17876 modi3.n277 modi3.n276 4.5
R17877 modi3.n226 modi3.n225 4.5
R17878 modi3.n94 modi3.n93 4.5
R17879 modi3.n106 modi3.n105 4.5
R17880 modi3.n86 modi3.n85 4.5
R17881 modi3.n116 modi3.n115 4.5
R17882 modi3.n84 modi3.n82 4.5
R17883 modi3.n140 modi3.n139 4.5
R17884 modi3.n145 modi3.n70 4.5
R17885 modi3.n158 modi3.n157 4.5
R17886 modi3.n170 modi3.n57 4.5
R17887 modi3.n177 modi3.n176 4.5
R17888 modi3.n178 modi3.n55 4.5
R17889 modi3.n52 modi3.n51 4.5
R17890 modi3.n199 modi3.n198 4.5
R17891 modi3.n203 modi3.n202 4.5
R17892 modi3.n47 modi3.n46 4.5
R17893 modi3.n192 modi3.n191 4.5
R17894 modi3.n169 modi3.n168 4.5
R17895 modi3.n113 modi3.n112 4.5
R17896 modi3.n83 modi3.n79 4.5
R17897 modi3.n138 modi3.n74 4.5
R17898 modi3.n81 modi3.n80 4.5
R17899 modi3.n122 modi3.n78 4.5
R17900 modi3.n135 modi3.n77 4.5
R17901 modi3.n130 modi3.n129 4.5
R17902 modi3.n153 modi3.n152 4.5
R17903 modi3.n149 modi3.n148 4.5
R17904 modi3.n147 modi3.n146 4.5
R17905 modi3.n88 modi3.n87 4.5
R17906 modi3.n184 modi3.n183 4.5
R17907 modi3.n54 modi3.n53 4.5
R17908 modi3.n50 modi3.n49 4.5
R17909 modi3.n166 modi3.n165 4.5
R17910 modi3.n159 modi3.n65 4.5
R17911 modi3.n155 modi3.n66 4.5
R17912 modi3.n175 modi3.n58 4.5
R17913 modi3.n210 modi3.n209 4.5
R17914 modi3.n92 modi3.n91 4.5
R17915 modi3.n101 modi3.n100 4.5
R17916 modi3.n289 modi3.n234 4.141
R17917 modi3.n110 modi3.n80 4.141
R17918 modi3.n150 modi3.n149 4.141
R17919 modi3.n194 modi3.n53 4.141
R17920 modi3.n232 modi3.n231 4.137
R17921 modi3.n270 modi3.n248 4.137
R17922 modi3.n225 modi3.n221 3.764
R17923 modi3.n229 modi3.n222 3.764
R17924 modi3.n256 modi3.n249 3.764
R17925 modi3.n120 modi3.n78 3.764
R17926 modi3.n165 modi3.n163 3.764
R17927 modi3.n126 modi3.n125 3.736
R17928 modi3.n6 modi3.n5 3.463
R17929 modi3.n238 modi3.n220 3.388
R17930 modi3.n268 modi3.n266 3.388
R17931 modi3.n271 modi3.n265 3.388
R17932 modi3.n96 modi3.n87 3.388
R17933 modi3.n135 modi3.n134 3.388
R17934 modi3.n183 modi3.n182 3.388
R17935 modi3.n205 modi3.n49 3.388
R17936 modi3.n173 modi3.n172 3.36
R17937 modi3.n293 modi3.n220 3.011
R17938 modi3.n239 modi3.n233 3.011
R17939 modi3.n266 modi3.n265 3.011
R17940 modi3.n108 modi3.n87 3.011
R17941 modi3.n136 modi3.n135 3.011
R17942 modi3.n131 modi3.n130 3.011
R17943 modi3.n172 modi3.n61 3.011
R17944 modi3.n183 modi3.n174 3.011
R17945 modi3.n196 modi3.n49 3.011
R17946 modi3.n225 modi3.n222 2.635
R17947 modi3.n257 modi3.n247 2.635
R17948 modi3.n279 modi3.n249 2.635
R17949 modi3.n124 modi3.n78 2.635
R17950 modi3.n127 modi3.n126 2.635
R17951 modi3.n161 modi3.n65 2.635
R17952 modi3.n165 modi3.n164 2.635
R17953 modi3.n272 modi3.n263 2.266
R17954 modi3.n223 modi3.n213 2.265
R17955 modi3.n239 modi3.n238 2.258
R17956 modi3.n257 modi3.n256 2.258
R17957 modi3.n118 modi3.n80 2.258
R17958 modi3.n180 modi3.n53 2.258
R17959 modi3.n301 modi3.n43 2.25
R17960 modi3.n131 modi3.n128 2.245
R17961 modi3.n162 modi3.n161 2.245
R17962 modi3 modi3.n301 2.02
R17963 modi3.n103 modi3.n102 1.755
R17964 modi3.n263 modi3.n262 1.755
R17965 modi3.n212 modi3.n211 1.705
R17966 modi3.n200 modi3.n44 1.705
R17967 modi3.n189 modi3.n188 1.705
R17968 modi3.n187 modi3.n186 1.705
R17969 modi3.n156 modi3.n56 1.705
R17970 modi3.n104 modi3.n103 1.705
R17971 modi3.n115 modi3.n72 1.705
R17972 modi3.n142 modi3.n141 1.705
R17973 modi3.n144 modi3.n143 1.705
R17974 modi3.n299 modi3.n213 1.705
R17975 modi3.n298 modi3.n297 1.705
R17976 modi3.n286 modi3.n214 1.705
R17977 modi3.n262 modi3.n261 1.705
R17978 modi3.n151 modi3.n65 1.505
R17979 modi3.n274 modi3.n273 1.5
R17980 modi3.n261 modi3.n251 1.5
R17981 modi3.n297 modi3.n215 1.5
R17982 modi3.n241 modi3.n216 1.5
R17983 modi3.n260 modi3.n259 1.5
R17984 modi3.n288 modi3.n287 1.5
R17985 modi3.n285 modi3.n284 1.5
R17986 modi3.n226 modi3.n224 1.5
R17987 modi3.n114 modi3.n81 1.5
R17988 modi3.n122 modi3.n73 1.5
R17989 modi3.n77 modi3.n76 1.5
R17990 modi3.n129 modi3.n71 1.5
R17991 modi3.n154 modi3.n153 1.5
R17992 modi3.n148 modi3.n67 1.5
R17993 modi3.n185 modi3.n184 1.5
R17994 modi3.n190 modi3.n54 1.5
R17995 modi3.n167 modi3.n166 1.5
R17996 modi3.n159 modi3.n63 1.5
R17997 modi3.n38 modi3.n36 1.402
R17998 modi3.n7 modi3.n6 1.355
R17999 modi3.n300 modi3.n212 1.284
R18000 modi3.n39 modi3.n38 1.141
R18001 modi3.n40 modi3.n39 1.137
R18002 modi3.n8 modi3.n7 1.137
R18003 modi3.n13 modi3.n12 1.137
R18004 modi3.n28 modi3.n27 1.137
R18005 modi3.n22 modi3.n21 1.137
R18006 modi3.n18 modi3.n17 1.137
R18007 modi3.n130 modi3.n69 1.129
R18008 modi3.n211 modi3.n45 1.127
R18009 modi3.n102 modi3.n90 1.127
R18010 modi3.n89 modi3.n88 1.125
R18011 modi3.n201 modi3.n50 1.125
R18012 modi3.n230 modi3.n219 0.752
R18013 modi3.n269 modi3.n250 0.752
R18014 modi3.n300 modi3.n299 0.719
R18015 modi3 modi3.n302 0.16
R18016 modi3.n98 modi3.n97 0.155
R18017 modi3.n207 modi3.n206 0.155
R18018 modi3.n302 modi3 0.155
R18019 modi3.n109 modi3.n108 0.144
R18020 modi3.n196 modi3.n195 0.144
R18021 modi3.n119 modi3.n118 0.133
R18022 modi3.n181 modi3.n180 0.133
R18023 modi3.n228 modi3.n218 0.053
R18024 modi3.n267 modi3.n252 0.053
R18025 modi3.n94 modi3.n92 0.053
R18026 modi3.n106 modi3.n86 0.053
R18027 modi3.n116 modi3.n82 0.053
R18028 modi3.n139 modi3.n75 0.053
R18029 modi3.n171 modi3.n170 0.053
R18030 modi3.n178 modi3.n177 0.053
R18031 modi3.n198 modi3.n52 0.053
R18032 modi3.n203 modi3.n47 0.053
R18033 modi3.n103 modi3.n72 0.05
R18034 modi3.n142 modi3.n72 0.05
R18035 modi3.n143 modi3.n142 0.05
R18036 modi3.n143 modi3.n56 0.05
R18037 modi3.n187 modi3.n56 0.05
R18038 modi3.n188 modi3.n187 0.05
R18039 modi3.n188 modi3.n44 0.05
R18040 modi3.n212 modi3.n44 0.05
R18041 modi3.n299 modi3.n298 0.05
R18042 modi3.n298 modi3.n214 0.05
R18043 modi3.n262 modi3.n214 0.05
R18044 modi3.n6 modi3.n4 0.048
R18045 modi3.n288 modi3.n235 0.045
R18046 modi3.n259 modi3.n254 0.045
R18047 modi3.n148 modi3.n147 0.045
R18048 modi3.n159 modi3.n158 0.045
R18049 modi3.n242 modi3.n241 0.043
R18050 modi3.n284 modi3.n246 0.043
R18051 modi3.n129 modi3.n70 0.043
R18052 modi3.n153 modi3.n66 0.043
R18053 modi3.n33 modi3.n32 0.037
R18054 modi3.n99 modi3.n92 0.034
R18055 modi3.n193 modi3.n52 0.032
R18056 modi3.n208 modi3.n47 0.032
R18057 modi3.n224 modi3.n217 0.03
R18058 modi3.n275 modi3.n274 0.03
R18059 modi3.n107 modi3.n106 0.03
R18060 modi3.n111 modi3.n86 0.03
R18061 modi3.n177 modi3.n175 0.03
R18062 modi3.n82 modi3.n79 0.028
R18063 modi3.n198 modi3.n197 0.028
R18064 modi3.n204 modi3.n203 0.028
R18065 modi3.n284 modi3.n236 0.025
R18066 modi3.n95 modi3.n94 0.025
R18067 modi3.n117 modi3.n116 0.025
R18068 modi3.n153 modi3.n68 0.025
R18069 modi3.n125 modi3.n124 0.024
R18070 modi3.n174 modi3.n173 0.024
R18071 modi3.n288 modi3.n236 0.023
R18072 modi3.n148 modi3.n68 0.023
R18073 modi3.n179 modi3.n178 0.023
R18074 modi3.n226 modi3.n223 0.021
R18075 modi3.n228 modi3.n227 0.021
R18076 modi3.n255 modi3.n251 0.021
R18077 modi3.n277 modi3.n252 0.021
R18078 modi3.n122 modi3.n121 0.021
R18079 modi3.n123 modi3.n75 0.021
R18080 modi3.n166 modi3.n64 0.021
R18081 modi3.n170 modi3.n169 0.021
R18082 modi3.n21 modi3.n20 0.021
R18083 modi3.n295 modi3.n218 0.019
R18084 modi3.n295 modi3.n294 0.019
R18085 modi3.n237 modi3.n215 0.019
R18086 modi3.n278 modi3.n277 0.019
R18087 modi3.n267 modi3.n264 0.019
R18088 modi3.n273 modi3.n272 0.019
R18089 modi3.n95 modi3.n88 0.019
R18090 modi3.n139 modi3.n138 0.019
R18091 modi3.n138 modi3.n137 0.019
R18092 modi3.n133 modi3.n77 0.019
R18093 modi3.n169 modi3.n62 0.019
R18094 modi3.n171 modi3.n59 0.019
R18095 modi3.n184 modi3.n60 0.019
R18096 modi3.n204 modi3.n50 0.019
R18097 modi3.n100 modi3.n90 0.019
R18098 modi3.n209 modi3.n45 0.019
R18099 modi3.n141 modi3.n73 0.018
R18100 modi3.n27 modi3.n26 0.018
R18101 modi3.n17 modi3.n16 0.018
R18102 modi3.n294 modi3.n215 0.017
R18103 modi3.n241 modi3.n240 0.017
R18104 modi3.n273 modi3.n264 0.017
R18105 modi3.n107 modi3.n88 0.017
R18106 modi3.n112 modi3.n81 0.017
R18107 modi3.n137 modi3.n77 0.017
R18108 modi3.n132 modi3.n129 0.017
R18109 modi3.n184 modi3.n59 0.017
R18110 modi3.n192 modi3.n54 0.017
R18111 modi3.n197 modi3.n50 0.017
R18112 modi3.n186 modi3.n185 0.017
R18113 modi3.n297 modi3.n216 0.016
R18114 modi3.n261 modi3.n260 0.016
R18115 modi3.n93 modi3.n91 0.016
R18116 modi3.n105 modi3.n85 0.016
R18117 modi3.n115 modi3.n84 0.016
R18118 modi3.n176 modi3.n55 0.016
R18119 modi3.n199 modi3.n51 0.016
R18120 modi3.n202 modi3.n46 0.016
R18121 modi3.n36 modi3.n35 0.016
R18122 modi3.n34 modi3.n33 0.016
R18123 modi3.n32 modi3.n31 0.016
R18124 modi3.n4 modi3.n3 0.016
R18125 modi3.n227 modi3.n226 0.015
R18126 modi3.n259 modi3.n258 0.015
R18127 modi3.n278 modi3.n251 0.015
R18128 modi3.n287 modi3.n244 0.015
R18129 modi3.n260 modi3.n253 0.015
R18130 modi3.n123 modi3.n122 0.015
R18131 modi3.n160 modi3.n159 0.015
R18132 modi3.n166 modi3.n62 0.015
R18133 modi3.n76 modi3.n71 0.015
R18134 modi3.n154 modi3.n67 0.015
R18135 modi3.n167 modi3.n63 0.015
R18136 modi3.n243 modi3.n216 0.014
R18137 modi3.n285 modi3.n245 0.014
R18138 modi3.n202 modi3.n201 0.014
R18139 modi3.n93 modi3.n89 0.013
R18140 modi3.n146 modi3.n67 0.013
R18141 modi3.n155 modi3.n154 0.013
R18142 modi3.n134 modi3.n128 0.012
R18143 modi3.n163 modi3.n162 0.012
R18144 modi3.n240 modi3.n237 0.012
R18145 modi3.n258 modi3.n255 0.012
R18146 modi3.n117 modi3.n81 0.012
R18147 modi3.n133 modi3.n132 0.012
R18148 modi3.n160 modi3.n64 0.012
R18149 modi3.n179 modi3.n54 0.012
R18150 modi3.n297 modi3.n296 0.011
R18151 modi3.n276 modi3.n261 0.011
R18152 modi3.n101 modi3.n91 0.011
R18153 modi3.n113 modi3.n85 0.011
R18154 modi3.n115 modi3.n114 0.011
R18155 modi3.n76 modi3.n74 0.011
R18156 modi3.n144 modi3.n71 0.011
R18157 modi3.n191 modi3.n51 0.011
R18158 modi3.n210 modi3.n46 0.011
R18159 modi3.n38 modi3.n37 0.011
R18160 modi3.n27 modi3.n24 0.011
R18161 modi3.n12 modi3.n11 0.011
R18162 modi3.n7 modi3.n2 0.011
R18163 modi3.n23 modi3.n22 0.011
R18164 modi3.n18 modi3.n14 0.011
R18165 modi3.n156 modi3.n63 0.01
R18166 modi3.n168 modi3.n167 0.01
R18167 modi3.n26 modi3.n25 0.01
R18168 modi3.n16 modi3.n15 0.01
R18169 modi3.n224 modi3.n213 0.009
R18170 modi3.n141 modi3.n140 0.009
R18171 modi3.n186 modi3.n57 0.009
R18172 modi3.n176 modi3.n58 0.009
R18173 modi3.n190 modi3.n189 0.009
R18174 modi3.n200 modi3.n199 0.009
R18175 modi3.n242 modi3.n235 0.008
R18176 modi3.n254 modi3.n246 0.008
R18177 modi3.n286 modi3.n285 0.008
R18178 modi3.n274 modi3.n263 0.008
R18179 modi3.n147 modi3.n70 0.008
R18180 modi3.n158 modi3.n66 0.008
R18181 modi3.n105 modi3.n104 0.008
R18182 modi3.n84 modi3.n83 0.008
R18183 modi3.n83 modi3.n73 0.008
R18184 modi3.n35 modi3.n34 0.008
R18185 modi3.n287 modi3.n286 0.007
R18186 modi3.n276 modi3.n275 0.007
R18187 modi3.n185 modi3.n58 0.007
R18188 modi3.n30 modi3.n29 0.007
R18189 modi3.n22 modi3.n19 0.007
R18190 modi3.n19 modi3.n18 0.007
R18191 modi3.n10 modi3.n9 0.007
R18192 modi3.n28 modi3.n23 0.007
R18193 modi3.n14 modi3.n13 0.007
R18194 modi3.n296 modi3.n217 0.006
R18195 modi3.n112 modi3.n111 0.006
R18196 modi3.n121 modi3.n79 0.006
R18197 modi3.n175 modi3.n60 0.006
R18198 modi3.n193 modi3.n192 0.006
R18199 modi3.n168 modi3.n57 0.006
R18200 modi3.n104 modi3.n89 0.005
R18201 modi3.n114 modi3.n113 0.005
R18202 modi3.n140 modi3.n74 0.005
R18203 modi3.n191 modi3.n190 0.005
R18204 modi3.n211 modi3.n210 0.005
R18205 modi3.n100 modi3.n99 0.004
R18206 modi3.n209 modi3.n208 0.004
R18207 modi3.n102 modi3.n101 0.004
R18208 modi3.n201 modi3.n200 0.004
R18209 modi3.n29 modi3.n28 0.004
R18210 modi3.n13 modi3.n10 0.004
R18211 modi3.n9 modi3.n8 0.004
R18212 modi3.n157 modi3.n156 0.003
R18213 modi3.n41 modi3.n40 0.002
R18214 modi3.n1 modi3.n0 0.002
R18215 modi3.n42 modi3.n41 0.002
R18216 modi3.n40 modi3.n1 0.002
R18217 modi3.n39 modi3.n30 0.002
R18218 modi3.n244 modi3.n243 0.002
R18219 modi3.n253 modi3.n245 0.002
R18220 modi3.n146 modi3.n145 0.002
R18221 modi3.n157 modi3.n155 0.002
R18222 modi3.n145 modi3.n144 0.001
R18223 modi3.n189 modi3.n55 0.001
R18224 modi.n2 modi.t1 1037.94
R18225 modi.n2 modi.t0 796.922
R18226 modi.n5 modi.n2 3.462
R18227 modi.n38 modi.n37 1.402
R18228 modi.n7 modi.n5 1.355
R18229 modi.n39 modi.n38 1.141
R18230 modi.n40 modi.n39 1.137
R18231 modi.n28 modi.n27 1.137
R18232 modi.n8 modi.n7 1.137
R18233 modi.n13 modi.n12 1.137
R18234 modi.n18 modi.n17 1.137
R18235 modi.n22 modi.n21 1.137
R18236 modi modi.n42 0.111
R18237 modi.n5 modi.n4 0.048
R18238 modi.n34 modi.n33 0.037
R18239 modi.n21 modi.n20 0.021
R18240 modi.n17 modi.n16 0.018
R18241 modi.n27 modi.n25 0.018
R18242 modi.n4 modi.n3 0.016
R18243 modi.n33 modi.n32 0.016
R18244 modi.n35 modi.n34 0.016
R18245 modi.n37 modi.n36 0.016
R18246 modi.n7 modi.n6 0.011
R18247 modi.n12 modi.n11 0.011
R18248 modi.n27 modi.n26 0.011
R18249 modi.n38 modi.n31 0.011
R18250 modi.n18 modi.n14 0.011
R18251 modi.n23 modi.n22 0.011
R18252 modi.n16 modi.n15 0.01
R18253 modi.n25 modi.n24 0.01
R18254 modi.n36 modi.n35 0.008
R18255 modi.n10 modi.n9 0.007
R18256 modi.n19 modi.n18 0.007
R18257 modi.n22 modi.n19 0.007
R18258 modi.n30 modi.n29 0.007
R18259 modi.n14 modi.n13 0.007
R18260 modi.n28 modi.n23 0.007
R18261 modi.n9 modi.n8 0.004
R18262 modi.n13 modi.n10 0.004
R18263 modi.n29 modi.n28 0.004
R18264 modi.n40 modi.n1 0.002
R18265 modi.n42 modi.n41 0.002
R18266 modi.n1 modi.n0 0.002
R18267 modi.n41 modi.n40 0.002
R18268 modi.n39 modi.n30 0.002
R18269 modo.n257 modo.t3 1037.29
R18270 modo modo.t2 796.136
R18271 modo.n30 modo.n29 92.5
R18272 modo.n46 modo.n45 92.5
R18273 modo.n45 modo.t1 70.344
R18274 modo.n8 modo.n7 31.034
R18275 modo.n65 modo.n64 31.034
R18276 modo.n113 modo.n112 9.3
R18277 modo.n190 modo.n189 9.3
R18278 modo.n15 modo.n14 9.3
R18279 modo.n66 modo.n65 9.3
R18280 modo.n9 modo.n8 9.3
R18281 modo.n77 modo.n76 9.3
R18282 modo.n229 modo.n228 9.154
R18283 modo.n257 modo.n256 8.715
R18284 modo.n31 modo.n30 8.282
R18285 modo.n47 modo.n46 8.282
R18286 modo.n228 modo.t0 7.141
R18287 modo.n149 modo.n148 7.033
R18288 modo.n92 modo.n91 7.033
R18289 modo.n9 modo.n5 5.647
R18290 modo.n66 modo.n62 5.647
R18291 modo.n230 modo.n229 4.65
R18292 modo.n44 modo.n43 4.65
R18293 modo.n176 modo.n175 4.5
R18294 modo.n196 modo.n195 4.5
R18295 modo.n209 modo.n208 4.5
R18296 modo.n216 modo.n213 4.5
R18297 modo.n225 modo.n224 4.5
R18298 modo.n231 modo.n227 4.5
R18299 modo.n100 modo.n97 4.5
R18300 modo.n107 modo.n106 4.5
R18301 modo.n119 modo.n118 4.5
R18302 modo.n129 modo.n128 4.5
R18303 modo.n139 modo.n138 4.5
R18304 modo.n163 modo.n162 4.5
R18305 modo.n83 modo.n81 4.5
R18306 modo.n70 modo.n67 4.5
R18307 modo.n57 modo.n55 4.5
R18308 modo.n32 modo.n31 4.5
R18309 modo.n39 modo.n38 4.5
R18310 modo.n48 modo.n47 4.5
R18311 modo.n12 modo.n11 4.5
R18312 modo.n20 modo.n19 4.5
R18313 modo.n128 modo.n125 4.141
R18314 modo.n162 modo.n161 4.141
R18315 modo.n7 modo.n6 4.137
R18316 modo.n64 modo.n63 4.137
R18317 modo.n118 modo.n115 3.764
R18318 modo.n208 modo.n206 3.764
R18319 modo.n19 modo.n17 3.764
R18320 modo.n67 modo.n60 3.764
R18321 modo.n138 modo.n135 3.388
R18322 modo.n106 modo.n105 3.388
R18323 modo.n195 modo.n194 3.388
R18324 modo.n175 modo.n174 3.388
R18325 modo.n11 modo.n10 3.388
R18326 modo.n81 modo.n80 3.388
R18327 modo.n138 modo.n137 3.011
R18328 modo.n106 modo.n103 3.011
R18329 modo.n97 modo.n95 3.011
R18330 modo.n189 modo.n188 3.011
R18331 modo.n195 modo.n193 3.011
R18332 modo.n175 modo.n173 3.011
R18333 modo.n11 modo.n9 3.011
R18334 modo.n31 modo.n28 3.011
R18335 modo.n81 modo.n79 3.011
R18336 modo.n118 modo.n117 2.635
R18337 modo.n112 modo.n111 2.635
R18338 modo.n213 modo.n212 2.635
R18339 modo.n208 modo.n207 2.635
R18340 modo.n19 modo.n18 2.635
R18341 modo.n55 modo.n54 2.635
R18342 modo.n67 modo.n66 2.635
R18343 modo.n128 modo.n127 2.258
R18344 modo.n162 modo.n160 2.258
R18345 modo.n25 modo.n0 1.754
R18346 modo.n179 modo.n150 1.754
R18347 modo.n25 modo.n24 1.705
R18348 modo.n42 modo.n41 1.705
R18349 modo.n72 modo.n71 1.705
R18350 modo.n86 modo.n85 1.705
R18351 modo.n255 modo.n144 1.705
R18352 modo.n199 modo.n198 1.705
R18353 modo.n219 modo.n218 1.705
R18354 modo.n248 modo.n247 1.705
R18355 modo.n254 modo.n253 1.705
R18356 modo.n242 modo.n241 1.705
R18357 modo.n236 modo.n235 1.705
R18358 modo.n185 modo.n184 1.705
R18359 modo.n179 modo.n178 1.705
R18360 modo.n213 modo.n211 1.505
R18361 modo.n197 modo.n196 1.5
R18362 modo.n210 modo.n209 1.5
R18363 modo.n217 modo.n216 1.5
R18364 modo.n226 modo.n225 1.5
R18365 modo.n232 modo.n231 1.5
R18366 modo.n84 modo.n83 1.5
R18367 modo.n71 modo.n70 1.5
R18368 modo.n33 modo.n32 1.5
R18369 modo.n58 modo.n57 1.5
R18370 modo.n40 modo.n39 1.5
R18371 modo.n49 modo.n48 1.5
R18372 modo.n24 modo.n12 1.5
R18373 modo.n21 modo.n20 1.5
R18374 modo modo.n257 1.439
R18375 modo.n256 modo.n255 1.268
R18376 modo.n97 modo.n96 1.129
R18377 modo.n150 modo.n149 1.127
R18378 modo.n144 modo.n92 1.127
R18379 modo.n140 modo.n139 1.125
R18380 modo.n177 modo.n176 1.125
R18381 modo.n5 modo.n4 0.752
R18382 modo.n62 modo.n61 0.752
R18383 modo.n256 modo.n86 0.709
R18384 modo.n91 modo.n90 0.155
R18385 modo.n148 modo.n147 0.155
R18386 modo.n137 modo.n136 0.144
R18387 modo.n173 modo.n172 0.144
R18388 modo.n127 modo.n126 0.133
R18389 modo.n160 modo.n159 0.132
R18390 modo.n133 modo.n132 0.053
R18391 modo.n123 modo.n122 0.053
R18392 modo.n113 modo.n110 0.053
R18393 modo.n157 modo.n156 0.053
R18394 modo.n167 modo.n166 0.053
R18395 modo.n170 modo.n169 0.053
R18396 modo.n77 modo.n75 0.053
R18397 modo.n42 modo.n25 0.049
R18398 modo.n72 modo.n42 0.049
R18399 modo.n86 modo.n72 0.049
R18400 modo.n255 modo.n254 0.049
R18401 modo.n254 modo.n248 0.049
R18402 modo.n248 modo.n242 0.049
R18403 modo.n242 modo.n236 0.049
R18404 modo.n236 modo.n219 0.049
R18405 modo.n219 modo.n199 0.049
R18406 modo.n199 modo.n185 0.049
R18407 modo.n185 modo.n179 0.049
R18408 modo.n39 modo.n37 0.045
R18409 modo.n57 modo.n53 0.045
R18410 modo.n100 modo.n99 0.043
R18411 modo.n225 modo.n223 0.043
R18412 modo.n88 modo.n87 0.034
R18413 modo.n166 modo.n165 0.032
R18414 modo.n134 modo.n133 0.03
R18415 modo.n132 modo.n131 0.03
R18416 modo.n156 modo.n155 0.03
R18417 modo.n22 modo.n21 0.03
R18418 modo.n84 modo.n74 0.03
R18419 modo.n122 modo.n121 0.028
R18420 modo.n168 modo.n167 0.028
R18421 modo.n171 modo.n170 0.028
R18422 modo.n94 modo.n93 0.025
R18423 modo.n124 modo.n123 0.025
R18424 modo.n48 modo.n44 0.025
R18425 modo.n117 modo.n116 0.024
R18426 modo.n193 modo.n192 0.024
R18427 modo.n231 modo.n230 0.023
R18428 modo.n158 modo.n157 0.023
R18429 modo.n120 modo.n119 0.021
R18430 modo.n114 modo.n113 0.021
R18431 modo.n203 modo.n202 0.021
R18432 modo.n20 modo.n13 0.021
R18433 modo.n16 modo.n15 0.021
R18434 modo.n70 modo.n59 0.021
R18435 modo.n139 modo.n94 0.019
R18436 modo.n110 modo.n109 0.019
R18437 modo.n109 modo.n108 0.019
R18438 modo.n107 modo.n102 0.019
R18439 modo.n204 modo.n203 0.019
R18440 modo.n191 modo.n190 0.019
R18441 modo.n176 modo.n171 0.019
R18442 modo.n2 modo.n1 0.019
R18443 modo.n3 modo.n2 0.019
R18444 modo.n69 modo.n68 0.019
R18445 modo.n78 modo.n77 0.019
R18446 modo.n83 modo.n82 0.019
R18447 modo.n92 modo.n89 0.019
R18448 modo.n149 modo.n146 0.019
R18449 modo.n198 modo.n197 0.018
R18450 modo.n139 modo.n134 0.017
R18451 modo.n130 modo.n129 0.017
R18452 modo.n108 modo.n107 0.017
R18453 modo.n101 modo.n100 0.017
R18454 modo.n196 modo.n191 0.017
R18455 modo.n164 modo.n163 0.017
R18456 modo.n176 modo.n168 0.017
R18457 modo.n12 modo.n3 0.017
R18458 modo.n32 modo.n27 0.017
R18459 modo.n83 modo.n78 0.017
R18460 modo.n142 modo.n141 0.016
R18461 modo.n252 modo.n251 0.016
R18462 modo.n246 modo.n245 0.016
R18463 modo.n181 modo.n180 0.016
R18464 modo.n153 modo.n152 0.016
R18465 modo.n71 modo.n58 0.016
R18466 modo.n119 modo.n114 0.015
R18467 modo.n216 modo.n215 0.015
R18468 modo.n209 modo.n204 0.015
R18469 modo.n238 modo.n237 0.015
R18470 modo.n232 modo.n226 0.015
R18471 modo.n217 modo.n210 0.015
R18472 modo.n20 modo.n16 0.015
R18473 modo.n57 modo.n56 0.015
R18474 modo.n70 modo.n69 0.015
R18475 modo.n40 modo.n35 0.015
R18476 modo.n58 modo.n51 0.015
R18477 modo.n177 modo.n153 0.014
R18478 modo.n34 modo.n33 0.014
R18479 modo.n50 modo.n49 0.014
R18480 modo.n141 modo.n140 0.013
R18481 modo.n233 modo.n232 0.013
R18482 modo.n226 modo.n221 0.013
R18483 modo.n105 modo.n104 0.012
R18484 modo.n206 modo.n205 0.012
R18485 modo.n129 modo.n124 0.012
R18486 modo.n102 modo.n101 0.012
R18487 modo.n215 modo.n214 0.012
R18488 modo.n163 modo.n158 0.012
R18489 modo.n27 modo.n26 0.012
R18490 modo.n143 modo.n142 0.011
R18491 modo.n251 modo.n250 0.011
R18492 modo.n239 modo.n238 0.011
R18493 modo.n218 modo.n217 0.011
R18494 modo.n182 modo.n181 0.011
R18495 modo.n152 modo.n151 0.011
R18496 modo.n24 modo.n23 0.011
R18497 modo.n210 modo.n201 0.01
R18498 modo.n184 modo.n183 0.01
R18499 modo.n253 modo.n252 0.009
R18500 modo.n241 modo.n240 0.009
R18501 modo.n187 modo.n186 0.009
R18502 modo.n99 modo.n98 0.008
R18503 modo.n223 modo.n222 0.008
R18504 modo.n245 modo.n244 0.008
R18505 modo.n244 modo.n243 0.008
R18506 modo.n37 modo.n36 0.008
R18507 modo.n53 modo.n52 0.008
R18508 modo.n85 modo.n84 0.008
R18509 modo.n197 modo.n187 0.007
R18510 modo.n41 modo.n40 0.007
R18511 modo.n74 modo.n73 0.007
R18512 modo.n131 modo.n130 0.006
R18513 modo.n121 modo.n120 0.006
R18514 modo.n155 modo.n154 0.006
R18515 modo.n165 modo.n164 0.006
R18516 modo.n201 modo.n200 0.006
R18517 modo.n23 modo.n22 0.006
R18518 modo.n144 modo.n143 0.005
R18519 modo.n250 modo.n249 0.005
R18520 modo.n240 modo.n239 0.005
R18521 modo.n183 modo.n182 0.005
R18522 modo.n178 modo.n177 0.005
R18523 modo.n89 modo.n88 0.004
R18524 modo.n146 modo.n145 0.004
R18525 modo.n235 modo.n234 0.002
R18526 modo.n234 modo.n233 0.002
R18527 modo.n221 modo.n220 0.002
R18528 modo.n35 modo.n34 0.002
R18529 modo.n51 modo.n50 0.002
R18530 modo.n247 modo.n246 0.001
R18531 P0 P0.t0 1038.51
R18532 P0 P0.t1 796.136
R18533 P6 P6.t0 1038.31
R18534 P6 P6.t1 796.506
R18535 P3 P3.t1 1038.7
R18536 P3 P3.t0 796.11
R18537 P2 P2.t0 1038.73
R18538 P2 P2.t1 796.136
R18539 P4 P4.t0 1038.31
R18540 P4 P4.t1 798.111
R18541 P5 P5.t1 1038.31
R18542 P5 P5.t0 796.506
C0 a_n10460_2476# a_n8769_2484# 0.03fF
C1 a_n15024_8436# fout0 0.03fF
C2 a_n5187_8439# VDD 1.44fF
C3 a_n11112_5995# fout4 0.04fF
C4 a_n10992_8440# a_n9840_8440# 0.06fF
C5 a_n11944_11462# a_n9159_8440# 0.06fF
C6 a_n5187_8439# a_n4036_12366# 0.03fF
C7 a_n6140_11462# a_n3749_8439# 0.43fF
C8 a_n16325_2475# modi5 0.27fF
C9 a_n17419_5897# a_n17674_2475# 0.08fF
C10 a_n5187_8439# modi2 0.10fF
C11 a_n12800_11551# fout1 0.03fF
C12 a_n18665_11548# a_n18465_11548# 0.97fF
C13 a_n17149_12355# modi0 0.02fF
C14 a_n16976_5994# VDD 1.02fF
C15 a_n4792_8439# a_n4035_8439# 0.02fF
C16 a_n4604_2477# a_n5954_2477# 0.03fF
C17 a_n4261_5899# a_n5273_2477# 0.03fF
C18 a_n16993_2475# a_n16237_2475# 0.01fF
C19 a_n16325_2475# a_n15538_5994# 0.11fF
C20 a_n3749_8439# modi3 0.05fF
C21 a_n17143_8436# VDD 0.94fF
C22 a_n3817_5996# fout4 0.03fF
C23 a_n14284_11547# modi1 0.07fF
C24 a_n21205_8431# fout0 0.15fF
C25 a_n21734_5903# fout 0.23fF
C26 a_n6652_2485# modi4 0.08fF
C27 a_n24251_11543# fin 0.04fF
C28 fout0 modi0 2.00fF
C29 VDD P2 0.32fF
C30 a_n4604_2477# a_n4498_5996# 0.73fF
C31 a_n13930_2482# P6 0.02fF
C32 a_n4261_5899# a_n3817_5996# 0.69fF
C33 a_n16468_12355# a_n15707_12363# 0.01fF
C34 a_n9674_5995# VDD 0.94fF
C35 VDD fout5 4.75fF
C36 a_n23172_5903# a_n21972_6000# 0.07fF
C37 a_n14130_2482# fout6 0.13fF
C38 a_n20386_2489# fout 1.05fF
C39 a_n4604_2477# fout3 1.64fF
C40 fout modi 0.72fF
C41 a_n15419_8436# a_n16462_8436# 0.07fF
C42 a_n22077_2481# a_n22746_2481# 0.06fF
C43 a_n21734_5903# a_n21989_2481# 0.08fF
C44 a_n11793_5995# a_n11112_5995# 0.02fF
C45 a_n11555_5898# a_n10460_2476# 0.49fF
C46 fout5 P6 0.56fF
C47 a_n17419_5897# modi6 0.05fF
C48 a_n17810_11459# fout1 0.43fF
C49 a_n8419_11550# modi1 0.04fF
C50 a_n15419_8436# fout0 0.79fF
C51 a_n8769_2484# fout5 1.05fF
C52 a_n23595_11454# a_n22928_8431# 0.09fF
C53 a_n12800_11551# a_n12600_11551# 0.97fF
C54 a_n5255_5996# modi3 0.06fF
C55 a_n22928_8431# fin 0.02fF
C56 a_n5954_2477# a_n5273_2477# 0.01fF
C57 a_n10460_2476# fout4 1.45fF
C58 a_n23172_5903# fout6 0.79fF
C59 a_n17419_5897# a_n16237_2475# 0.04fF
C60 a_n6353_11550# modi2 0.09fF
C61 a_n11944_11462# fout1 1.50fF
C62 a_n16325_2475# VDD 1.39fF
C63 a_n3835_2477# fout4 0.04fF
C64 a_n11277_8440# fout2 0.02fF
C65 a_n4035_8439# a_n3354_8439# 0.02fF
C66 a_n16237_2475# a_n15556_2475# 0.01fF
C67 a_n4604_2477# a_n4516_2477# 0.34fF
C68 a_n4261_5899# a_n3835_2477# 0.35fF
C69 a_n10602_12359# a_n9841_12367# 0.01fF
C70 a_n15024_8436# modi0 0.64fF
C71 a_n11112_5995# modi4 0.06fF
C72 a_n24451_11543# a_n23808_11542# 0.02fF
C73 a_n23595_11454# a_n22643_8431# 0.85fF
C74 a_n5273_2477# fout3 0.04fF
C75 a_n15705_8436# VDD 1.03fF
C76 a_n22928_8431# a_n22247_8431# 0.02fF
C77 a_n5187_8439# a_n5473_8439# 0.66fF
C78 a_n6140_11462# a_n4792_8439# 0.67fF
C79 a_n12800_11551# modi1 0.09fF
C80 a_n15981_5897# fout6 0.29fF
C81 a_n22643_8431# fin 0.87fF
C82 a_n4498_5996# a_n3817_5996# 0.02fF
C83 a_n22728_6000# a_n22077_2481# 0.12fF
C84 a_n19682_2488# fout 0.12fF
C85 a_n3817_5996# fout3 0.04fF
C86 a_n15419_8436# a_n15024_8436# 0.15fF
C87 a_n6995_11551# a_n6795_11551# 0.97fF
C88 a_n6652_2485# modi3 0.04fF
C89 a_n11793_5995# a_n10460_2476# 0.06fF
C90 a_n11112_5995# a_n10117_5898# 0.06fF
C91 a_n6795_11551# fout3 0.13fF
C92 a_n21734_5903# a_n20386_2489# 0.04fF
C93 a_n22077_2481# a_n21308_2481# 0.04fF
C94 a_n11555_5898# fout5 0.17fF
C95 a_n21492_12358# a_n20815_12350# 0.01fF
C96 a_n21205_8431# modi0 0.05fF
C97 a_n24251_11543# modo 0.09fF
C98 a_n22728_6000# VDD 1.03fF
C99 VDD fout2 4.38fF
C100 fout0 P1 0.68fF
C101 a_n4036_12366# fout2 0.04fF
C102 VDD modi5 1.37fF
C103 fout2 modi2 1.99fF
C104 a_n8066_2483# fout5 0.12fF
C105 a_n22643_8431# a_n22247_8431# 0.15fF
C106 a_n23595_11454# a_n21491_8431# 0.12fF
C107 a_n4604_2477# modi3 0.27fF
C108 fout fout6 2.92fF
C109 a_n5273_2477# a_n4516_2477# 0.01fF
C110 a_n21491_8431# fin 0.03fF
C111 a_n9674_5995# fout4 0.04fF
C112 a_n4797_12358# a_n4036_12366# 0.01fF
C113 fout5 fout4 3.03fF
C114 modi5 P6 0.13fF
C115 a_n23409_6000# fout6 0.02fF
C116 a_n4797_12358# modi2 0.02fF
C117 a_n17810_11459# a_n16857_8436# 0.85fF
C118 a_n18665_11548# a_n18023_11547# 0.02fF
C119 a_n15419_8436# modi0 0.80fF
C120 a_n2409_2484# fout4 0.13fF
C121 a_n15538_5994# VDD 0.94fF
C122 a_n4604_2477# a_n2913_2485# 0.03fF
C123 a_n10460_2476# modi4 0.27fF
C124 a_n23172_5903# modi6 0.82fF
C125 a_n23595_11454# a_n23808_11542# 0.03fF
C126 a_n3835_2477# fout3 0.03fF
C127 a_n11277_8440# VDD 0.91fF
C128 a_n22247_8431# a_n21491_8431# 0.02fF
C129 a_n5187_8439# a_n4035_8439# 0.06fF
C130 a_n6140_11462# a_n3354_8439# 0.06fF
C131 a_n11944_11462# modi1 0.25fF
C132 a_n23808_11542# fin 0.05fF
C133 a_n11555_5898# a_n11810_2476# 0.08fF
C134 a_n16993_2475# fout5 0.05fF
C135 a_n23427_2481# modi6 0.36fF
C136 a_n15707_12363# a_n15030_12355# 0.01fF
C137 a_n5699_5899# VDD 1.32fF
C138 a_n21734_5903# a_n21972_6000# 0.15fF
C139 a_n5273_2477# modi3 0.05fF
C140 a_n5187_8439# fout3 0.27fF
C141 a_n11112_5995# a_n10355_5995# 0.02fF
C142 a_n10117_5898# a_n10460_2476# 0.85fF
C143 a_n12800_11551# P2 0.02fF
C144 a_n17149_12355# fout1 0.04fF
C145 a_n22643_8431# modo 0.10fF
C146 a_n22077_2481# VDD 1.30fF
C147 a_n18372_2483# modi5 0.04fF
C148 a_n20386_2489# a_n19682_2488# 0.02fF
C149 a_n12800_11551# a_n12157_11550# 0.02fF
C150 a_n11944_11462# a_n10992_8440# 0.85fF
C151 a_n17419_5897# a_n16976_5994# 0.70fF
C152 a_n4516_2477# a_n3835_2477# 0.01fF
C153 a_n11555_5898# modi5 0.05fF
C154 a_n9554_8440# a_n10596_8440# 0.07fF
C155 a_n21734_5903# fout6 0.86fF
C156 modi0 P1 0.11fF
C157 fout0 fout1 2.91fF
C158 VDD modi2 1.30fF
C159 a_n24251_11543# fout0 0.13fF
C160 a_n16325_2475# a_n16993_2475# 0.06fF
C161 a_n15981_5897# a_n16237_2475# 0.08fF
C162 a_n4036_12366# modi2 0.05fF
C163 a_n5699_5899# a_n5936_5996# 0.15fF
C164 a_n11283_12359# fout1 0.06fF
C165 a_n17810_11459# a_n18023_11547# 0.03fF
C166 VDD P6 0.34fF
C167 fout2 P3 0.68fF
C168 a_n5473_8439# fout2 0.03fF
C169 a_n20386_2489# fout6 0.05fF
C170 a_n14633_2483# a_n14130_2482# 0.02fF
C171 modi fout6 0.13fF
C172 fout modi6 0.54fF
C173 a_n17810_11459# a_n17143_8436# 0.10fF
C174 a_n9841_12367# a_n9164_12359# 0.01fF
C175 a_n21491_8431# modo 0.06fF
C176 fout5 modi4 0.57fF
C177 modi5 fout4 0.13fF
C178 a_n17419_5897# fout5 0.79fF
C179 a_n22643_8431# a_n22934_12350# 0.35fF
C180 a_n23595_11454# a_n22253_12350# 0.34fF
C181 a_n23409_6000# modi6 0.68fF
C182 a_n2409_2484# fout3 0.04fF
C183 a_n9840_8440# VDD 1.02fF
C184 a_n21491_8431# a_n20810_8431# 0.02fF
C185 a_n8419_11550# fout2 0.05fF
C186 a_n18465_11548# fout0 0.04fF
C187 a_n11555_5898# a_n10372_2476# 0.04fF
C188 a_n15556_2475# fout5 0.06fF
C189 a_n21989_2481# modi6 0.02fF
C190 a_n5936_5996# VDD 1.10fF
C191 a_n22077_2481# a_n21291_6000# 0.10fF
C192 a_n22928_8431# fout0 0.03fF
C193 a_n6995_11551# a_n6353_11550# 0.02fF
C194 a_n6140_11462# a_n5187_8439# 0.85fF
C195 a_n3835_2477# modi3 0.02fF
C196 a_n10460_2476# a_n10355_5995# 0.73fF
C197 a_n10117_5898# a_n9674_5995# 0.69fF
C198 a_n6353_11550# fout3 1.08fF
C199 a_n10117_5898# fout5 0.27fF
C200 a_n21291_6000# VDD 0.94fF
C201 a_n23808_11542# modo 0.08fF
C202 a_n16993_2475# modi5 0.05fF
C203 a_n11944_11462# a_n12157_11550# 0.03fF
C204 a_n17419_5897# a_n16325_2475# 0.50fF
C205 a_n17657_5994# a_n16976_5994# 0.02fF
C206 a_n5699_5899# fout4 0.14fF
C207 a_n12800_11551# fout2 0.12fF
C208 a_n4036_12366# a_n3360_12358# 0.01fF
C209 a_n9554_8440# a_n9159_8440# 0.15fF
C210 a_n21972_6000# fout6 0.02fF
C211 a_n22643_8431# fout0 0.25fF
C212 a_n11810_2476# modi4 0.36fF
C213 a_n15981_5897# a_n14633_2483# 0.04fF
C214 a_n16325_2475# a_n15556_2475# 0.04fF
C215 a_n5699_5899# a_n4261_5899# 0.09fF
C216 a_n3360_12358# modi2 0.35fF
C217 a_n16857_8436# a_n17149_12355# 0.35fF
C218 a_n17810_11459# a_n16468_12355# 0.34fF
C219 a_n11555_5898# VDD 1.39fF
C220 a_n4035_8439# fout2 0.03fF
C221 a_n19682_2488# fout6 0.03fF
C222 a_n14130_2482# a_n13930_2482# 0.97fF
C223 a_n16857_8436# a_n16462_8436# 0.15fF
C224 a_n17810_11459# a_n15705_8436# 0.12fF
C225 VDD P0 0.25fF
C226 a_n23172_5903# a_n24125_2489# 0.06fF
C227 a_n17657_5994# fout5 0.02fF
C228 a_n21734_5903# modi6 0.11fF
C229 a_n23595_11454# a_n21492_12358# 0.06fF
C230 modi0 fout1 0.56fF
C231 VDD P3 0.32fF
C232 fout0 modi1 0.12fF
C233 a_n5473_8439# VDD 0.94fF
C234 a_n6995_11551# fout2 0.03fF
C235 a_n11283_12359# modi1 0.02fF
C236 a_n16857_8436# fout0 0.81fF
C237 modi2 P3 0.11fF
C238 a_n21492_12358# fin 0.05fF
C239 fout2 fout3 2.94fF
C240 VDD fout4 4.84fF
C241 a_n14130_2482# fout5 0.04fF
C242 a_n20386_2489# modi6 0.10fF
C243 a_n4261_5899# VDD 1.43fF
C244 modi modi6 0.07fF
C245 fout P7 0.04fF
C246 a_n8769_2484# a_n8066_2483# 0.02fF
C247 modi5 modi4 0.07fF
C248 fout5 P5 0.04fF
C249 a_n6140_11462# a_n6353_11550# 0.03fF
C250 a_n17419_5897# modi5 0.82fF
C251 a_n2409_2484# modi3 0.09fF
C252 a_n10355_5995# a_n9674_5995# 0.02fF
C253 a_n8419_11550# modi2 0.07fF
C254 a_n15419_8436# fout1 0.17fF
C255 a_n18465_11548# modi0 0.11fF
C256 a_n8769_2484# fout4 0.04fF
C257 a_n22253_12350# modo 0.02fF
C258 a_n15556_2475# modi5 0.02fF
C259 a_n5699_5899# a_n5954_2477# 0.08fF
C260 a_n11944_11462# a_n10602_12359# 0.34fF
C261 a_n10992_8440# a_n11283_12359# 0.35fF
C262 a_n10596_8440# fout1 0.03fF
C263 a_n17657_5994# a_n16325_2475# 0.06fF
C264 a_n16976_5994# a_n15981_5897# 0.06fF
C265 a_n2913_2485# a_n2409_2484# 0.02fF
C266 a_n11944_11462# fout2 0.40fF
C267 a_n23808_11542# fout0 1.07fF
C268 a_n10372_2476# modi4 0.02fF
C269 a_n5699_5899# a_n4498_5996# 0.07fF
C270 a_n2614_11550# modi2 0.04fF
C271 a_n17810_11459# a_n15707_12363# 0.06fF
C272 a_n9554_8440# fout1 0.73fF
C273 a_n11793_5995# VDD 1.13fF
C274 a_n24125_2489# fout 0.04fF
C275 a_n5699_5899# fout3 0.84fF
C276 a_n5699_5899# modi4 0.05fF
C277 a_n23172_5903# a_n22746_2481# 0.35fF
C278 a_n15981_5897# fout5 0.86fF
C279 a_n22934_12350# a_n22253_12350# 0.01fF
C280 a_n23595_11454# a_n20815_12350# 0.03fF
C281 a_n22643_8431# a_n21205_8431# 0.09fF
C282 a_n4035_8439# VDD 1.03fF
C283 a_n6140_11462# fout2 1.51fF
C284 a_n3749_8439# a_n4792_8439# 0.07fF
C285 a_n17143_8436# a_n16462_8436# 0.02fF
C286 a_n18023_11547# fout0 0.05fF
C287 a_n10460_2476# a_n11129_2476# 0.06fF
C288 a_n23427_2481# a_n22746_2481# 0.01fF
C289 a_n10117_5898# a_n10372_2476# 0.08fF
C290 a_n4035_8439# modi2 0.06fF
C291 a_n23595_11454# VDD 1.27fF
C292 a_n12508_2484# fout5 0.04fF
C293 a_n19682_2488# modi6 0.10fF
C294 a_n4498_5996# VDD 1.01fF
C295 VDD fin 1.32fF
C296 a_n17143_8436# fout0 0.03fF
C297 a_n11555_5898# fout4 0.82fF
C298 a_n17657_5994# modi5 0.68fF
C299 a_n5187_8439# a_n5478_12358# 0.35fF
C300 a_n11944_11462# a_n11277_8440# 0.09fF
C301 a_n6140_11462# a_n4797_12358# 0.34fF
C302 P1 fout1 0.04fF
C303 modi0 modi1 0.07fF
C304 VDD fout3 5.72fF
C305 a_n6995_11551# modi2 0.09fF
C306 fout2 modi3 0.12fF
C307 VDD modi4 1.37fF
C308 a_n16857_8436# modi0 0.10fF
C309 modi2 fout3 0.60fF
C310 a_n8066_2483# fout4 0.03fF
C311 a_n17419_5897# VDD 1.37fF
C312 a_n21492_12358# modo 0.05fF
C313 a_n14130_2482# modi5 0.12fF
C314 a_n24451_11543# P0 0.02fF
C315 fout6 modi6 2.24fF
C316 a_n17810_11459# VDD 1.30fF
C317 a_n5699_5899# a_n4516_2477# 0.04fF
C318 a_n9159_8440# fout1 0.03fF
C319 a_n11944_11462# a_n9841_12367# 0.06fF
C320 a_n21205_8431# a_n21491_8431# 0.66fF
C321 a_n16976_5994# a_n16219_5994# 0.02fF
C322 a_n15981_5897# a_n16325_2475# 0.85fF
C323 a_n2409_2484# a_n2209_2484# 0.97fF
C324 a_n22247_8431# VDD 1.01fF
C325 a_n4261_5899# fout4 0.23fF
C326 a_n15419_8436# modi1 0.05fF
C327 a_n8769_2484# modi4 0.10fF
C328 a_n5255_5996# a_n4604_2477# 0.12fF
C329 a_n17810_11459# a_n15030_12355# 0.03fF
C330 a_n16857_8436# a_n15419_8436# 0.09fF
C331 a_n17149_12355# a_n16468_12355# 0.01fF
C332 a_n10117_5898# VDD 1.46fF
C333 a_n23172_5903# a_n22728_6000# 0.70fF
C334 a_n5936_5996# fout3 0.04fF
C335 a_n11944_11462# VDD 1.28fF
C336 a_n11555_5898# a_n11793_5995# 0.15fF
C337 a_n16219_5994# fout5 0.02fF
C338 a_n3749_8439# a_n3354_8439# 0.15fF
C339 a_n16462_8436# a_n15705_8436# 0.02fF
C340 a_n9554_8440# modi1 0.81fF
C341 a_n22746_2481# a_n21989_2481# 0.01fF
C342 a_n10460_2476# a_n9691_2476# 0.04fF
C343 a_n10117_5898# a_n8769_2484# 0.04fF
C344 a_n24125_2489# modi 0.07fF
C345 a_n5699_5899# modi3 0.82fF
C346 a_n15705_8436# fout0 0.03fF
C347 a_n6140_11462# VDD 1.27fF
C348 a_n11793_5995# fout4 0.04fF
C349 a_n11944_11462# a_n9840_8440# 0.12fF
C350 a_n15981_5897# modi5 0.11fF
C351 a_n6140_11462# a_n4036_12366# 0.06fF
C352 a_n10992_8440# a_n10596_8440# 0.15fF
C353 a_n17419_5897# a_n18372_2483# 0.06fF
C354 a_n6140_11462# modi2 0.26fF
C355 a_n18023_11547# modi0 0.09fF
C356 a_n20815_12350# modo 0.35fF
C357 a_n17657_5994# VDD 1.10fF
C358 a_n12508_2484# modi5 0.08fF
C359 a_n19682_2488# P7 0.02fF
C360 a_n11283_12359# a_n10602_12359# 0.01fF
C361 a_n10992_8440# a_n9554_8440# 0.09fF
C362 VDD modo 1.03fF
C363 P0 fin 0.65fF
C364 a_n11944_11462# a_n9164_12359# 0.03fF
C365 a_n11555_5898# modi4 0.82fF
C366 a_n15981_5897# a_n15538_5994# 0.69fF
C367 a_n16325_2475# a_n16219_5994# 0.73fF
C368 VDD modi3 1.57fF
C369 a_n20810_8431# VDD 1.07fF
C370 a_n6995_11551# P3 0.02fF
C371 a_n11283_12359# fout2 0.04fF
C372 P3 fout3 0.04fF
C373 modi2 modi3 0.07fF
C374 VDD P5 0.34fF
C375 a_n24451_11543# fin 0.03fF
C376 a_n8066_2483# modi4 0.10fF
C377 a_n5473_8439# fout3 0.03fF
C378 a_n4261_5899# a_n4498_5996# 0.15fF
C379 a_n10355_5995# VDD 1.01fF
C380 fout6 P7 0.41fF
C381 fout3 fout4 2.95fF
C382 a_n23409_6000# a_n22728_6000# 0.02fF
C383 a_n23172_5903# a_n22077_2481# 0.43fF
C384 a_n9159_8440# modi1 0.64fF
C385 a_n14633_2483# fout6 1.07fF
C386 a_n21308_2481# fout 0.04fF
C387 a_n11810_2476# a_n11129_2476# 0.01fF
C388 fout4 modi4 2.14fF
C389 a_n4261_5899# fout3 0.91fF
C390 a_n21734_5903# a_n22746_2481# 0.03fF
C391 a_n22077_2481# a_n23427_2481# 0.03fF
C392 a_n11555_5898# a_n10117_5898# 0.09fF
C393 a_n18465_11548# fout1 0.13fF
C394 a_n22253_12350# a_n21205_8431# 0.04fF
C395 a_n23172_5903# VDD 1.34fF
C396 a_n15705_8436# a_n15024_8436# 0.02fF
C397 a_n5478_12358# fout2 0.03fF
C398 a_n15707_12363# fout0 0.04fF
C399 a_n21989_2481# a_n21308_2481# 0.01fF
C400 a_n9691_2476# fout5 0.04fF
C401 a_n5936_5996# modi3 0.68fF
C402 a_n10117_5898# fout4 0.89fF
C403 a_n6140_11462# a_n3360_12358# 0.03fF
C404 a_n5478_12358# a_n4797_12358# 0.01fF
C405 a_n5187_8439# a_n3749_8439# 0.09fF
C406 a_n17419_5897# a_n16993_2475# 0.35fF
C407 a_n2614_11550# fout3 0.06fF
C408 a_n12600_11551# fout1 0.04fF
C409 a_n16468_12355# modi0 0.02fF
C410 a_n15981_5897# VDD 1.45fF
C411 a_n20070_11542# modo 0.04fF
C412 a_n4604_2477# a_n5273_2477# 0.06fF
C413 a_n4261_5899# a_n4516_2477# 0.08fF
C414 a_n15705_8436# modi0 0.06fF
C415 a_n11793_5995# modi4 0.68fF
C416 a_n16219_5994# a_n15538_5994# 0.02fF
C417 a_n16462_8436# VDD 1.02fF
C418 a_n6140_11462# a_n5473_8439# 0.10fF
C419 a_n22077_2481# fout 0.38fF
C420 a_n23595_11454# fin 1.51fF
C421 a_n4604_2477# a_n3817_5996# 0.11fF
C422 a_n16468_12355# a_n15419_8436# 0.04fF
C423 a_n23409_6000# a_n22077_2481# 0.06fF
C424 a_n22728_6000# a_n21734_5903# 0.06fF
C425 VDD fout0 4.42fF
C426 P0 modo 0.06fF
C427 a_n13930_2482# fout6 0.12fF
C428 a_n19882_2488# fout 0.13fF
C429 a_n11129_2476# a_n10372_2476# 0.01fF
C430 a_n4498_5996# fout3 0.04fF
C431 a_n15419_8436# a_n15705_8436# 0.66fF
C432 fout1 modi1 1.98fF
C433 VDD fout 2.98fF
C434 a_n6995_11551# fout3 0.12fF
C435 a_n11555_5898# a_n10355_5995# 0.07fF
C436 a_n22077_2481# a_n21989_2481# 0.34fF
C437 a_n21734_5903# a_n21308_2481# 0.35fF
C438 a_n21492_12358# a_n21205_8431# 0.33fF
C439 a_n16857_8436# fout1 0.26fF
C440 VDD P4 0.29fF
C441 a_n8066_2483# P5 0.02fF
C442 a_n24451_11543# modo 0.06fF
C443 a_n23409_6000# VDD 1.10fF
C444 fout6 fout5 2.98fF
C445 modi6 P7 0.14fF
C446 modi3 fout4 0.51fF
C447 fout3 modi4 0.13fF
C448 a_n8266_2483# fout5 0.13fF
C449 a_n23595_11454# a_n22247_8431# 0.67fF
C450 a_n22643_8431# a_n22928_8431# 0.66fF
C451 a_n4261_5899# modi3 0.11fF
C452 fout4 P5 0.56fF
C453 a_n22247_8431# fin 0.03fF
C454 a_n10355_5995# fout4 0.04fF
C455 a_n5478_12358# modi2 0.02fF
C456 a_n10992_8440# fout1 0.86fF
C457 a_n15707_12363# modi0 0.05fF
C458 a_n16219_5994# VDD 1.01fF
C459 a_n2913_2485# fout4 1.05fF
C460 a_n22746_2481# fout6 0.04fF
C461 a_n4261_5899# a_n2913_2485# 0.04fF
C462 a_n4604_2477# a_n3835_2477# 0.04fF
C463 a_n10602_12359# a_n9554_8440# 0.04fF
C464 a_n10117_5898# modi4 0.11fF
C465 a_n24251_11543# a_n23808_11542# 0.02fF
C466 a_n2614_11550# modi3 0.07fF
C467 a_n15024_8436# VDD 1.14fF
C468 a_n9554_8440# fout2 0.16fF
C469 a_n5187_8439# a_n4792_8439# 0.15fF
C470 a_n6140_11462# a_n4035_8439# 0.12fF
C471 a_n12600_11551# modi1 0.11fF
C472 a_n16325_2475# fout6 0.49fF
C473 a_n21291_6000# fout 0.03fF
C474 a_n20070_11542# fout0 0.05fF
C475 a_n11555_5898# a_n12508_2484# 0.06fF
C476 a_n15707_12363# a_n15419_8436# 0.33fF
C477 a_n24125_2489# modi6 0.04fF
C478 a_n21734_5903# a_n22077_2481# 0.83fF
C479 a_n22728_6000# a_n21972_6000# 0.02fF
C480 a_n10372_2476# a_n9691_2476# 0.01fF
C481 a_n5954_2477# modi3 0.36fF
C482 a_n6140_11462# fout3 0.44fF
C483 a_n11112_5995# a_n10460_2476# 0.12fF
C484 a_n22077_2481# a_n20386_2489# 0.03fF
C485 a_n21205_8431# a_n20815_12350# 0.08fF
C486 a_n18023_11547# fout1 1.07fF
C487 a_n21734_5903# VDD 1.45fF
C488 a_n23595_11454# modo 0.25fF
C489 a_n3749_8439# fout2 0.74fF
C490 a_n11277_8440# a_n10596_8440# 0.02fF
C491 a_n20386_2489# a_n19882_2488# 0.02fF
C492 a_n21205_8431# VDD 1.34fF
C493 P0 fout0 0.04fF
C494 fin modo 1.14fF
C495 a_n17143_8436# fout1 0.03fF
C496 VDD modi0 1.38fF
C497 a_n23595_11454# a_n20810_8431# 0.06fF
C498 a_n22643_8431# a_n21491_8431# 0.06fF
C499 a_n17419_5897# a_n17657_5994# 0.15fF
C500 VDD modi 0.25fF
C501 fout1 P2 0.67fF
C502 a_n20810_8431# fin 0.03fF
C503 a_n4797_12358# a_n3749_8439# 0.04fF
C504 a_n22728_6000# fout6 0.02fF
C505 fout3 modi3 3.35fF
C506 a_n24451_11543# fout0 0.12fF
C507 a_n16325_2475# a_n17674_2475# 0.03fF
C508 a_n15981_5897# a_n16993_2475# 0.03fF
C509 a_n12157_11550# fout1 0.05fF
C510 a_n18465_11548# a_n18023_11547# 0.02fF
C511 modi6 fout5 0.13fF
C512 a_n15030_12355# modi0 0.35fF
C513 fout6 modi5 0.65fF
C514 modi3 modi4 0.07fF
C515 a_n2209_2484# fout4 0.12fF
C516 a_n21308_2481# fout6 0.03fF
C517 fout4 P4 0.04fF
C518 modi4 P5 0.13fF
C519 a_n15419_8436# VDD 1.40fF
C520 a_n9841_12367# a_n9554_8440# 0.33fF
C521 a_n23595_11454# a_n22934_12350# 0.04fF
C522 a_n22643_8431# a_n23808_11542# 0.04fF
C523 a_n2913_2485# fout3 0.05fF
C524 a_n10596_8440# VDD 1.01fF
C525 a_n10992_8440# modi1 0.10fF
C526 a_n15538_5994# fout6 0.03fF
C527 a_n18665_11548# fout0 0.03fF
C528 a_n22934_12350# fin 0.06fF
C529 a_n11555_5898# a_n11129_2476# 0.35fF
C530 a_n22746_2481# modi6 0.05fF
C531 a_n15419_8436# a_n15030_12355# 0.08fF
C532 a_n22077_2481# a_n21972_6000# 0.71fF
C533 a_n21734_5903# a_n21291_6000# 0.69fF
C534 a_n9554_8440# VDD 1.38fF
C535 a_n4516_2477# modi3 0.02fF
C536 a_n10117_5898# a_n10355_5995# 0.15fF
C537 a_n9554_8440# modi2 0.05fF
C538 a_n21205_8431# a_n20070_11542# 0.06fF
C539 a_n20070_11542# modi0 0.07fF
C540 a_n11129_2476# fout4 0.05fF
C541 a_n21972_6000# VDD 1.02fF
C542 a_n17674_2475# modi5 0.36fF
C543 a_n10596_8440# a_n9840_8440# 0.02fF
C544 a_n19882_2488# a_n19682_2488# 0.97fF
C545 a_n12600_11551# a_n12157_11550# 0.02fF
C546 a_n17419_5897# a_n15981_5897# 0.09fF
C547 a_n3749_8439# VDD 1.32fF
C548 a_n9554_8440# a_n9840_8440# 0.66fF
C549 a_n4036_12366# a_n3749_8439# 0.33fF
C550 a_n22077_2481# fout6 1.38fF
C551 a_n12508_2484# modi4 0.04fF
C552 a_n23595_11454# fout0 0.40fF
C553 a_n3749_8439# modi2 0.80fF
C554 a_n16325_2475# a_n16237_2475# 0.34fF
C555 a_n15981_5897# a_n15556_2475# 0.35fF
C556 a_n5699_5899# a_n5255_5996# 0.70fF
C557 a_n17810_11459# a_n17149_12355# 0.04fF
C558 a_n16857_8436# a_n18023_11547# 0.04fF
C559 a_n14284_11547# modi0 0.04fF
C560 VDD P1 0.33fF
C561 fin fout0 2.82fF
C562 a_n4792_8439# fout2 0.03fF
C563 a_n19882_2488# fout6 0.04fF
C564 a_n14633_2483# a_n13930_2482# 0.02fF
C565 a_n16857_8436# a_n17143_8436# 0.66fF
C566 modi1 P2 0.11fF
C567 a_n17810_11459# a_n16462_8436# 0.67fF
C568 fout1 fout2 2.85fF
C569 a_n9554_8440# a_n9164_12359# 0.08fF
C570 VDD fout6 4.57fF
C571 a_n20810_8431# modo 0.64fF
C572 a_n22728_6000# modi6 0.06fF
C573 a_n22643_8431# a_n22253_12350# 0.08fF
C574 a_n2209_2484# fout3 0.03fF
C575 a_n9159_8440# VDD 1.14fF
C576 a_n12157_11550# modi1 0.09fF
C577 fout6 P6 0.04fF
C578 fout3 P4 0.57fF
C579 modi6 modi5 0.07fF
C580 a_n17810_11459# fout0 1.51fF
C581 a_n14633_2483# fout5 0.05fF
C582 a_n21308_2481# modi6 0.02fF
C583 a_n15419_8436# a_n14284_11547# 0.06fF
C584 a_n5255_5996# VDD 1.02fF
C585 a_n21972_6000# a_n21291_6000# 0.02fF
C586 a_n8769_2484# a_n8266_2483# 0.02fF
C587 a_n6795_11551# a_n6353_11550# 0.02fF
C588 a_n2913_2485# modi3 0.09fF
C589 a_n5478_12358# fout3 0.04fF
C590 a_n10460_2476# a_n9674_5995# 0.11fF
C591 a_n10460_2476# fout5 0.46fF
C592 a_n18665_11548# modi0 0.09fF
C593 a_n9691_2476# fout4 0.05fF
C594 a_n22934_12350# modo 0.02fF
C595 a_n16237_2475# modi5 0.02fF
C596 a_n9840_8440# a_n9159_8440# 0.02fF
C597 a_n5699_5899# a_n6652_2485# 0.06fF
C598 a_n11277_8440# fout1 0.02fF
C599 a_n10992_8440# a_n12157_11550# 0.04fF
C600 a_n11944_11462# a_n11283_12359# 0.04fF
C601 a_n17419_5897# a_n16219_5994# 0.07fF
C602 a_n3749_8439# a_n3360_12358# 0.08fF
C603 a_n12600_11551# fout2 0.13fF
C604 a_n21291_6000# fout6 0.02fF
C605 a_n11129_2476# modi4 0.05fF
C606 a_n16325_2475# a_n14633_2483# 0.03fF
C607 a_n5699_5899# a_n4604_2477# 0.46fF
C608 a_n5936_5996# a_n5255_5996# 0.02fF
C609 a_n9841_12367# fout1 0.05fF
C610 a_n16857_8436# a_n16468_12355# 0.09fF
C611 a_n3354_8439# fout2 0.03fF
C612 a_n18372_2483# fout6 0.06fF
C613 a_n16857_8436# a_n15705_8436# 0.06fF
C614 a_n9554_8440# a_n8419_11550# 0.06fF
C615 a_n17810_11459# a_n15024_8436# 0.06fF
C616 a_n23172_5903# a_n23427_2481# 0.08fF
C617 a_n16976_5994# fout5 0.02fF
C618 a_n22643_8431# a_n21492_12358# 0.03fF
C619 a_n22077_2481# modi6 0.27fF
C620 a_n23595_11454# a_n21205_8431# 0.50fF
C621 a_n4792_8439# VDD 1.03fF
C622 a_n6795_11551# fout2 0.04fF
C623 a_n10602_12359# modi1 0.02fF
C624 a_n10460_2476# a_n11810_2476# 0.03fF
C625 a_n10117_5898# a_n11129_2476# 0.03fF
C626 a_n21205_8431# fin 0.73fF
C627 fin modi0 0.12fF
C628 VDD fout1 4.56fF
C629 modo fout0 0.51fF
C630 a_n13930_2482# fout5 0.03fF
C631 a_n19882_2488# modi6 0.12fF
C632 a_n4604_2477# VDD 1.37fF
C633 fout1 modi2 0.12fF
C634 VDD modi6 1.37fF
C635 modi1 fout2 0.54fF
C636 a_n8266_2483# a_n8066_2483# 0.97fF
C637 a_n5187_8439# a_n6353_11550# 0.04fF
C638 a_n6140_11462# a_n5478_12358# 0.04fF
C639 a_n2209_2484# modi3 0.07fF
C640 a_n9674_5995# fout5 0.03fF
C641 modi3 P4 0.10fF
C642 a_n17810_11459# modi0 0.26fF
C643 a_n8266_2483# fout4 0.04fF
C644 a_n14633_2483# modi5 0.10fF
C645 a_n5699_5899# a_n5273_2477# 0.35fF
C646 a_n21205_8431# a_n22247_8431# 0.07fF
C647 a_n10992_8440# a_n10602_12359# 0.08fF
C648 a_n9840_8440# fout1 0.03fF
C649 a_n16976_5994# a_n16325_2475# 0.12fF
C650 a_n2913_2485# a_n2209_2484# 0.02fF
C651 a_n22928_8431# VDD 0.91fF
C652 a_n10992_8440# fout2 0.25fF
C653 a_n3749_8439# a_n2614_11550# 0.06fF
C654 a_n18665_11548# P1 0.02fF
C655 a_n22934_12350# fout0 0.04fF
C656 a_n23172_5903# fout 0.14fF
C657 a_n9691_2476# modi4 0.02fF
C658 a_n5936_5996# a_n4604_2477# 0.06fF
C659 a_n5255_5996# a_n4261_5899# 0.06fF
C660 a_n17810_11459# a_n15419_8436# 0.43fF
C661 a_n16857_8436# a_n15707_12363# 0.03fF
C662 a_n11112_5995# VDD 1.02fF
C663 a_n23172_5903# a_n23409_6000# 0.15fF
C664 a_n23172_5903# a_n21989_2481# 0.04fF
C665 a_n16325_2475# fout5 1.40fF
C666 a_n3354_8439# VDD 1.07fF
C667 a_n5187_8439# fout2 0.81fF
C668 a_n3749_8439# a_n4035_8439# 0.66fF
C669 a_n9841_12367# modi1 0.05fF
C670 a_n17149_12355# fout0 0.03fF
C671 a_n10460_2476# a_n10372_2476# 0.34fF
C672 a_n10117_5898# a_n9691_2476# 0.35fF
C673 a_n3354_8439# modi2 0.64fF
C674 a_n22643_8431# VDD 1.43fF
C675 a_n18372_2483# modi6 0.07fF
C676 a_n3817_5996# VDD 0.94fF
C677 a_n16462_8436# fout0 0.03fF
C678 a_n5187_8439# a_n4797_12358# 0.08fF
C679 a_n11944_11462# a_n10596_8440# 0.67fF
C680 a_n16976_5994# modi5 0.06fF
C681 a_n10992_8440# a_n11277_8440# 0.66fF
C682 a_n3749_8439# fout3 0.18fF
C683 a_n6795_11551# modi2 0.11fF
C684 a_n14284_11547# fout1 0.05fF
C685 a_n21205_8431# modo 0.81fF
C686 a_n6652_2485# fout4 0.04fF
C687 VDD modi1 1.37fF
C688 a_n13930_2482# modi5 0.10fF
C689 modo modi0 0.07fF
C690 a_n5473_8439# a_n4792_8439# 0.02fF
C691 a_n16857_8436# VDD 1.47fF
C692 a_n17674_2475# a_n16993_2475# 0.01fF
C693 modi1 modi2 0.07fF
C694 VDD P7 0.35fF
C695 P2 fout2 0.04fF
C696 a_n10992_8440# a_n9841_12367# 0.03fF
C697 a_n21205_8431# a_n20810_8431# 0.15fF
C698 a_n11944_11462# a_n9554_8440# 0.50fF
C699 a_n15981_5897# a_n16219_5994# 0.15fF
C700 a_n24451_11543# a_n24251_11543# 0.97fF
C701 a_n4604_2477# fout4 0.39fF
C702 a_n21491_8431# VDD 1.03fF
C703 a_n12157_11550# fout2 1.07fF
C704 fout5 modi5 2.23fF
C705 a_n17419_5897# fout6 0.20fF
C706 a_n2209_2484# P4 0.02fF
C707 a_n8266_2483# modi4 0.12fF
C708 a_n5255_5996# a_n4498_5996# 0.02fF
C709 a_n4261_5899# a_n4604_2477# 0.85fF
C710 a_n10460_2476# VDD 1.40fF
C711 a_n23172_5903# a_n21734_5903# 0.09fF
C712 a_n9840_8440# modi1 0.06fF
C713 a_n15556_2475# fout6 0.04fF
C714 a_n5255_5996# fout3 0.04fF
C715 a_n10992_8440# VDD 1.45fF
C716 a_n11555_5898# a_n11112_5995# 0.70fF
C717 a_n15538_5994# fout5 0.02fF
C718 a_n18665_11548# fout1 0.12fF
C719 a_n22253_12350# a_n21492_12358# 0.01fF
C720 a_n23172_5903# modi 0.05fF
C721 a_n6353_11550# fout2 0.05fF
C722 a_n9164_12359# modi1 0.35fF
.ends

