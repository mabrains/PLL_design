** sch_path: /home/ahmed/PLL_Internship/Ahmed Elshahat LC VCO/CMOS_LC_VCO/CMOS_VCO_tb1.sch
**.subckt CMOS_VCO_tb1

XM1 net2 net2 GND GND sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1

XM2 net1 net2 GND GND sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=50 m=50

XM3 vn vp net1 net1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=43.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3

XM4 vp vn net1 net1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=43.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3

XM5 vn vp VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=30.117 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=30 m=30

XM6 vp vn VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=30.117 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=30 m=30

XM7 V_ctrl vn V_ctrl V_ctrl sky130_fd_pr__nfet_01v8_lvt L=2.7 W=49.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=2

XM8 V_ctrl vp V_ctrl V_ctrl sky130_fd_pr__nfet_01v8_lvt L=2.7 W=49.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=2

*sources
VDD VDD GND V_supply
*I0 VDD net2 dc=5.4m $ideal current source
X1 net2 GND VDD BGR_Banba $non-ideal current source
VTuner V_ctrl GND dc=0.7

*inductor model
L1 vn net3 1.6n m=1
R1 vp net3 1.6 m=1
R2 vp vn 400 m=1
XCF vp vn sky130_fd_pr__cap_mim_m3_1 W=10 L=2.3 MF=1 m=1
XC3 vn GND sky130_fd_pr__cap_mim_m3_1 W=1 L=1.95 MF=1 m=1
XC2 vp GND sky130_fd_pr__cap_mim_m3_1 W=1 L=1.95 MF=1 m=1
*XC_load vp vn sky130_fd_pr__cap_mim_m3_1 W=30 L=38.6 MF=1 m=1

*load cap
C_load vp vn 0.6p m=1


**** begin user architecture code
.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice

* corners parameters
.temp 27
.options tnom=27
.param V_supply = 1.8
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

.subckt BGR_Banba  Iref GND VDD
*.iopin VDD
*.iopin GND
*.opin Iref
XM13 net3 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM14 VBE net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XQ10 GND GND VBE sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ2 GND GND net2 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ3 GND GND net2 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ4 GND GND net2 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ5 GND GND net2 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ6 GND GND net2 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ7 GND GND net2 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ8 GND GND net2 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XQ9 GND GND net2 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XR3 net2 net3 GND sky130_fd_pr__res_xhigh_po_1p41 L=20 mult=1 m=1
XM15 net5 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM16 net1 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=44 m=44
XM17 net6 net3 net5 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6
XM18 net4 VBE net5 VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6
XM19 net1 net6 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
XM20 net6 net4 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM21 net4 net4 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM22 net7 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM23 net7 net1 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=20 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM24 VBE net7 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XR4 GND net3 GND sky130_fd_pr__res_xhigh_po_1p41 L=70 mult=1 m=1
XR5 GND VBE GND sky130_fd_pr__res_xhigh_po_1p41 L=70 mult=1 m=1
XM25 Iref net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=40 m=40
.ends



.GLOBAL GND
.GLOBAL VDD


.save all
.tran 0.01ns 100ns
.control
op
save  @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
 save  @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gm]
 save  @m.xm3.msky130_fd_pr__nfet_01v8_lvt[gm]
 save  @m.xm4.msky130_fd_pr__nfet_01v8_lvt[gm]
 save  @m.xm5.msky130_fd_pr__pfet_01v8_lvt[gm]
 save  @m.xm6.msky130_fd_pr__pfet_01v8_lvt[gm]
 save  @m.xm7.msky130_fd_pr__nfet_01v8_lvt[gm]
 save  @m.xm8.msky130_fd_pr__nfet_01v8_lvt[gm]
 save  @m.x1.xm13.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm14.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm15.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm16.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm17.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm18.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm19.msky130_fd_pr__nfet_g5v0d10v5[gm]
 save  @m.x1.xm20.msky130_fd_pr__nfet_g5v0d10v5[gm]
 save  @m.x1.xm21.msky130_fd_pr__nfet_g5v0d10v5[gm]
 save  @m.x1.xm22.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm23.msky130_fd_pr__nfet_g5v0d10v5[gm]
 save  @m.x1.xm24.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm25.msky130_fd_pr__pfet_g5v0d10v5[gm]
 run
save  @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
 save  @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gm]
 save  @m.xm3.msky130_fd_pr__nfet_01v8_lvt[gm]
 save  @m.xm4.msky130_fd_pr__nfet_01v8_lvt[gm]
 save  @m.xm5.msky130_fd_pr__pfet_01v8_lvt[gm]
 save  @m.xm6.msky130_fd_pr__pfet_01v8_lvt[gm]
 save  @m.xm7.msky130_fd_pr__nfet_01v8_lvt[gm]
 save  @m.xm8.msky130_fd_pr__nfet_01v8_lvt[gm]
 save  @m.x1.xm13.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm14.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm15.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm16.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm17.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm18.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm19.msky130_fd_pr__nfet_g5v0d10v5[gm]
 save  @m.x1.xm20.msky130_fd_pr__nfet_g5v0d10v5[gm]
 save  @m.x1.xm21.msky130_fd_pr__nfet_g5v0d10v5[gm]
 save  @m.x1.xm22.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm23.msky130_fd_pr__nfet_g5v0d10v5[gm]
 save  @m.x1.xm24.msky130_fd_pr__pfet_g5v0d10v5[gm]
 save  @m.x1.xm25.msky130_fd_pr__pfet_g5v0d10v5[gm]
 let vdiff = vp-vn
save vdiff
plot vdiff
linearize vdiff
fft vdiff
wrdata csv_files/gm_xm1.csv tran1.@m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
 wrdata csv_files/gm_xm2.csv tran1.@m.xm2.msky130_fd_pr__nfet_01v8_lvt[gm]
 wrdata csv_files/gm_xm3.csv tran1.@m.xm3.msky130_fd_pr__nfet_01v8_lvt[gm]
 wrdata csv_files/gm_xm4.csv tran1.@m.xm4.msky130_fd_pr__nfet_01v8_lvt[gm]
 wrdata csv_files/gm_xm5.csv tran1.@m.xm5.msky130_fd_pr__pfet_01v8_lvt[gm]
 wrdata csv_files/gm_xm6.csv tran1.@m.xm6.msky130_fd_pr__pfet_01v8_lvt[gm]
 wrdata csv_files/gm_xm7.csv tran1.@m.xm7.msky130_fd_pr__nfet_01v8_lvt[gm]
 wrdata csv_files/gm_xm8.csv tran1.@m.xm8.msky130_fd_pr__nfet_01v8_lvt[gm]
 wrdata csv_files/gm_bgr_banba_xm13.csv tran1.@m.x1.xm13.msky130_fd_pr__pfet_g5v0d10v5[gm]
 wrdata csv_files/gm_bgr_banba_xm14.csv tran1.@m.x1.xm14.msky130_fd_pr__pfet_g5v0d10v5[gm]
 wrdata csv_files/gm_bgr_banba_xm15.csv tran1.@m.x1.xm15.msky130_fd_pr__pfet_g5v0d10v5[gm]
 wrdata csv_files/gm_bgr_banba_xm16.csv tran1.@m.x1.xm16.msky130_fd_pr__pfet_g5v0d10v5[gm]
 wrdata csv_files/gm_bgr_banba_xm17.csv tran1.@m.x1.xm17.msky130_fd_pr__pfet_g5v0d10v5[gm]
 wrdata csv_files/gm_bgr_banba_xm18.csv tran1.@m.x1.xm18.msky130_fd_pr__pfet_g5v0d10v5[gm]
 wrdata csv_files/gm_bgr_banba_xm19.csv tran1.@m.x1.xm19.msky130_fd_pr__nfet_g5v0d10v5[gm]
 wrdata csv_files/gm_bgr_banba_xm20.csv tran1.@m.x1.xm20.msky130_fd_pr__nfet_g5v0d10v5[gm]
 wrdata csv_files/gm_bgr_banba_xm21.csv tran1.@m.x1.xm21.msky130_fd_pr__nfet_g5v0d10v5[gm]
 wrdata csv_files/gm_bgr_banba_xm22.csv tran1.@m.x1.xm22.msky130_fd_pr__pfet_g5v0d10v5[gm]
 wrdata csv_files/gm_bgr_banba_xm23.csv tran1.@m.x1.xm23.msky130_fd_pr__nfet_g5v0d10v5[gm]
 wrdata csv_files/gm_bgr_banba_xm24.csv tran1.@m.x1.xm24.msky130_fd_pr__pfet_g5v0d10v5[gm]
 wrdata csv_files/gm_bgr_banba_xm25.csv tran1.@m.x1.xm25.msky130_fd_pr__pfet_g5v0d10v5[gm]
 plot mag(sp2.vdiff)
wrdata csv_files/vdiff_fft_before_noise.csv mag(sp2.vdiff)
quit
.endc
.end
