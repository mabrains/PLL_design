* Circuit Model for Charge Pump



.subckt charge_pump_behav up dn out vdd gnd +
    voff_up=0.1 von_up=1.7 ron_up=1 roff_up=1Meg i_up=100u +
    voff_dn=0.1 von_dn=1.7 ron_dn=1 roff_dn=1Meg i_dn=100u

    .model cp_switch_up aswitch(cntl_off=voff_up cntl_on=von_up r_off=roff_up r_on=ron_up log=TRUE limit=TRUE)
    .model cp_switch_dn aswitch(cntl_off=voff_dn cntl_on=von_dn r_off=roff_dn r_on=ron_dn log=TRUE limit=TRUE)

    Iup vdd nup_sw i_up
    Aup_sw up %gd(nup_sw out) cp_switch_up
    
    Idn ndn_sw gnd i_dn
    Adn_sw dn %gd(ndn_sw out) cp_switch_dn
.ends