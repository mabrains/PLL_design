* Extracted by KLayout with SKY130 LVS runset on : 07/10/2022 16:21

.SUBCKT TOP
X$1 VDD \$2 via_new$7
X$2 VDD \$2 via_new$2
X$3 VDD \$2 via_new$2
X$4 VDD \$2 via_new$2
X$5 VDD \$2 via_new$2
X$6 VDD \$2 via_new$2
X$7 VDD \$2 via_new$2
X$8 VDD \$2 via_new$2
X$9 net5 \$16 via_new
X$10 net5 \$16 via_new
X$11 \$8 \$15 via_new
X$12 \$8 \$15 via_new
X$13 up \$19 via_new
X$14 up \$19 via_new
X$15 net2 \$20 via_new
X$16 net2 \$20 via_new
X$17 RST via_new$5
X$18 RST via_new$5
X$19 \$47 \$23 via_new$4
X$20 \$47 \$23 via_new$4
X$21 net6 \$52 via_new$2
X$22 net6 \$52 via_new$2
X$23 net3 \$54 via_new$2
X$24 net3 \$54 via_new$2
X$25 \$47 via_new$5
X$26 GND \$57 via_new$6
X$27 GND \$86 via_new$9
X$28 GND \$57 via_new$4
X$29 GND \$86 via_new$2
X$30 GND \$86 via_new$2
X$31 GND \$86 via_new$2
X$32 GND \$86 via_new$2
X$33 GND \$86 via_new$2
X$34 GND \$86 via_new$2
X$35 FB \$56 via_new$3
X$36 FB \$56 via_new$3
X$37 REF \$59 via_new$3
X$38 REF \$59 via_new$3
M$1 \$47 dn_b net7 \$24 sky130_fd_pr__pfet_01v8 L=0.2 W=4 AS=1.16 AD=0.58
+ PS=8.58 PD=4.29
M$2 net7 up_b VDD \$24 sky130_fd_pr__pfet_01v8 L=0.2 W=4 AS=0.58 AD=1.16
+ PS=4.29 PD=8.58
M$3 net1 REF net2 \$71 sky130_fd_pr__pfet_01v8 L=0.2 W=4 AS=1.16 AD=1.16
+ PS=8.58 PD=8.58
M$4 up_b REF net3 \$73 sky130_fd_pr__pfet_01v8 L=0.2 W=4 AS=1.16 AD=1.16
+ PS=8.58 PD=8.58
M$5 net6 FB dn_b \$74 sky130_fd_pr__pfet_01v8 L=0.2 W=4 AS=1.16 AD=1.16 PS=8.58
+ PD=8.58
M$6 net5 FB net4 \$72 sky130_fd_pr__pfet_01v8 L=0.2 W=4 AS=1.16 AD=1.16 PS=8.58
+ PD=8.58
M$7 VDD RST net5 \$28 sky130_fd_pr__pfet_01v8 L=0.15 W=5 AS=1.45 AD=1.45
+ PS=10.58 PD=10.58
M$8 VDD net4 dn_b \$30 sky130_fd_pr__pfet_01v8 L=0.15 W=5 AS=1.45 AD=1.45
+ PS=10.58 PD=10.58
M$9 VDD dn_b \$8 \$34 sky130_fd_pr__pfet_01v8 L=0.15 W=5 AS=1.45 AD=1.45
+ PS=10.58 PD=10.58
M$10 net2 RST VDD \$29 sky130_fd_pr__pfet_01v8 L=0.15 W=5 AS=1.45 AD=1.45
+ PS=10.58 PD=10.58
M$11 up up_b VDD \$38 sky130_fd_pr__pfet_01v8 L=0.15 W=5 AS=1.45 AD=1.45
+ PS=10.58 PD=10.58
M$12 up_b net1 VDD \$35 sky130_fd_pr__pfet_01v8 L=0.15 W=5 AS=1.45 AD=1.45
+ PS=10.58 PD=10.58
M$13 net1 RST GND sky130_gnd sky130_fd_pr__nfet_01v8 L=0.15 W=2.5 AS=0.725
+ AD=0.725 PS=5.58 PD=5.58
M$14 \$47 dn_b GND sky130_gnd sky130_fd_pr__nfet_01v8 L=0.2 W=2 AS=0.58 AD=0.29
+ PS=4.58 PD=2.29
M$15 GND up_b \$47 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.2 W=2 AS=0.29 AD=0.58
+ PS=2.29 PD=4.58
M$16 net6 net4 GND sky130_gnd sky130_fd_pr__nfet_01v8 L=0.15 W=2.5 AS=0.725
+ AD=0.725 PS=5.58 PD=5.58
M$17 GND net1 net3 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.15 W=2.5 AS=0.725
+ AD=0.725 PS=5.58 PD=5.58
M$18 up up_b GND sky130_gnd sky130_fd_pr__nfet_01v8 L=0.15 W=2.5 AS=0.725
+ AD=0.725 PS=5.58 PD=5.58
M$19 GND RST net4 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.15 W=2.5 AS=0.725
+ AD=0.725 PS=5.58 PD=5.58
M$20 GND dn_b \$8 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.15 W=2.5 AS=0.725
+ AD=0.725 PS=5.58 PD=5.58
.ENDS TOP

.SUBCKT via_new$7 \$1 \$4
.ENDS via_new$7

.SUBCKT via_new$9 \$1 \$4
.ENDS via_new$9

.SUBCKT via_new$6 \$1 \$2
.ENDS via_new$6

.SUBCKT via_new$5 \$1
.ENDS via_new$5

.SUBCKT via_new$4 \$1 \$2
.ENDS via_new$4

.SUBCKT via_new$3 \$1 \$2
.ENDS via_new$3

.SUBCKT via_new \$1 \$2
.ENDS via_new

.SUBCKT via_new$2 \$1 \$3
.ENDS via_new$2
