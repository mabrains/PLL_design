** conventional pfd test bench

.include CONV_PFD.ckt
* .lib /open_design_environment/foundry/pdks/skywaters/sky130A/libs.tech/ngspice/sky130.lib.spice "tt"
.lib /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice "tt"
* .Include /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/corners/tt.spice

.temp 27
.options tnom=27
VDD VDD GND 1.8

Xconventional_pfd  REF VDD GND FB up dn conventional_pfd

V4 REF GND pulse(0 1.8 50n 1n 1n 50ns 100ns)
V5 FB GND pulse(0 1.8 0 1n 1n 50ns 100ns)


.control
set wr_singlescale
set wr_vecnames
option numdgt = 3
save all 
print all

tran 0.01ns 400ns 

meas tran tup_check FIND v(up) AT=25n
print tup_check
plot REF FB up dn
wrdata ../csv_files/pfd_ckt{{ corner_string }}.csv v(up) v(dn) v(FB) v(REF)
.endc

.GLOBAL GND
.GLOBAL VDD
.end