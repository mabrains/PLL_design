* NGSPICE file created from vco.ext - technology: sky130A

.subckt cm_p a_2090_700# a_1142_700# a_7462_700# a_6514_700# a_n84_603# a_3670_700#
+ a_2722_700# w_n501_n3475# a_9042_700# a_5250_700# a_4302_700# a_36_700# a_6198_700#
+ a_94_603# a_1458_700# a_6830_700# a_510_700# a_7778_700# a_3986_700# a_3038_700#
+ a_8410_700# a_9594_603# a_9358_700# a_194_700# a_5566_700# a_4618_700# a_1774_700#
+ a_826_700# a_8094_700# a_7146_700# a_3354_700# a_2406_700# a_8726_700# a_5882_700#
+ a_4934_700# VSUBS
X0 a_826_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=5.8e+12p pd=4.058e+07u as=1.508e+14p ps=1.05508e+09u w=2e+07u l=500000u
X1 a_5566_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X2 a_7778_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X3 a_36_700# a_94_603# a_194_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X4 a_36_700# a_94_603# a_1142_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X5 a_94_603# a_94_603# a_3354_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=2.9e+13p pd=2.029e+08u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X6 a_36_700# a_94_603# a_5566_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X7 a_510_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X8 a_5250_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X9 a_7462_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X10 a_94_603# a_94_603# a_7778_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X11 a_36_700# a_94_603# a_7462_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X12 a_36_700# a_94_603# a_5250_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X13 a_7146_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X14 a_36_700# a_94_603# a_2722_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X15 a_36_700# a_94_603# a_4934_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X16 a_9358_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X17 a_36_700# a_94_603# a_7146_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X18 a_194_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X19 a_36_700# a_94_603# a_9358_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X20 a_3038_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X21 a_36_700# a_94_603# a_2406_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X22 a_94_603# a_94_603# a_4618_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X23 a_36_700# a_94_603# a_9042_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X24 a_36_700# a_94_603# a_6830_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X25 a_2722_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X26 a_36_700# a_94_603# a_4302_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X27 a_4934_700# a_94_603# a_94_603# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X28 a_36_700# a_94_603# a_2090_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X29 a_36_700# a_94_603# a_6514_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X30 a_36_700# a_94_603# a_8726_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X31 a_6198_700# a_94_603# a_94_603# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X32 a_2406_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X33 a_4618_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X34 a_6830_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X35 a_9042_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X36 a_36_700# a_94_603# a_3986_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X37 a_36_700# a_94_603# a_6198_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X38 a_2090_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X39 a_36_700# a_94_603# a_8410_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X40 a_4302_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X41 a_6514_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X42 a_8726_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X43 a_36_700# a_94_603# a_8094_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.058e+07u w=2e+07u l=500000u
X44 a_1774_700# a_94_603# a_94_603# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X45 a_3986_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X46 a_8410_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X47 a_36_700# a_94_603# a_826_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X48 a_36_700# a_94_603# a_1774_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X49 a_3670_700# a_94_603# a_94_603# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X50 a_1458_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X51 a_5882_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=5.8e+12p pd=4.058e+07u as=0p ps=0u w=2e+07u l=500000u
X52 a_8094_700# a_94_603# a_94_603# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X53 a_36_700# a_94_603# a_3038_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X54 a_36_700# a_94_603# a_510_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X55 a_94_603# a_94_603# a_1458_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X56 a_94_603# a_94_603# a_5882_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X57 a_1142_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X58 a_3354_700# a_94_603# a_36_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
X59 a_36_700# a_94_603# a_3670_700# w_n501_n3475# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=500000u
C0 a_826_700# a_194_700# 0.12fF
C1 a_3986_700# a_3670_700# 0.23fF
C2 a_1458_700# a_2406_700# 0.09fF
C3 a_9594_603# a_8726_700# 0.07fF
C4 a_8410_700# a_8726_700# 0.23fF
C5 a_94_603# a_1142_700# 0.76fF
C6 w_n501_n3475# a_3986_700# 0.11fF
C7 a_3986_700# a_36_700# 10.75fF
C8 a_3354_700# a_4302_700# 0.09fF
C9 a_2722_700# a_2406_700# 0.23fF
C10 a_1458_700# a_n84_603# 0.01fF
C11 a_4302_700# a_3038_700# 0.05fF
C12 a_1142_700# a_2090_700# 0.09fF
C13 a_8410_700# a_7462_700# 0.09fF
C14 a_6830_700# w_n501_n3475# 0.11fF
C15 a_6830_700# a_36_700# 10.81fF
C16 a_6198_700# a_7146_700# 0.09fF
C17 a_1774_700# a_3038_700# 0.05fF
C18 a_3354_700# a_3038_700# 0.23fF
C19 a_8410_700# a_7778_700# 0.12fF
C20 a_1774_700# a_826_700# 0.09fF
C21 a_194_700# a_510_700# 0.23fF
C22 a_94_603# a_9594_603# 0.04fF
C23 a_7462_700# a_8726_700# 0.05fF
C24 a_5250_700# a_6514_700# 0.05fF
C25 a_8410_700# a_94_603# 0.76fF
C26 a_1142_700# w_n501_n3475# 0.19fF
C27 a_1142_700# a_36_700# 10.83fF
C28 a_7778_700# a_8726_700# 0.09fF
C29 a_94_603# a_8726_700# 0.68fF
C30 a_8094_700# a_7146_700# 0.09fF
C31 a_5250_700# a_3986_700# 0.05fF
C32 a_n84_603# a_194_700# 0.10fF
C33 a_2722_700# a_3986_700# 0.05fF
C34 a_7778_700# a_7462_700# 0.23fF
C35 a_3986_700# a_4934_700# 0.09fF
C36 a_4618_700# a_3986_700# 0.12fF
C37 a_94_603# a_5882_700# 5.84fF
C38 a_1774_700# a_510_700# 0.05fF
C39 a_94_603# a_7462_700# 0.82fF
C40 a_6514_700# a_6198_700# 0.23fF
C41 w_n501_n3475# a_9594_603# 2.32fF
C42 a_9594_603# a_36_700# 0.70fF
C43 a_8410_700# w_n501_n3475# 0.19fF
C44 a_8410_700# a_36_700# 10.83fF
C45 a_6514_700# a_5566_700# 0.09fF
C46 a_826_700# a_510_700# 0.23fF
C47 a_1774_700# a_2406_700# 0.12fF
C48 a_7778_700# a_94_603# 5.76fF
C49 a_3354_700# a_2406_700# 0.09fF
C50 a_1458_700# a_1142_700# 0.23fF
C51 a_2406_700# a_3038_700# 0.12fF
C52 w_n501_n3475# a_8726_700# 0.25fF
C53 a_8726_700# a_36_700# 10.78fF
C54 a_94_603# a_2090_700# 0.82fF
C55 a_826_700# a_n84_603# 0.07fF
C56 a_6830_700# a_6198_700# 0.12fF
C57 w_n501_n3475# a_5882_700# 0.12fF
C58 w_n501_n3475# a_7462_700# 0.11fF
C59 a_36_700# a_5882_700# 5.79fF
C60 a_7462_700# a_36_700# 10.83fF
C61 a_6830_700# a_5566_700# 0.05fF
C62 a_3986_700# a_4302_700# 0.23fF
C63 a_94_603# a_3670_700# 5.84fF
C64 a_7778_700# w_n501_n3475# 0.12fF
C65 a_7778_700# a_36_700# 5.86fF
C66 a_94_603# w_n501_n3475# 28.61fF
C67 a_3354_700# a_3986_700# 0.12fF
C68 a_94_603# a_36_700# 40.39fF
C69 a_1142_700# a_194_700# 0.09fF
C70 a_3986_700# a_3038_700# 0.09fF
C71 a_n84_603# a_510_700# 0.09fF
C72 a_6830_700# a_8094_700# 0.05fF
C73 w_n501_n3475# a_2090_700# 0.11fF
C74 a_9042_700# a_9594_603# 0.09fF
C75 a_2090_700# a_36_700# 10.83fF
C76 a_8410_700# a_9042_700# 0.12fF
C77 a_6514_700# a_7146_700# 0.12fF
C78 a_5250_700# a_5882_700# 0.12fF
C79 a_9042_700# a_8726_700# 0.23fF
C80 w_n501_n3475# a_3670_700# 0.12fF
C81 a_3670_700# a_36_700# 5.79fF
C82 a_9358_700# a_9594_603# 0.10fF
C83 a_1774_700# a_1142_700# 0.12fF
C84 a_1458_700# a_94_603# 5.76fF
C85 a_8410_700# a_9358_700# 0.09fF
C86 a_5882_700# a_4934_700# 0.09fF
C87 w_n501_n3475# a_36_700# 10.64fF
C88 a_4618_700# a_5882_700# 0.05fF
C89 a_5250_700# a_94_603# 0.90fF
C90 a_94_603# a_2722_700# 0.84fF
C91 a_826_700# a_1142_700# 0.23fF
C92 a_6830_700# a_7146_700# 0.23fF
C93 a_1458_700# a_2090_700# 0.12fF
C94 a_9358_700# a_8726_700# 0.12fF
C95 a_94_603# a_4934_700# 5.87fF
C96 a_4618_700# a_94_603# 5.87fF
C97 a_7778_700# a_9042_700# 0.05fF
C98 a_2722_700# a_2090_700# 0.12fF
C99 a_8094_700# a_9594_603# 0.01fF
C100 a_9042_700# a_94_603# 0.57fF
C101 a_8410_700# a_8094_700# 0.23fF
C102 a_6198_700# a_5882_700# 0.23fF
C103 a_6198_700# a_7462_700# 0.05fF
C104 a_5566_700# a_5882_700# 0.23fF
C105 a_1458_700# w_n501_n3475# 0.13fF
C106 a_1458_700# a_36_700# 5.86fF
C107 a_8094_700# a_8726_700# 0.12fF
C108 a_2722_700# a_3670_700# 0.09fF
C109 a_94_603# a_194_700# 0.44fF
C110 a_6198_700# a_94_603# 5.79fF
C111 a_1142_700# a_510_700# 0.12fF
C112 a_5250_700# w_n501_n3475# 0.11fF
C113 a_9358_700# a_94_603# 0.44fF
C114 a_5250_700# a_36_700# 10.75fF
C115 a_94_603# a_5566_700# 0.90fF
C116 w_n501_n3475# a_2722_700# 0.11fF
C117 a_2722_700# a_36_700# 10.81fF
C118 a_3670_700# a_4934_700# 0.05fF
C119 a_4618_700# a_3670_700# 0.09fF
C120 a_1142_700# a_2406_700# 0.05fF
C121 a_8094_700# a_7462_700# 0.12fF
C122 w_n501_n3475# a_4934_700# 0.12fF
C123 a_4618_700# w_n501_n3475# 0.12fF
C124 a_36_700# a_4934_700# 5.76fF
C125 a_4618_700# a_36_700# 5.76fF
C126 a_6830_700# a_6514_700# 0.23fF
C127 a_9042_700# w_n501_n3475# 0.31fF
C128 a_94_603# a_4302_700# 0.90fF
C129 a_8410_700# a_7146_700# 0.05fF
C130 a_9042_700# a_36_700# 10.71fF
C131 a_1142_700# a_n84_603# 0.04fF
C132 a_7778_700# a_8094_700# 0.23fF
C133 a_94_603# a_8094_700# 5.76fF
C134 a_1774_700# a_94_603# 5.76fF
C135 a_3354_700# a_94_603# 5.79fF
C136 w_n501_n3475# a_194_700# 0.31fF
C137 a_194_700# a_36_700# 10.62fF
C138 a_6198_700# w_n501_n3475# 0.12fF
C139 a_94_603# a_3038_700# 0.82fF
C140 a_6198_700# a_36_700# 5.83fF
C141 w_n501_n3475# a_5566_700# 0.11fF
C142 a_1458_700# a_2722_700# 0.05fF
C143 a_9358_700# w_n501_n3475# 0.43fF
C144 a_9358_700# a_36_700# 10.62fF
C145 a_5566_700# a_36_700# 10.75fF
C146 a_94_603# a_826_700# 0.68fF
C147 a_3354_700# a_2090_700# 0.05fF
C148 a_1774_700# a_2090_700# 0.23fF
C149 a_7146_700# a_5882_700# 0.05fF
C150 a_7462_700# a_7146_700# 0.23fF
C151 a_3670_700# a_4302_700# 0.12fF
C152 a_2090_700# a_3038_700# 0.09fF
C153 a_826_700# a_2090_700# 0.05fF
C154 a_5250_700# a_4934_700# 0.23fF
C155 w_n501_n3475# a_4302_700# 0.11fF
C156 a_4618_700# a_5250_700# 0.12fF
C157 a_4302_700# a_36_700# 10.75fF
C158 a_7778_700# a_7146_700# 0.12fF
C159 a_3354_700# a_3670_700# 0.23fF
C160 a_94_603# a_7146_700# 0.84fF
C161 w_n501_n3475# a_8094_700# 0.13fF
C162 a_8094_700# a_36_700# 5.86fF
C163 a_4618_700# a_4934_700# 0.23fF
C164 a_1774_700# w_n501_n3475# 0.12fF
C165 a_3354_700# w_n501_n3475# 0.12fF
C166 a_3354_700# a_36_700# 5.83fF
C167 a_3670_700# a_3038_700# 0.12fF
C168 a_1774_700# a_36_700# 5.86fF
C169 a_1458_700# a_194_700# 0.05fF
C170 a_94_603# a_510_700# 0.57fF
C171 w_n501_n3475# a_3038_700# 0.11fF
C172 a_3038_700# a_36_700# 10.83fF
C173 a_826_700# w_n501_n3475# 0.25fF
C174 a_826_700# a_36_700# 10.78fF
C175 a_5250_700# a_6198_700# 0.09fF
C176 a_5250_700# a_5566_700# 0.23fF
C177 a_94_603# a_2406_700# 0.84fF
C178 a_6198_700# a_4934_700# 0.05fF
C179 a_94_603# a_n84_603# 0.04fF
C180 a_5566_700# a_4934_700# 0.12fF
C181 a_4618_700# a_5566_700# 0.09fF
C182 a_6514_700# a_5882_700# 0.12fF
C183 a_6514_700# a_7462_700# 0.09fF
C184 a_2090_700# a_2406_700# 0.23fF
C185 a_5250_700# a_4302_700# 0.09fF
C186 a_9358_700# a_9042_700# 0.23fF
C187 w_n501_n3475# a_7146_700# 0.11fF
C188 a_7146_700# a_36_700# 10.81fF
C189 a_1458_700# a_1774_700# 0.23fF
C190 a_7778_700# a_6514_700# 0.05fF
C191 a_4302_700# a_4934_700# 0.12fF
C192 w_n501_n3475# a_510_700# 0.28fF
C193 a_4618_700# a_4302_700# 0.23fF
C194 a_6514_700# a_94_603# 0.82fF
C195 a_510_700# a_36_700# 10.71fF
C196 a_3354_700# a_2722_700# 0.12fF
C197 a_1774_700# a_2722_700# 0.09fF
C198 a_1458_700# a_826_700# 0.12fF
C199 a_2406_700# a_3670_700# 0.05fF
C200 a_6198_700# a_5566_700# 0.12fF
C201 a_2722_700# a_3038_700# 0.23fF
C202 a_4618_700# a_3354_700# 0.05fF
C203 w_n501_n3475# a_2406_700# 0.11fF
C204 a_2406_700# a_36_700# 10.81fF
C205 a_6830_700# a_5882_700# 0.09fF
C206 a_9042_700# a_8094_700# 0.09fF
C207 a_6830_700# a_7462_700# 0.12fF
C208 a_94_603# a_3986_700# 0.90fF
C209 w_n501_n3475# a_n84_603# 1.63fF
C210 a_n84_603# a_36_700# 0.70fF
C211 a_6830_700# a_7778_700# 0.09fF
C212 a_5566_700# a_4302_700# 0.05fF
C213 a_6830_700# a_94_603# 0.84fF
C214 a_8410_700# a_9594_603# 0.04fF
C215 a_9358_700# a_8094_700# 0.05fF
C216 a_1458_700# a_510_700# 0.09fF
C217 a_6514_700# w_n501_n3475# 0.11fF
C218 a_6514_700# a_36_700# 10.83fF
C219 a_9358_700# VSUBS -0.17fF
C220 a_9042_700# VSUBS -0.24fF
C221 a_8726_700# VSUBS -0.28fF
C222 a_8410_700# VSUBS -0.29fF
C223 a_8094_700# VSUBS -0.26fF
C224 a_7778_700# VSUBS -0.25fF
C225 a_7462_700# VSUBS -0.25fF
C226 a_7146_700# VSUBS -0.25fF
C227 a_6830_700# VSUBS -0.25fF
C228 a_6514_700# VSUBS -0.25fF
C229 a_6198_700# VSUBS -0.25fF
C230 a_5882_700# VSUBS -0.25fF
C231 a_5566_700# VSUBS -0.25fF
C232 a_5250_700# VSUBS -0.25fF
C233 a_4934_700# VSUBS -0.25fF
C234 a_4618_700# VSUBS -0.25fF
C235 a_4302_700# VSUBS -0.25fF
C236 a_3986_700# VSUBS -0.25fF
C237 a_3670_700# VSUBS -0.25fF
C238 a_3354_700# VSUBS -0.25fF
C239 a_3038_700# VSUBS -0.25fF
C240 a_2722_700# VSUBS -0.25fF
C241 a_2406_700# VSUBS -0.25fF
C242 a_2090_700# VSUBS -0.25fF
C243 a_1774_700# VSUBS -0.25fF
C244 a_1458_700# VSUBS -0.26fF
C245 a_1142_700# VSUBS -0.29fF
C246 a_826_700# VSUBS -0.28fF
C247 a_510_700# VSUBS -0.20fF
C248 a_194_700# VSUBS -0.05fF
C249 a_36_700# VSUBS -5.21fF
C250 a_94_603# VSUBS -0.60fF
C251 a_n84_603# VSUBS 0.70fF
C252 w_n501_n3475# VSUBS 428.25fF
.ends

.subckt cm_n a_2638_n1800# a_1348_n1800# a_258_n1712# a_2122_n1800# a_1606_n1800#
+ a_574_n1800# a_58_n1800# a_3174_n1800# a_2896_n1800# a_0_n1712# a_n220_n1800# m4_n8380_3913#
+ a_832_n1800# a_1548_n1712# a_2380_n1800# a_1864_n1800# a_316_n1800# a_1090_n1800#
+ VSUBS
X0 a_0_n1712# a_316_n1800# a_258_n1712# VSUBS sky130_fd_pr__nfet_01v8 ad=4.35e+13p pd=3.0348e+08u as=4.35e+13p ps=3.0348e+08u w=2.5e+07u l=1e+06u
X1 a_258_n1712# a_2122_n1800# a_0_n1712# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+07u l=1e+06u
X2 a_258_n1712# a_1090_n1800# a_0_n1712# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+07u l=1e+06u
X3 a_258_n1712# a_58_n1800# a_0_n1712# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+07u l=1e+06u
X4 a_0_n1712# a_832_n1800# a_258_n1712# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+07u l=1e+06u
X5 a_0_n1712# a_2896_n1800# a_258_n1712# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+07u l=1e+06u
X6 a_258_n1712# a_2638_n1800# a_0_n1712# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+07u l=1e+06u
X7 a_1548_n1712# a_1348_n1800# a_258_n1712# VSUBS sky130_fd_pr__nfet_01v8 ad=7.25e+12p pd=5.058e+07u as=0p ps=0u w=2.5e+07u l=1e+06u
X8 a_0_n1712# a_1864_n1800# a_258_n1712# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+07u l=1e+06u
X9 a_258_n1712# a_1606_n1800# a_1548_n1712# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+07u l=1e+06u
X10 a_258_n1712# a_574_n1800# a_0_n1712# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+07u l=1e+06u
X11 a_0_n1712# a_2380_n1800# a_258_n1712# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+07u l=1e+06u
C0 a_0_n1712# a_258_n1712# 45.11fF
C1 a_574_n1800# a_0_n1712# 0.80fF
C2 a_58_n1800# a_316_n1800# 0.36fF
C3 a_1090_n1800# a_1348_n1800# 0.36fF
C4 a_2380_n1800# a_0_n1712# 0.80fF
C5 a_832_n1800# a_0_n1712# 0.82fF
C6 a_1864_n1800# a_0_n1712# 0.78fF
C7 a_2638_n1800# a_1548_n1712# 0.11fF
C8 a_2638_n1800# a_258_n1712# 0.64fF
C9 a_n220_n1800# a_0_n1712# 1.34fF
C10 m4_n8380_3913# a_0_n1712# 1.99fF
C11 a_0_n1712# a_3174_n1800# 1.34fF
C12 a_2896_n1800# a_1548_n1712# 0.05fF
C13 a_2638_n1800# a_2380_n1800# 0.36fF
C14 a_2896_n1800# a_258_n1712# 0.53fF
C15 m4_n8380_3913# a_2638_n1800# 0.04fF
C16 a_1548_n1712# a_1090_n1800# 0.23fF
C17 a_58_n1800# a_1548_n1712# 0.05fF
C18 a_1090_n1800# a_258_n1712# 0.88fF
C19 a_58_n1800# a_258_n1712# 0.53fF
C20 a_2896_n1800# m4_n8380_3913# 0.05fF
C21 a_1548_n1712# a_316_n1800# 0.11fF
C22 a_2638_n1800# a_0_n1712# 0.76fF
C23 a_2896_n1800# a_3174_n1800# 0.04fF
C24 a_316_n1800# a_258_n1712# 0.64fF
C25 a_1606_n1800# a_1348_n1800# 0.36fF
C26 a_1548_n1712# a_2122_n1800# 0.20fF
C27 a_1548_n1712# a_1348_n1800# 0.27fF
C28 a_574_n1800# a_316_n1800# 0.36fF
C29 a_832_n1800# a_1090_n1800# 0.36fF
C30 a_2122_n1800# a_258_n1712# 0.82fF
C31 a_1348_n1800# a_258_n1712# 0.92fF
C32 a_2896_n1800# a_0_n1712# 0.74fF
C33 a_58_n1800# a_n220_n1800# 0.04fF
C34 a_2380_n1800# a_2122_n1800# 0.36fF
C35 m4_n8380_3913# a_1090_n1800# 0.04fF
C36 a_58_n1800# m4_n8380_3913# 0.06fF
C37 a_1864_n1800# a_2122_n1800# 0.36fF
C38 m4_n8380_3913# a_316_n1800# 0.04fF
C39 m4_n8380_3913# a_2122_n1800# 0.04fF
C40 m4_n8380_3913# a_1348_n1800# 0.04fF
C41 a_2896_n1800# a_2638_n1800# 0.36fF
C42 a_1090_n1800# a_0_n1712# 0.78fF
C43 a_58_n1800# a_0_n1712# 0.74fF
C44 a_0_n1712# a_316_n1800# 0.76fF
C45 a_1606_n1800# a_1548_n1712# 0.27fF
C46 a_0_n1712# a_2122_n1800# 0.82fF
C47 a_1348_n1800# a_0_n1712# 0.75fF
C48 a_1606_n1800# a_258_n1712# 0.92fF
C49 a_1548_n1712# a_258_n1712# 9.12fF
C50 a_574_n1800# a_1548_n1712# 0.16fF
C51 a_574_n1800# a_258_n1712# 0.73fF
C52 a_2380_n1800# a_1548_n1712# 0.16fF
C53 a_1606_n1800# a_1864_n1800# 0.36fF
C54 a_832_n1800# a_1548_n1712# 0.20fF
C55 a_1864_n1800# a_1548_n1712# 0.23fF
C56 a_2380_n1800# a_258_n1712# 0.73fF
C57 a_832_n1800# a_258_n1712# 0.82fF
C58 a_1864_n1800# a_258_n1712# 0.88fF
C59 a_832_n1800# a_574_n1800# 0.36fF
C60 a_1606_n1800# m4_n8380_3913# 0.04fF
C61 m4_n8380_3913# a_1548_n1712# 0.14fF
C62 a_n220_n1800# a_258_n1712# 0.48fF
C63 m4_n8380_3913# a_258_n1712# 0.09fF
C64 a_574_n1800# m4_n8380_3913# 0.04fF
C65 a_3174_n1800# a_258_n1712# 0.48fF
C66 a_1606_n1800# a_0_n1712# 0.75fF
C67 a_1548_n1712# a_0_n1712# 1.38fF
C68 m4_n8380_3913# a_2380_n1800# 0.04fF
C69 a_832_n1800# m4_n8380_3913# 0.04fF
C70 m4_n8380_3913# a_1864_n1800# 0.04fF
C71 m4_n8380_3913# VSUBS 5.39fF
C72 a_3174_n1800# VSUBS 5.67fF
C73 a_1548_n1712# VSUBS -0.24fF
C74 a_258_n1712# VSUBS 2.69fF
C75 a_0_n1712# VSUBS 8.24fF
C76 a_2896_n1800# VSUBS 0.66fF
C77 a_2638_n1800# VSUBS 0.51fF
C78 a_2380_n1800# VSUBS 0.51fF
C79 a_2122_n1800# VSUBS 0.51fF
C80 a_1864_n1800# VSUBS 0.51fF
C81 a_1606_n1800# VSUBS 0.51fF
C82 a_1348_n1800# VSUBS 0.51fF
C83 a_1090_n1800# VSUBS 0.51fF
C84 a_832_n1800# VSUBS 0.51fF
C85 a_574_n1800# VSUBS 0.51fF
C86 a_316_n1800# VSUBS 0.51fF
C87 a_58_n1800# VSUBS 0.66fF
C88 a_n220_n1800# VSUBS 5.67fF
.ends

.subckt cross_p w_n2129_n555# a_n18_607# a_36_700# a_80_10731# a_1078_600# a_128_700#
+ VSUBS
X0 a_128_700# a_80_10731# a_36_700# w_n2129_n555# sky130_fd_pr__pfet_01v8 ad=8.25e+13p pd=5.033e+08u as=4.85e+13p ps=3.0194e+08u w=5e+07u l=150000u
X1 a_128_700# a_36_700# a_80_10731# w_n2129_n555# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.85e+13p ps=3.0194e+08u w=5e+07u l=150000u
X2 a_80_10731# a_36_700# a_128_700# w_n2129_n555# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=150000u
X3 a_36_700# a_80_10731# a_128_700# w_n2129_n555# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=150000u
X4 a_128_700# a_80_10731# a_36_700# w_n2129_n555# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=150000u
X5 a_128_700# a_36_700# a_80_10731# w_n2129_n555# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=150000u
X6 a_36_700# a_80_10731# a_128_700# w_n2129_n555# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=150000u
X7 a_80_10731# a_36_700# a_128_700# w_n2129_n555# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=150000u
X8 a_80_10731# a_36_700# a_128_700# w_n2129_n555# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=150000u
X9 a_128_700# a_80_10731# a_36_700# w_n2129_n555# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+07u l=150000u
C0 a_36_700# a_80_10731# 3.38fF
C1 a_n18_607# a_128_700# 0.49fF
C2 a_128_700# w_n2129_n555# 5.00fF
C3 a_n18_607# w_n2129_n555# 5.58fF
C4 a_1078_600# a_36_700# 0.34fF
C5 a_36_700# a_128_700# 54.63fF
C6 a_n18_607# a_36_700# 0.52fF
C7 a_36_700# w_n2129_n555# 9.69fF
C8 a_1078_600# a_80_10731# 0.53fF
C9 a_80_10731# a_128_700# 38.95fF
C10 a_n18_607# a_80_10731# 0.38fF
C11 a_80_10731# w_n2129_n555# 9.33fF
C12 a_1078_600# a_128_700# 0.52fF
C13 a_1078_600# a_n18_607# 0.15fF
C14 a_1078_600# w_n2129_n555# 5.58fF
C15 a_1078_600# VSUBS 0.03fF
C16 a_128_700# VSUBS -0.58fF
C17 a_36_700# VSUBS 1.79fF
C18 a_80_10731# VSUBS 1.83fF
C19 a_n18_607# VSUBS 0.03fF
C20 w_n2129_n555# VSUBS 181.15fF
.ends

.subckt cap m3_0_0# c1_100_100# VSUBS
X0 c1_100_100# m3_0_0# sky130_fd_pr__cap_mim_m3_1 l=1.3e+07u w=1.4e+07u
C0 c1_100_100# m3_0_0# 15.76fF
C1 c1_100_100# VSUBS 1.31fF
C2 m3_0_0# VSUBS 5.64fF
.ends

.subckt var a_n48_0# a_1610_0# a_n106_88# VSUBS
X0 a_n106_88# a_n48_0# a_n106_88# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.479e+13p pd=1.0374e+08u as=0p ps=0u w=1.7e+07u l=8e+06u
X1 a_n106_88# a_1610_0# a_n106_88# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.7e+07u l=8e+06u
C0 a_1610_0# a_n48_0# 0.39fF
C1 a_1610_0# a_n106_88# 11.26fF
C2 a_n106_88# a_n48_0# 8.80fF
C3 a_n106_88# VSUBS 7.55fF
C4 a_1610_0# VSUBS 4.90fF
C5 a_n48_0# VSUBS 4.73fF
.ends

.subckt cross_n a_92_n512# a_1042_n600# a_0_n512# a_n54_n600# a_44_3510# VSUBS
X0 a_0_n512# a_44_3510# a_92_n512# VSUBS sky130_fd_pr__nfet_01v8 ad=1.94e+13p pd=1.2194e+08u as=3.3e+13p ps=2.033e+08u w=2e+07u l=150000u
X1 a_92_n512# a_0_n512# a_44_3510# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.94e+13p ps=1.2194e+08u w=2e+07u l=150000u
X2 a_44_3510# a_0_n512# a_92_n512# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X3 a_92_n512# a_44_3510# a_0_n512# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X4 a_44_3510# a_0_n512# a_92_n512# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X5 a_92_n512# a_44_3510# a_0_n512# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X6 a_92_n512# a_44_3510# a_0_n512# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X7 a_0_n512# a_44_3510# a_92_n512# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X8 a_92_n512# a_0_n512# a_44_3510# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
X9 a_44_3510# a_0_n512# a_92_n512# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+07u l=150000u
C0 a_92_n512# a_0_n512# 26.69fF
C1 a_44_3510# a_1042_n600# 0.23fF
C2 a_1042_n600# a_n54_n600# 0.06fF
C3 a_44_3510# a_n54_n600# 0.18fF
C4 a_92_n512# a_1042_n600# 0.22fF
C5 a_44_3510# a_92_n512# 16.08fF
C6 a_92_n512# a_n54_n600# 0.21fF
C7 a_0_n512# a_1042_n600# 0.15fF
C8 a_44_3510# a_0_n512# 1.88fF
C9 a_0_n512# a_n54_n600# 0.22fF
C10 a_1042_n600# VSUBS 2.61fF
C11 a_92_n512# VSUBS 3.47fF
C12 a_0_n512# VSUBS 8.23fF
C13 a_44_3510# VSUBS 7.36fF
C14 a_n54_n600# VSUBS 2.61fF
.ends

.subckt vco VDD GND vp vn ibias vctrl net2 net1
Xcm_p_0 VDD VDD VDD VDD cm_p_0/a_n84_603# VDD VDD VDD VDD VDD VDD net2 VDD net1 VDD
+ VDD VDD VDD VDD VDD VDD cm_p_0/a_9594_603# VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD
+ VDD VDD VDD GND cm_p
Xcm_n_0 ibias ibias GND ibias ibias ibias ibias cm_n_0/a_3174_n1800# ibias net1 cm_n_0/a_n220_n1800#
+ ibias ibias ibias ibias ibias ibias ibias GND cm_n
Xcross_p_0 net2 cross_p_0/a_n18_607# vp vn cross_p_0/a_1078_600# net2 GND cross_p
Xcap_0 vn vp GND cap
Xvar_0 vn vp vctrl GND var
Xcross_n_0 GND cross_n_0/a_1042_n600# vp cross_n_0/a_n54_n600# vn GND cross_n
C0 net1 ibias 0.85fF
C1 vn vp 21.59fF
C2 net1 vp 2.67fF
C3 vp cross_n_0/a_n54_n600# -0.07fF
C4 net1 vn 5.17fF
C5 vn cross_n_0/a_n54_n600# -0.02fF
C6 cm_p_0/a_n84_603# VDD 0.09fF
C7 net2 cross_p_0/a_n18_607# 1.64fF
C8 net2 VDD 6.56fF
C9 vn cross_n_0/a_1042_n600# -0.07fF
C10 vp vctrl 0.67fF
C11 net1 cm_n_0/a_n220_n1800# -0.69fF
C12 net1 cm_n_0/a_3174_n1800# -0.69fF
C13 vp cross_p_0/a_n18_607# -0.18fF
C14 vp VDD 0.13fF
C15 net2 cross_p_0/a_1078_600# 1.63fF
C16 vn cross_p_0/a_n18_607# -0.04fF
C17 net2 vp 4.67fF
C18 vn VDD 1.17fF
C19 net2 vn 18.15fF
C20 net1 VDD 18.58fF
C21 net2 net1 0.62fF
C22 cm_p_0/a_9594_603# VDD 0.10fF
C23 vn ibias 0.85fF
C24 cross_p_0/a_1078_600# vp -0.02fF
C25 cross_p_0/a_1078_600# vn -0.17fF
C26 VDD GND 669.20fF
C27 net2 GND 240.85fF
C28 cross_n_0/a_1042_n600# GND 3.26fF
C29 vn GND 99.84fF
C30 cross_n_0/a_n54_n600# GND 3.27fF
C31 vctrl GND 15.49fF
C32 vp GND 85.13fF
C33 cross_p_0/a_1078_600# GND 0.03fF
C34 cross_p_0/a_n18_607# GND 0.03fF
C35 cm_n_0/a_3174_n1800# GND 6.55fF
C36 net1 GND 26.70fF
C37 ibias GND 24.19fF
C38 cm_n_0/a_n220_n1800# GND 6.55fF
C39 cm_p_0/a_n84_603# GND 0.70fF
.ends

