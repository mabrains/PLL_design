
 V1 net8 vp DC 0 trnoise (6.949344748800417e-10 0.03n 1 6.949344748800417e-10)
 V2 net7 vn DC 0 trnoise (5.810405225373581e-10 0.03n 1 5.810405225373582e-10)
 V4 net3 net2 DC 0 trnoise (8.140844938214757e-10 0.03n 1 8.140844938214759e-10)
 V5 net5 net2 DC 0 trnoise (7.164133635857781e-10 0.03n 1 7.164133635857781e-10)
 V7 net6 vp DC 0 trnoise (5.835983832218721e-10 0.03n 1 5.835983832218721e-10)
 V11 net9 vn DC 0 trnoise (6.908184444313312e-10 0.03n 1 6.908184444313311e-10)
 V3 net11 vp DC 0 trnoise (0 0 0 0)
 V10 net10 vn DC 0 trnoise (0 0 0 0)
 VR1 net12 vp DC 0 trnoise (4.424242308011621e-09 0.03n 0 0)
VR2 net13 net14 DC 0 trnoise (2.228901074520805e-10 0.03n 0 0)

 V1 net8 vp DC 0 trnoise (6.835090128649205e-10 0.03n 1 6.835090128649205e-10)
 V2 net7 vn DC 0 trnoise (5.785427398132504e-10 0.03n 1 5.785427398132504e-10)
 V4 net3 net2 DC 0 trnoise (7.927040635837875e-10 0.03n 1 7.927040635837876e-10)
 V5 net5 net2 DC 0 trnoise (7.158307893455211e-10 0.03n 1 7.158307893455212e-10)
 V7 net6 vp DC 0 trnoise (5.615748424773629e-10 0.03n 1 5.615748424773628e-10)
 V11 net9 vn DC 0 trnoise (6.874629010540658e-10 0.03n 1 6.874629010540658e-10)
 V3 net11 vp DC 0 trnoise (0 0 0 0)
 V10 net10 vn DC 0 trnoise (0 0 0 0)
 VR1 net12 vp DC 0 trnoise (4.424242308011621e-09 0.03n 0 0)
VR2 net13 net14 DC 0 trnoise (2.228901074520805e-10 0.03n 0 0)


** sch_path: /home/ahmed/Mabrains_internship/VCO_Try1/VCO_try7.sch
**.subckt VCO_try7
XM11 vp net9 net1 net1 sky130_fd_pr__pfet_01v8 L=0.15 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
XM1 vn net8 net1 net1 sky130_fd_pr__pfet_01v8 L=0.15 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
XM2 vp net7 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
L1 vp net14 4n m=1
I0 net2 GND 5m
R1 net12 vn 1182 m=1
VDD VDD GND 1.8
R2 net13 vn 3 m=1
XM4 net1 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
XM5 net2 net5 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
XM7 vn net6 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
C1 vp vn 5f m=10
C3 vp GND 5f m=5
C2 vn GND 5f m=5
Vctrl net4 GND 1.7
XM10 net4 net10 net4 GND sky130_fd_pr__pfet_01v8_lvt L=1.3 W=12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
XM3 net4 net11 net4 GND sky130_fd_pr__pfet_01v8_lvt L=1.3 W=12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
C13 vp vn 10f m=10

**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foundry/pdks/skywaters/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


.tran 0.04n 200u
.save all
.control
  run

 
  let vdiff = v(vp)-v(vn)
  save vdiff
  *plot vdiff
  linearize vdiff
  *save vdiff
  *fft (v(vp)-v(vn))
  fft vdiff
  *spec 0.5 1.5e9 210e3 vout
  
 


  plot mag(sp2.vdiff)
  wrdata vdiff_fft.csv mag(sp2.vdiff)
  
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
