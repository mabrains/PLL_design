** Test bench for ring

.include ../spice_files/ring_cir.ckt


.lib /foundry/pdks/skywaters/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice ff
.temp 125.00
.options tnom=125.00
VDD VDD GND 1.62

xring Vin out VDD GND ring

**** begin user architecture code

.control

    op 
    save all
        
    print all

    tran 2ns 5us uic
    plot out
    meas tran tperiod TRIG out VAL=0.4 RISE=15 TARG out VAL=0.4 RISE=16
    let freq = 1/(tperiod*1000000)
    print freq
    
.endc

.GLOBAL GND
.GLOBAL VDD
.end