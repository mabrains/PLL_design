* NGSPICE file created from c2.ext - technology: sky130A


* Top level circuit c2

X0 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X1 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X2 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X3 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X4 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X5 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X6 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X7 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X8 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X9 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X10 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X11 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X12 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X13 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X14 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X15 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X16 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X17 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X18 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X19 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X20 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X21 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X22 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X23 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X24 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X25 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X26 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X27 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X28 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X29 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X30 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X31 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X32 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X33 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X34 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X35 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X36 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X37 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X38 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X39 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X40 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X41 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X42 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X43 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X44 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X45 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X46 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X47 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X48 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X49 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X50 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X51 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X52 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X53 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X54 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X55 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X56 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X57 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X58 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X59 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X60 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X61 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X62 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X63 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X64 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X65 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X66 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X67 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X68 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X69 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X70 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X71 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X72 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X73 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X74 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X75 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X76 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X77 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X78 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X79 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X80 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X81 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X82 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X83 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X84 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X85 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X86 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X87 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X88 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X89 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X90 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X91 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X92 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X93 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X94 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X95 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X96 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X97 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X98 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X99 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X100 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X101 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X102 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X103 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X104 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X105 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X106 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X107 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X108 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X109 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X110 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X111 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X112 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X113 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X114 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X115 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X116 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X117 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X118 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X119 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X120 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X121 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X122 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X123 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X124 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X125 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X126 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X127 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X128 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X129 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X130 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X131 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X132 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X133 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X134 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X135 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X136 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X137 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X138 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X139 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X140 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X141 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X142 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X143 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X144 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X145 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X146 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X147 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X148 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X149 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X150 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X151 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X152 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X153 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X154 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X155 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X156 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X157 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X158 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X159 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X160 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X161 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X162 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X163 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X164 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X165 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X166 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X167 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X168 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X169 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X170 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X171 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X172 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X173 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X174 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X175 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X176 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X177 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X178 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X179 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X180 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X181 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X182 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X183 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X184 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X185 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X186 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X187 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X188 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X189 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X190 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X191 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X192 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X193 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X194 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X195 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X196 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X197 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X198 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X199 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X200 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X201 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X202 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X203 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X204 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X205 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X206 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X207 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X208 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X209 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X210 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X211 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X212 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X213 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X214 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X215 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X216 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X217 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X218 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X219 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X220 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X221 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X222 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X223 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X224 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X225 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X226 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X227 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X228 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X229 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X230 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X231 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X232 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X233 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X234 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X235 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X236 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X237 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X238 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X239 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X240 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X241 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X242 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X243 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X244 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X245 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X246 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X247 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X248 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X249 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X250 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X251 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X252 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X253 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X254 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X255 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X256 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X257 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X258 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X259 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X260 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X261 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X262 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X263 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X264 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X265 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X266 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X267 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X268 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X269 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X270 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X271 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X272 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X273 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X274 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X275 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X276 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X277 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X278 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X279 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X280 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X281 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X282 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X283 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X284 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X285 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X286 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X287 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X288 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X289 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X290 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X291 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X292 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X293 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X294 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X295 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X296 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X297 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X298 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X299 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X300 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X301 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X302 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X303 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X304 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X305 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X306 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X307 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X308 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X309 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X310 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X311 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X312 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X313 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X314 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X315 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X316 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X317 m3_51_6723 m3_n2557_n3135 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X318 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
X319 m3_n2557_n3135 m3_51_6723 sky130_fd_pr__cap_mim_m3_1 l=2.788e+07u w=2.787e+07u
.end

