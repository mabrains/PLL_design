** Test bench for BGR

.include ../spice_files/BGR_cir.ckt


.lib /open_design_environment/foundry/pdks/skywaters/sky130A/libs.tech/ngspice/sky130.lib.spice ss
.temp 50.00
.options tnom=50.00

VDD VDD GND 1.62
VTuner out GND 0.90


xvco out GND VDD BGR_Banba

**** begin user architecture code

.control
    set wr_singlescale
    set wr_vecnames
    set appendwrite

    op
    let Iref = i(VTuner)*1000000
    print Iref
    print all

   
    
.endc

.GLOBAL GND
.GLOBAL VDD
.end