* NGSPICE file created from DIV_CELL.ext - technology: sky130A

.subckt DIV_CELL fin P modo net1 net1_nand3 net2 net2_nand3 net1_ff1 net2_ff1 net4_ff1
+ net5_ff1 net4_ff2 net2_ff2 net5_ff2 2 1 3 modi fout 31 finb net3_ff1 net3_ff2 VDD
+ GND
X0 VDD 2 fout VDD sky130_fd_pr__pfet_01v8 ad=1.508e+13p pd=1.1154e+08u as=2.32e+12p ps=1.716e+07u w=4 l=0.15
X1 net1_ff1 fout VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u w=4 l=0.15
X2 GND modo net2_nand3 GND sky130_fd_pr__nfet_01v8 ad=8.7e+12p pd=6.522e+07u as=3.48e+12p ps=2.516e+07u w=6 l=0.15
X3 net2 modi 31 GND sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=1.74e+12p ps=1.258e+07u w=6 l=0.15
X4 net4_ff1 net3_ff1 VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=1.716e+07u as=0p ps=0u w=4 l=0.15
X5 net1_nand3 P 2 GND sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=1.74e+12p ps=1.258e+07u w=6 l=0.15
X6 net5_ff2 net3_ff2 GND GND sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2 l=0.15
X7 GND 31 3 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2 l=0.15
X8 net3_ff1 finb net1_ff1 VDD sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4 l=0.15
X9 VDD modi 31 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.32e+12p ps=1.716e+07u w=4 l=0.15
X10 net1 2 fout GND sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=2.516e+07u as=1.74e+12p ps=1.258e+07u w=6 l=0.15
X11 GND fin finb GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2 l=0.15
X12 VDD 1 fout VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4 l=0.15
X13 net3_ff1 fin net2_ff1 GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=1.16e+12p ps=9.16e+06u w=2 l=0.15
X14 modo finb net5_ff2 GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2 l=0.15
X15 VDD fin 2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.48e+12p ps=2.574e+07u w=4 l=0.15
X16 GND 1 net1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6 l=0.15
X17 modo fin net4_ff2 VDD sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=4.64e+12p ps=3.432e+07u w=4 l=0.15
X18 net3_ff2 fin net2_ff2 GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=1.16e+12p ps=9.16e+06u w=2 l=0.15
X19 1 fin net4_ff1 VDD sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4 l=0.15
X20 net2_ff1 fout GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2 l=0.15
X21 GND fout net2 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6 l=0.15
X22 1 finb net5_ff1 GND sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=1.16e+12p ps=9.16e+06u w=2 l=0.15
X23 net2_nand3 fin net1_nand3 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6 l=0.15
X24 net5_ff1 net3_ff1 GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2 l=0.15
X25 net3_ff2 finb net4_ff2 VDD sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4 l=0.15
X26 finb fin VDD VDD sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4 l=0.15
X27 net4_ff2 net3_ff2 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4 l=0.15
X28 VDD modo 2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4 l=0.15
X29 net4_ff2 3 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4 l=0.15
X30 net2_ff2 3 GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2 l=0.15
X31 VDD P 2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4 l=0.15
X32 VDD fout 31 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4 l=0.15
X33 3 31 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4 l=0.15
C0 net3_ff1 2 0.02fF
C1 net4_ff2 1 0.18fF
C2 fin fout 2.86fF
C3 net4_ff1 net3_ff2 0.07fF
C4 finb net2_nand3 0.05fF
C5 modo net5_ff1 0.02fF
C6 finb 31 0.18fF
C7 net3_ff1 net4_ff2 0.06fF
C8 fin 3 0.37fF
C9 fin net1_ff1 0.03fF
C10 finb modi 0.14fF
C11 P VDD 0.27fF
C12 fin 1 1.54fF
C13 P fout 0.09fF
C14 finb net2 0.01fF
C15 fin net3_ff1 0.90fF
C16 net4_ff2 net3_ff2 0.81fF
C17 P 1 0.01fF
C18 modo VDD 0.90fF
C19 modo fout 0.51fF
C20 net1 net2_nand3 0.02fF
C21 fin net3_ff2 0.76fF
C22 finb net2_ff2 0.01fF
C23 modo 3 0.53fF
C24 modo 1 0.25fF
C25 finb net2_ff1 0.07fF
C26 net5_ff1 1 0.34fF
C27 net2_nand3 net1_nand3 0.97fF
C28 modo net3_ff1 0.10fF
C29 net2_nand3 2 0.12fF
C30 net3_ff1 net5_ff1 0.08fF
C31 VDD fout 3.21fF
C32 VDD 3 1.67fF
C33 VDD net1_ff1 0.91fF
C34 modo net3_ff2 0.81fF
C35 net4_ff2 31 0.05fF
C36 VDD 1 1.24fF
C37 fout 3 1.06fF
C38 net1_ff1 fout 0.03fF
C39 net5_ff1 net3_ff2 0.04fF
C40 1 fout 0.41fF
C41 fin net2_nand3 0.04fF
C42 net3_ff1 VDD 1.34fF
C43 fin 31 0.17fF
C44 1 3 0.09fF
C45 net1_ff1 1 0.09fF
C46 fin modi 0.12fF
C47 net3_ff1 fout 0.25fF
C48 modo net5_ff2 0.35fF
C49 net3_ff1 3 0.05fF
C50 net3_ff1 net1_ff1 0.66fF
C51 VDD net3_ff2 1.31fF
C52 net3_ff1 1 0.85fF
C53 fout net3_ff2 0.16fF
C54 net1 finb 0.08fF
C55 net3_ff2 3 0.22fF
C56 modo net2_nand3 0.09fF
C57 1 net3_ff2 0.50fF
C58 fin net2_ff2 0.05fF
C59 modo 31 1.43fF
C60 finb net4_ff1 0.06fF
C61 modo modi 0.06fF
C62 net3_ff1 net3_ff2 0.09fF
C63 fin net2_ff1 0.06fF
C64 finb net1_nand3 0.04fF
C65 net5_ff2 3 0.03fF
C66 modo net2 0.04fF
C67 finb 2 0.20fF
C68 net5_ff2 1 0.03fF
C69 finb net4_ff2 0.01fF
C70 net2_nand3 fout 0.13fF
C71 VDD 31 2.52fF
C72 VDD modi 0.24fF
C73 modo net2_ff2 0.05fF
C74 31 fout 1.16fF
C75 fout modi 0.96fF
C76 finb fin 2.10fF
C77 net5_ff1 net2_ff2 0.01fF
C78 31 3 1.51fF
C79 modo net2_ff1 0.02fF
C80 net5_ff2 net3_ff2 0.08fF
C81 modi 3 0.74fF
C82 net1 net1_nand3 0.02fF
C83 net1 2 0.13fF
C84 fout net2 0.05fF
C85 net2_ff1 net5_ff1 0.01fF
C86 finb P 0.04fF
C87 net2 3 0.11fF
C88 net4_ff2 net4_ff1 0.02fF
C89 net1_nand3 2 1.00fF
C90 modo finb 0.74fF
C91 net1 fin 0.05fF
C92 31 net3_ff2 0.19fF
C93 modi net3_ff2 0.05fF
C94 net2_ff2 3 0.01fF
C95 net2_ff1 fout 0.04fF
C96 finb net5_ff1 0.05fF
C97 1 net2_ff2 0.06fF
C98 fin net4_ff1 0.04fF
C99 net2 net3_ff2 0.06fF
C100 net2_ff1 1 0.04fF
C101 net3_ff1 net2_ff2 0.03fF
C102 fin net1_nand3 0.03fF
C103 31 net5_ff2 0.03fF
C104 fin 2 0.60fF
C105 net2_ff1 net3_ff1 0.35fF
C106 finb VDD 2.31fF
C107 fin net4_ff2 0.08fF
C108 net3_ff2 net2_ff2 0.33fF
C109 net1 modo 0.08fF
C110 P net1_nand3 0.03fF
C111 finb fout 2.72fF
C112 P 2 0.40fF
C113 finb 3 0.79fF
C114 finb net1_ff1 0.12fF
C115 finb 1 0.62fF
C116 31 modi 0.46fF
C117 modo net1_nand3 0.07fF
C118 net5_ff2 net2_ff2 0.01fF
C119 finb net3_ff1 0.88fF
C120 modo 2 0.80fF
C121 fin P 0.89fF
C122 31 net2 1.06fF
C123 modi net2 0.06fF
C124 modo net4_ff2 0.71fF
C125 net1 fout 1.07fF
C126 VDD net4_ff1 1.01fF
C127 finb net3_ff2 0.45fF
C128 net1 1 0.03fF
C129 modo fin 1.17fF
C130 31 net2_ff2 0.01fF
C131 net1_ff1 net4_ff1 0.02fF
C132 VDD 2 4.59fF
C133 net1_nand3 fout 0.12fF
C134 1 net4_ff1 0.67fF
C135 net1 net3_ff1 0.04fF
C136 2 fout 0.84fF
C137 finb net5_ff2 0.02fF
C138 VDD net4_ff2 2.02fF
C139 modo P 0.56fF
C140 net3_ff1 net4_ff1 0.15fF
C141 2 1 0.44fF
C142 net4_ff2 3 0.08fF
C143 fin VDD 1.51fF
.ends
