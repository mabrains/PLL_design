*VCO*behave

.subckt VCO CtrL_Signal OUT

	* Maybe needs an array parsing with too many values 
    asine CtrL_Signal OUT in_sine
    .model in_sine sine(cntl_array = [0.3 0.5 0.7 1.3]
    + freq_array=[2.4e9 2.43e9 2.46e9 2.48e9] out_low = -1.8
    + out_high = 1.8)
    
.ends VCO
