** Test bench for VCO

.include ../spice_files/vco_cir.ckt

{{ corner_setup }}

xvco vp vn vctrl ibias VDD GND vco

**** begin user architecture code

.control
    set wr_singlescale
    set wr_vecnames
    set appendwrite

    op
    print all

    ** tran 0.01ns 100ns
    ** let vdiff = v(vp)-v(vn)
    ** let vdiff_max =  vecmax(vp-vn)
    ** meas tran tperiod TRIG vdiff VAL=0.4 RISE=30 TARG vdiff VAL=0.4 RISE=31
    ** let freq = 1/tperiod
    ** print(freq)
.endc

.GLOBAL GND
.GLOBAL VDD
.end
