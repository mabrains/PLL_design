** sch_path: /home/mohammed/Desktop/RO/untitled.sch
**.subckt untitled
**.ends
.end
