* PLL subckt

.include ../../PFD/circuit/pfd_cir.ckt
.include ../../CP/circuit/cp_cir.ckt
.include ../../VCO/circuit/vco_sch.ckt
.include ../../VCO/circuit/inductor_model_cct.ckt
.include ../../VCO/circuit/vco_inverter.ckt
.include ../../BGR/circuit/bgr_sch.ckt
.include ../../LPF/circuit/lf_cir.ckt
.include ../../Divider/circuit/divider.ckt

.subckt pll ref p0 p1 p2 p3 p4 p5 p6 p7 vco_out VDD GND

Xconventional_pfd  ref VDD GND fb up dn conventional_pfd
Xcp up lf_input dn VDD GND CP_with_buffer 
Xloop_filter_3rd_order lf_input vctrl GND loop_filter_3rd_order 
*************************VCO********************
xvco vp vn vctrl ibias VDD GND vco_sch
xind1 vp vn ind_model
XC_load vp vn sky130_fd_pr__cap_mim_m3_1 W=13 L=9 MF=1 m=1  $mim cap
xbgr ibias GND VDD bgr_sch
** Isource VDD ibias 90u
xinverter vp vco_out VDD GND vco_inverter     w_p=60 w_n=4.2 l=0.15
xinverter2 vn fout_dummy VDD GND vco_inverter w_p=60 w_n=4.2 l=0.15
*************************************************
xdivider VDD fb GND p2 p7 p1 p6 p5 p4 p3 p0 vco_out float divider

.ends
.GLOBAL GND
.GLOBAL VDD


* Xconventional_pfd  ref VDD GND fb up dn conventional_pfd
* Xcp up VOP dn VDD GND CP_with_buffer 
* Vtest VOP lf_input DC 0 $ to measure the cuurent of the charge pump
* Xloop_filter_3rd_order lf_input vctrl GND loop_filter_3rd_order 

* *************************VCO********************
* xvco vp vn vctrl ibias VDD GND vco_sch
* xind1 vp vn ind_model
* XC_load vp vn sky130_fd_pr__cap_mim_m3_1 W=13 L=9 MF=1 m=1  $mim cap
* ** xbgr ibias GND VDD bgr_sch
* Isource VDD ibias 90u
* xinverter vp vco_out VDD GND vco_inverter     w_p=60 w_n=4.2 l=0.15
* xinverter2 vn fout_dummy VDD GND vco_inverter w_p=60 w_n=4.2 l=0.15
* *************************************************
* xdivider VDD fb GND p2 p7 p1 p6 p5 p4 p3 p0 vco_out float divider